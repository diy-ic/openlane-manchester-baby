magic
tech sky130A
magscale 1 2
timestamp 1700924122
<< viali >>
rect 13185 29257 13219 29291
rect 15669 29257 15703 29291
rect 18245 29257 18279 29291
rect 13093 29121 13127 29155
rect 15945 29121 15979 29155
rect 18521 29121 18555 29155
rect 14565 26945 14599 26979
rect 14749 26945 14783 26979
rect 15485 26945 15519 26979
rect 16957 26945 16991 26979
rect 17509 26877 17543 26911
rect 17969 26877 18003 26911
rect 18061 26877 18095 26911
rect 18705 26877 18739 26911
rect 17693 26809 17727 26843
rect 14657 26741 14691 26775
rect 15301 26741 15335 26775
rect 17141 26741 17175 26775
rect 19901 26537 19935 26571
rect 18613 26469 18647 26503
rect 15393 26401 15427 26435
rect 16313 26401 16347 26435
rect 19257 26401 19291 26435
rect 14105 26333 14139 26367
rect 15025 26333 15059 26367
rect 15301 26333 15335 26367
rect 15485 26333 15519 26367
rect 16221 26333 16255 26367
rect 17233 26333 17267 26367
rect 17489 26333 17523 26367
rect 14749 26265 14783 26299
rect 14841 26265 14875 26299
rect 15209 26197 15243 26231
rect 15577 26197 15611 26231
rect 16957 26197 16991 26231
rect 13093 25993 13127 26027
rect 14565 25993 14599 26027
rect 16221 25993 16255 26027
rect 18061 25993 18095 26027
rect 14228 25925 14262 25959
rect 16948 25925 16982 25959
rect 11888 25857 11922 25891
rect 14565 25857 14599 25891
rect 14749 25857 14783 25891
rect 14841 25857 14875 25891
rect 15108 25857 15142 25891
rect 16681 25857 16715 25891
rect 19717 25857 19751 25891
rect 11621 25789 11655 25823
rect 14473 25789 14507 25823
rect 19165 25789 19199 25823
rect 19257 25789 19291 25823
rect 13001 25653 13035 25687
rect 18521 25653 18555 25687
rect 19625 25653 19659 25687
rect 12817 25449 12851 25483
rect 13645 25449 13679 25483
rect 15301 25449 15335 25483
rect 18061 25381 18095 25415
rect 19257 25381 19291 25415
rect 10609 25313 10643 25347
rect 13001 25313 13035 25347
rect 17785 25313 17819 25347
rect 18797 25313 18831 25347
rect 9321 25245 9355 25279
rect 12909 25245 12943 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 17693 25245 17727 25279
rect 20637 25245 20671 25279
rect 10885 25177 10919 25211
rect 20370 25177 20404 25211
rect 9413 25109 9447 25143
rect 12357 25109 12391 25143
rect 18153 25109 18187 25143
rect 10977 24905 11011 24939
rect 11805 24905 11839 24939
rect 16948 24837 16982 24871
rect 10425 24769 10459 24803
rect 10609 24769 10643 24803
rect 10701 24769 10735 24803
rect 10793 24769 10827 24803
rect 11897 24769 11931 24803
rect 12265 24769 12299 24803
rect 14749 24769 14783 24803
rect 14841 24769 14875 24803
rect 16681 24769 16715 24803
rect 19073 24769 19107 24803
rect 6377 24701 6411 24735
rect 6653 24701 6687 24735
rect 8309 24701 8343 24735
rect 10057 24701 10091 24735
rect 10333 24701 10367 24735
rect 12817 24701 12851 24735
rect 13093 24701 13127 24735
rect 18705 24701 18739 24735
rect 14565 24633 14599 24667
rect 18061 24633 18095 24667
rect 8125 24565 8159 24599
rect 12081 24565 12115 24599
rect 18153 24565 18187 24599
rect 18889 24565 18923 24599
rect 6561 24361 6595 24395
rect 8401 24361 8435 24395
rect 9505 24361 9539 24395
rect 17049 24361 17083 24395
rect 18981 24361 19015 24395
rect 16773 24293 16807 24327
rect 18797 24293 18831 24327
rect 6469 24225 6503 24259
rect 10425 24225 10459 24259
rect 14565 24225 14599 24259
rect 16405 24225 16439 24259
rect 18521 24225 18555 24259
rect 6745 24157 6779 24191
rect 7113 24157 7147 24191
rect 8125 24157 8159 24191
rect 8493 24157 8527 24191
rect 8953 24157 8987 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 12449 24157 12483 24191
rect 13369 24157 13403 24191
rect 14289 24157 14323 24191
rect 18429 24157 18463 24191
rect 4445 24089 4479 24123
rect 6193 24089 6227 24123
rect 6837 24089 6871 24123
rect 6929 24089 6963 24123
rect 9137 24089 9171 24123
rect 10701 24089 10735 24123
rect 12357 24089 12391 24123
rect 14841 24089 14875 24123
rect 18162 24089 18196 24123
rect 7573 24021 7607 24055
rect 12173 24021 12207 24055
rect 13461 24021 13495 24055
rect 14473 24021 14507 24055
rect 16313 24021 16347 24055
rect 16865 24021 16899 24055
rect 5825 23817 5859 23851
rect 6377 23817 6411 23851
rect 7849 23817 7883 23851
rect 10517 23817 10551 23851
rect 14565 23817 14599 23851
rect 15577 23817 15611 23851
rect 6745 23749 6779 23783
rect 10149 23749 10183 23783
rect 18604 23749 18638 23783
rect 5917 23681 5951 23715
rect 6561 23681 6595 23715
rect 6653 23681 6687 23715
rect 6929 23681 6963 23715
rect 8125 23681 8159 23715
rect 8217 23681 8251 23715
rect 9965 23681 9999 23715
rect 10241 23681 10275 23715
rect 10333 23681 10367 23715
rect 13553 23681 13587 23715
rect 13737 23681 13771 23715
rect 14657 23681 14691 23715
rect 14841 23681 14875 23715
rect 15485 23681 15519 23715
rect 15945 23681 15979 23715
rect 20821 23681 20855 23715
rect 23489 23681 23523 23715
rect 14105 23613 14139 23647
rect 18337 23613 18371 23647
rect 24501 23613 24535 23647
rect 24777 23613 24811 23647
rect 14473 23545 14507 23579
rect 15761 23545 15795 23579
rect 8217 23477 8251 23511
rect 13553 23477 13587 23511
rect 14749 23477 14783 23511
rect 19717 23477 19751 23511
rect 20637 23477 20671 23511
rect 23581 23477 23615 23511
rect 26249 23477 26283 23511
rect 6377 23273 6411 23307
rect 9321 23273 9355 23307
rect 12081 23273 12115 23307
rect 13185 23273 13219 23307
rect 24961 23273 24995 23307
rect 25421 23273 25455 23307
rect 27721 23273 27755 23307
rect 7757 23205 7791 23239
rect 7849 23205 7883 23239
rect 8217 23205 8251 23239
rect 13001 23205 13035 23239
rect 6653 23137 6687 23171
rect 6745 23137 6779 23171
rect 12403 23137 12437 23171
rect 13553 23137 13587 23171
rect 20361 23137 20395 23171
rect 22477 23137 22511 23171
rect 6561 23069 6595 23103
rect 6837 23069 6871 23103
rect 7021 23069 7055 23103
rect 7665 23069 7699 23103
rect 7953 23069 7987 23103
rect 11989 23069 12023 23103
rect 12265 23069 12299 23103
rect 15117 23069 15151 23103
rect 15761 23069 15795 23103
rect 22385 23069 22419 23103
rect 25145 23069 25179 23103
rect 25329 23069 25363 23103
rect 27629 23069 27663 23103
rect 7113 23001 7147 23035
rect 8585 23001 8619 23035
rect 9505 23001 9539 23035
rect 20637 23001 20671 23035
rect 22293 23001 22327 23035
rect 22753 23001 22787 23035
rect 7481 22933 7515 22967
rect 8125 22933 8159 22967
rect 9137 22933 9171 22967
rect 9305 22933 9339 22967
rect 11805 22933 11839 22967
rect 12725 22933 12759 22967
rect 13185 22933 13219 22967
rect 14933 22933 14967 22967
rect 15669 22933 15703 22967
rect 22109 22933 22143 22967
rect 24225 22933 24259 22967
rect 28089 22933 28123 22967
rect 4445 22729 4479 22763
rect 6377 22729 6411 22763
rect 6653 22729 6687 22763
rect 7113 22729 7147 22763
rect 7757 22729 7791 22763
rect 9045 22729 9079 22763
rect 10517 22729 10551 22763
rect 10701 22729 10735 22763
rect 10793 22729 10827 22763
rect 12541 22729 12575 22763
rect 20729 22729 20763 22763
rect 21097 22729 21131 22763
rect 23029 22729 23063 22763
rect 23581 22729 23615 22763
rect 25145 22729 25179 22763
rect 25605 22729 25639 22763
rect 6193 22661 6227 22695
rect 9597 22661 9631 22695
rect 12357 22661 12391 22695
rect 14749 22661 14783 22695
rect 23949 22661 23983 22695
rect 28733 22661 28767 22695
rect 4077 22593 4111 22627
rect 4997 22593 5031 22627
rect 5457 22593 5491 22627
rect 5917 22593 5951 22627
rect 6009 22593 6043 22627
rect 6745 22593 6779 22627
rect 7021 22593 7055 22627
rect 7297 22593 7331 22627
rect 7665 22593 7699 22627
rect 7941 22593 7975 22627
rect 8401 22593 8435 22627
rect 8494 22593 8528 22627
rect 8677 22593 8711 22627
rect 8769 22593 8803 22627
rect 8866 22593 8900 22627
rect 9781 22593 9815 22627
rect 9965 22593 9999 22627
rect 10057 22593 10091 22627
rect 10977 22593 11011 22627
rect 11069 22593 11103 22627
rect 11253 22593 11287 22627
rect 11345 22593 11379 22627
rect 11529 22593 11563 22627
rect 11713 22593 11747 22627
rect 11805 22593 11839 22627
rect 11897 22593 11931 22627
rect 12015 22593 12049 22627
rect 12265 22593 12299 22627
rect 12442 22593 12476 22627
rect 12725 22593 12759 22627
rect 13001 22593 13035 22627
rect 14473 22593 14507 22627
rect 19533 22593 19567 22627
rect 23213 22593 23247 22627
rect 24041 22593 24075 22627
rect 25513 22593 25547 22627
rect 27997 22593 28031 22627
rect 28181 22593 28215 22627
rect 28457 22593 28491 22627
rect 28917 22593 28951 22627
rect 29193 22593 29227 22627
rect 29377 22593 29411 22627
rect 4169 22525 4203 22559
rect 4721 22525 4755 22559
rect 5273 22525 5307 22559
rect 5641 22525 5675 22559
rect 6536 22525 6570 22559
rect 8217 22525 8251 22559
rect 10149 22525 10183 22559
rect 12173 22525 12207 22559
rect 16497 22525 16531 22559
rect 16681 22525 16715 22559
rect 16957 22525 16991 22559
rect 19441 22525 19475 22559
rect 21189 22525 21223 22559
rect 21281 22525 21315 22559
rect 24133 22525 24167 22559
rect 25697 22525 25731 22559
rect 26341 22525 26375 22559
rect 26801 22525 26835 22559
rect 26985 22525 27019 22559
rect 6193 22457 6227 22491
rect 8125 22457 8159 22491
rect 19073 22457 19107 22491
rect 19809 22457 19843 22491
rect 26709 22457 26743 22491
rect 27261 22457 27295 22491
rect 4813 22389 4847 22423
rect 5181 22389 5215 22423
rect 7481 22389 7515 22423
rect 10517 22389 10551 22423
rect 12909 22389 12943 22423
rect 18429 22389 18463 22423
rect 18981 22389 19015 22423
rect 19993 22389 20027 22423
rect 27445 22389 27479 22423
rect 28641 22389 28675 22423
rect 29101 22389 29135 22423
rect 29285 22389 29319 22423
rect 4169 22185 4203 22219
rect 4905 22185 4939 22219
rect 8953 22185 8987 22219
rect 11621 22185 11655 22219
rect 15669 22185 15703 22219
rect 16957 22185 16991 22219
rect 18153 22185 18187 22219
rect 18981 22185 19015 22219
rect 19257 22185 19291 22219
rect 21465 22185 21499 22219
rect 25973 22185 26007 22219
rect 27905 22185 27939 22219
rect 17233 22117 17267 22151
rect 22293 22117 22327 22151
rect 25421 22117 25455 22151
rect 28089 22117 28123 22151
rect 29561 22117 29595 22151
rect 10517 22049 10551 22083
rect 13461 22049 13495 22083
rect 13670 22049 13704 22083
rect 17785 22049 17819 22083
rect 19717 22049 19751 22083
rect 22845 22049 22879 22083
rect 28733 22049 28767 22083
rect 29837 22049 29871 22083
rect 4353 21981 4387 22015
rect 4629 21981 4663 22015
rect 4721 21981 4755 22015
rect 4905 21981 4939 22015
rect 9137 21981 9171 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 9873 21981 9907 22015
rect 10425 21981 10459 22015
rect 12633 21981 12667 22015
rect 12817 21981 12851 22015
rect 13001 21981 13035 22015
rect 13185 21981 13219 22015
rect 14473 21981 14507 22015
rect 14749 21981 14783 22015
rect 15209 21981 15243 22015
rect 15485 21981 15519 22015
rect 17141 21981 17175 22015
rect 17601 21981 17635 22015
rect 18061 21981 18095 22015
rect 19073 21981 19107 22015
rect 19441 21981 19475 22015
rect 19533 21981 19567 22015
rect 19809 21981 19843 22015
rect 20545 21981 20579 22015
rect 20729 21981 20763 22015
rect 21649 21981 21683 22015
rect 22109 21981 22143 22015
rect 22753 21981 22787 22015
rect 22937 21981 22971 22015
rect 24409 21981 24443 22015
rect 24685 21981 24719 22015
rect 26157 21981 26191 22015
rect 26354 21981 26388 22015
rect 26571 21981 26605 22015
rect 26709 21981 26743 22015
rect 26893 21981 26927 22015
rect 27629 21981 27663 22015
rect 28641 21981 28675 22015
rect 28825 21981 28859 22015
rect 29101 21981 29135 22015
rect 29929 21981 29963 22015
rect 11805 21913 11839 21947
rect 11989 21913 12023 21947
rect 15301 21913 15335 21947
rect 20637 21913 20671 21947
rect 21189 21913 21223 21947
rect 21373 21913 21407 21947
rect 21741 21913 21775 21947
rect 21833 21913 21867 21947
rect 21971 21913 22005 21947
rect 22661 21913 22695 21947
rect 26249 21913 26283 21947
rect 26479 21913 26513 21947
rect 29285 21913 29319 21947
rect 4537 21845 4571 21879
rect 9321 21845 9355 21879
rect 9505 21845 9539 21879
rect 12541 21845 12575 21879
rect 13553 21845 13587 21879
rect 13829 21845 13863 21879
rect 17693 21845 17727 21879
rect 18613 21845 18647 21879
rect 21005 21845 21039 21879
rect 22201 21845 22235 21879
rect 26709 21845 26743 21879
rect 28917 21845 28951 21879
rect 5273 21641 5307 21675
rect 6929 21641 6963 21675
rect 9597 21641 9631 21675
rect 9689 21641 9723 21675
rect 10149 21641 10183 21675
rect 13185 21641 13219 21675
rect 15209 21641 15243 21675
rect 17509 21641 17543 21675
rect 19717 21641 19751 21675
rect 20085 21641 20119 21675
rect 23029 21641 23063 21675
rect 17877 21573 17911 21607
rect 18015 21573 18049 21607
rect 27813 21573 27847 21607
rect 1685 21505 1719 21539
rect 4813 21505 4847 21539
rect 5457 21505 5491 21539
rect 5733 21505 5767 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 6653 21505 6687 21539
rect 6745 21505 6779 21539
rect 9413 21505 9447 21539
rect 9505 21505 9539 21539
rect 10328 21505 10362 21539
rect 10425 21505 10459 21539
rect 10517 21505 10551 21539
rect 10700 21505 10734 21539
rect 10793 21505 10827 21539
rect 14013 21505 14047 21539
rect 15393 21505 15427 21539
rect 16681 21505 16715 21539
rect 17693 21505 17727 21539
rect 17785 21505 17819 21539
rect 18245 21505 18279 21539
rect 20269 21505 20303 21539
rect 20361 21505 20395 21539
rect 20545 21505 20579 21539
rect 21557 21505 21591 21539
rect 22937 21505 22971 21539
rect 23121 21505 23155 21539
rect 23673 21505 23707 21539
rect 25881 21505 25915 21539
rect 27353 21505 27387 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 4905 21437 4939 21471
rect 5641 21437 5675 21471
rect 9965 21437 9999 21471
rect 13645 21437 13679 21471
rect 14197 21437 14231 21471
rect 15025 21437 15059 21471
rect 15577 21437 15611 21471
rect 18153 21437 18187 21471
rect 21465 21437 21499 21471
rect 23857 21437 23891 21471
rect 25513 21437 25547 21471
rect 25605 21437 25639 21471
rect 27261 21437 27295 21471
rect 13369 21369 13403 21403
rect 26617 21369 26651 21403
rect 1501 21301 1535 21335
rect 5089 21301 5123 21335
rect 8125 21301 8159 21335
rect 13829 21301 13863 21335
rect 14473 21301 14507 21335
rect 16773 21301 16807 21335
rect 20545 21301 20579 21335
rect 21189 21301 21223 21335
rect 21373 21301 21407 21335
rect 26985 21301 27019 21335
rect 27261 21301 27295 21335
rect 5733 21097 5767 21131
rect 8033 21097 8067 21131
rect 9689 21097 9723 21131
rect 10517 21097 10551 21131
rect 10701 21097 10735 21131
rect 11989 21097 12023 21131
rect 12173 21097 12207 21131
rect 12817 21097 12851 21131
rect 14841 21097 14875 21131
rect 19441 21097 19475 21131
rect 23581 21097 23615 21131
rect 23765 21097 23799 21131
rect 27261 21097 27295 21131
rect 28089 21097 28123 21131
rect 6929 21029 6963 21063
rect 9229 21029 9263 21063
rect 9873 21029 9907 21063
rect 10241 21029 10275 21063
rect 12633 21029 12667 21063
rect 18705 21029 18739 21063
rect 22293 21029 22327 21063
rect 23029 21029 23063 21063
rect 27445 21029 27479 21063
rect 5365 20961 5399 20995
rect 7021 20961 7055 20995
rect 7573 20961 7607 20995
rect 7849 20961 7883 20995
rect 11345 20961 11379 20995
rect 14197 20961 14231 20995
rect 15577 20961 15611 20995
rect 15669 20961 15703 20995
rect 19257 20961 19291 20995
rect 19809 20961 19843 20995
rect 20729 20961 20763 20995
rect 23489 20961 23523 20995
rect 24869 20961 24903 20995
rect 26709 20961 26743 20995
rect 27629 20961 27663 20995
rect 27721 20961 27755 20995
rect 27813 20961 27847 20995
rect 1685 20893 1719 20927
rect 5089 20893 5123 20927
rect 5535 20893 5569 20927
rect 6469 20893 6503 20927
rect 6653 20893 6687 20927
rect 6745 20893 6779 20927
rect 6837 20893 6871 20927
rect 7481 20893 7515 20927
rect 8217 20893 8251 20927
rect 8401 20893 8435 20927
rect 8585 20893 8619 20927
rect 8953 20893 8987 20927
rect 9413 20893 9447 20927
rect 9965 20893 9999 20927
rect 10057 20893 10091 20927
rect 10333 20893 10367 20927
rect 10517 20893 10551 20927
rect 10885 20893 10919 20927
rect 11805 20893 11839 20927
rect 12541 20893 12575 20927
rect 13185 20893 13219 20927
rect 14565 20893 14599 20927
rect 14657 20893 14691 20927
rect 14933 20893 14967 20927
rect 18613 20893 18647 20927
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 19073 20893 19107 20927
rect 19717 20893 19751 20927
rect 22661 20893 22695 20927
rect 22937 20893 22971 20927
rect 23305 20893 23339 20927
rect 26801 20893 26835 20927
rect 26985 20893 27019 20927
rect 27905 20893 27939 20927
rect 28365 20893 28399 20927
rect 28549 20893 28583 20927
rect 28641 20893 28675 20927
rect 8309 20825 8343 20859
rect 9045 20825 9079 20859
rect 9505 20825 9539 20859
rect 10241 20825 10275 20859
rect 10977 20825 11011 20859
rect 11069 20825 11103 20859
rect 11187 20825 11221 20859
rect 11621 20825 11655 20859
rect 12817 20825 12851 20859
rect 14289 20825 14323 20859
rect 15945 20825 15979 20859
rect 17693 20825 17727 20859
rect 19993 20825 20027 20859
rect 21925 20825 21959 20859
rect 22477 20825 22511 20859
rect 22845 20825 22879 20859
rect 23949 20825 23983 20859
rect 25053 20825 25087 20859
rect 27077 20825 27111 20859
rect 28181 20825 28215 20859
rect 1501 20757 1535 20791
rect 4537 20757 4571 20791
rect 6561 20757 6595 20791
rect 9705 20757 9739 20791
rect 11437 20757 11471 20791
rect 12173 20757 12207 20791
rect 14381 20757 14415 20791
rect 18429 20757 18463 20791
rect 22385 20757 22419 20791
rect 23749 20757 23783 20791
rect 26985 20757 27019 20791
rect 27277 20757 27311 20791
rect 4261 20553 4295 20587
rect 4721 20553 4755 20587
rect 7573 20553 7607 20587
rect 11529 20553 11563 20587
rect 12081 20553 12115 20587
rect 16221 20553 16255 20587
rect 16681 20553 16715 20587
rect 20085 20553 20119 20587
rect 22845 20553 22879 20587
rect 28549 20553 28583 20587
rect 4813 20485 4847 20519
rect 5457 20485 5491 20519
rect 7757 20485 7791 20519
rect 12633 20485 12667 20519
rect 13001 20485 13035 20519
rect 14197 20485 14231 20519
rect 15853 20485 15887 20519
rect 19441 20485 19475 20519
rect 28917 20485 28951 20519
rect 29653 20485 29687 20519
rect 12403 20451 12437 20485
rect 5365 20417 5399 20451
rect 5549 20417 5583 20451
rect 5733 20417 5767 20451
rect 6929 20417 6963 20451
rect 7113 20417 7147 20451
rect 7297 20417 7331 20451
rect 7389 20417 7423 20451
rect 7573 20417 7607 20451
rect 7665 20417 7699 20451
rect 7849 20417 7883 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 11989 20417 12023 20451
rect 12173 20417 12207 20451
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 13277 20417 13311 20451
rect 13829 20417 13863 20451
rect 13921 20417 13955 20451
rect 15761 20417 15795 20451
rect 16405 20417 16439 20451
rect 17049 20417 17083 20451
rect 18705 20417 18739 20451
rect 18981 20417 19015 20451
rect 19165 20417 19199 20451
rect 19257 20417 19291 20451
rect 20821 20417 20855 20451
rect 22109 20417 22143 20451
rect 23305 20417 23339 20451
rect 23581 20417 23615 20451
rect 23857 20417 23891 20451
rect 24869 20417 24903 20451
rect 28733 20417 28767 20451
rect 28825 20417 28859 20451
rect 29101 20417 29135 20451
rect 29193 20407 29227 20441
rect 29469 20417 29503 20451
rect 29745 20417 29779 20451
rect 29837 20417 29871 20451
rect 2513 20349 2547 20383
rect 2789 20349 2823 20383
rect 4997 20349 5031 20383
rect 15669 20349 15703 20383
rect 17141 20349 17175 20383
rect 17325 20349 17359 20383
rect 18797 20349 18831 20383
rect 21097 20349 21131 20383
rect 21833 20349 21867 20383
rect 22937 20349 22971 20383
rect 5181 20281 5215 20315
rect 18889 20281 18923 20315
rect 23397 20281 23431 20315
rect 4353 20213 4387 20247
rect 12265 20213 12299 20247
rect 12449 20213 12483 20247
rect 12725 20213 12759 20247
rect 13645 20213 13679 20247
rect 19625 20213 19659 20247
rect 24961 20213 24995 20247
rect 29285 20213 29319 20247
rect 29929 20213 29963 20247
rect 30297 20213 30331 20247
rect 3065 20009 3099 20043
rect 3893 20009 3927 20043
rect 8217 20009 8251 20043
rect 11161 20009 11195 20043
rect 13093 20009 13127 20043
rect 17141 20009 17175 20043
rect 17233 20009 17267 20043
rect 19349 20009 19383 20043
rect 20177 20009 20211 20043
rect 23397 20009 23431 20043
rect 27997 20009 28031 20043
rect 28181 20009 28215 20043
rect 28733 20009 28767 20043
rect 8953 19941 8987 19975
rect 11069 19941 11103 19975
rect 24777 19941 24811 19975
rect 28549 19941 28583 19975
rect 29101 19941 29135 19975
rect 29193 19941 29227 19975
rect 7481 19873 7515 19907
rect 9597 19873 9631 19907
rect 10609 19873 10643 19907
rect 11621 19873 11655 19907
rect 16405 19873 16439 19907
rect 17141 19873 17175 19907
rect 21005 19873 21039 19907
rect 21189 19873 21223 19907
rect 22937 19873 22971 19907
rect 25329 19873 25363 19907
rect 25605 19873 25639 19907
rect 27445 19873 27479 19907
rect 28917 19873 28951 19907
rect 29009 19873 29043 19907
rect 1685 19805 1719 19839
rect 3249 19805 3283 19839
rect 3985 19805 4019 19839
rect 4905 19805 4939 19839
rect 5273 19805 5307 19839
rect 7757 19805 7791 19839
rect 8125 19805 8159 19839
rect 8401 19805 8435 19839
rect 9137 19805 9171 19839
rect 9505 19805 9539 19839
rect 10241 19805 10275 19839
rect 10701 19805 10735 19839
rect 11529 19805 11563 19839
rect 12541 19805 12575 19839
rect 12725 19805 12759 19839
rect 12909 19805 12943 19839
rect 16037 19805 16071 19839
rect 16221 19805 16255 19839
rect 17325 19805 17359 19839
rect 18613 19805 18647 19839
rect 18797 19805 18831 19839
rect 19441 19805 19475 19839
rect 19901 19805 19935 19839
rect 20453 19805 20487 19839
rect 20637 19805 20671 19839
rect 20821 19805 20855 19839
rect 22845 19805 22879 19839
rect 23305 19805 23339 19839
rect 23581 19805 23615 19839
rect 23857 19805 23891 19839
rect 24685 19805 24719 19839
rect 25145 19805 25179 19839
rect 27721 19805 27755 19839
rect 28273 19805 28307 19839
rect 29283 19783 29317 19817
rect 4997 19737 5031 19771
rect 5089 19737 5123 19771
rect 7849 19737 7883 19771
rect 7941 19737 7975 19771
rect 9229 19737 9263 19771
rect 9321 19737 9355 19771
rect 12817 19737 12851 19771
rect 16957 19737 16991 19771
rect 25789 19737 25823 19771
rect 1501 19669 1535 19703
rect 4721 19669 4755 19703
rect 6837 19669 6871 19703
rect 7573 19669 7607 19703
rect 18705 19669 18739 19703
rect 24501 19669 24535 19703
rect 25237 19669 25271 19703
rect 6377 19465 6411 19499
rect 6745 19465 6779 19499
rect 9781 19465 9815 19499
rect 17417 19465 17451 19499
rect 19441 19465 19475 19499
rect 26157 19465 26191 19499
rect 29469 19465 29503 19499
rect 7849 19397 7883 19431
rect 14473 19397 14507 19431
rect 17049 19397 17083 19431
rect 18981 19397 19015 19431
rect 24317 19397 24351 19431
rect 26525 19397 26559 19431
rect 26663 19397 26697 19431
rect 1685 19329 1719 19363
rect 5733 19329 5767 19363
rect 6837 19329 6871 19363
rect 7573 19329 7607 19363
rect 12449 19329 12483 19363
rect 12541 19329 12575 19363
rect 12633 19329 12667 19363
rect 14289 19329 14323 19363
rect 16221 19329 16255 19363
rect 16405 19329 16439 19363
rect 16931 19329 16965 19363
rect 17141 19329 17175 19363
rect 17233 19329 17267 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 18153 19329 18187 19363
rect 18245 19329 18279 19363
rect 18363 19329 18397 19363
rect 18797 19329 18831 19363
rect 19073 19329 19107 19363
rect 19257 19329 19291 19363
rect 20085 19329 20119 19363
rect 20361 19329 20395 19363
rect 20637 19329 20671 19363
rect 21005 19329 21039 19363
rect 21097 19329 21131 19363
rect 22565 19329 22599 19363
rect 23029 19329 23063 19363
rect 23305 19329 23339 19363
rect 23489 19329 23523 19363
rect 24041 19329 24075 19363
rect 26341 19329 26375 19363
rect 26433 19329 26467 19363
rect 27261 19329 27295 19363
rect 29101 19329 29135 19363
rect 29193 19329 29227 19363
rect 29377 19329 29411 19363
rect 29837 19329 29871 19363
rect 30113 19329 30147 19363
rect 30297 19329 30331 19363
rect 4997 19261 5031 19295
rect 7021 19261 7055 19295
rect 9321 19261 9355 19295
rect 9873 19261 9907 19295
rect 9965 19261 9999 19295
rect 14013 19261 14047 19295
rect 15117 19261 15151 19295
rect 16773 19261 16807 19295
rect 18521 19261 18555 19295
rect 21189 19261 21223 19295
rect 21649 19261 21683 19295
rect 23397 19261 23431 19295
rect 25789 19261 25823 19295
rect 26801 19261 26835 19295
rect 26985 19261 27019 19295
rect 29929 19261 29963 19295
rect 30205 19261 30239 19295
rect 9413 19193 9447 19227
rect 16221 19193 16255 19227
rect 18613 19193 18647 19227
rect 1501 19125 1535 19159
rect 4445 19125 4479 19159
rect 5549 19125 5583 19159
rect 13369 19125 13403 19159
rect 27997 19125 28031 19159
rect 28917 19125 28951 19159
rect 29101 19125 29135 19159
rect 6837 18921 6871 18955
rect 8677 18921 8711 18955
rect 13921 18921 13955 18955
rect 16313 18921 16347 18955
rect 17325 18921 17359 18955
rect 17601 18921 17635 18955
rect 18061 18921 18095 18955
rect 19073 18921 19107 18955
rect 19257 18921 19291 18955
rect 27537 18921 27571 18955
rect 12081 18853 12115 18887
rect 15669 18853 15703 18887
rect 18981 18853 19015 18887
rect 19349 18853 19383 18887
rect 29285 18853 29319 18887
rect 4537 18785 4571 18819
rect 5089 18785 5123 18819
rect 12173 18785 12207 18819
rect 12449 18785 12483 18819
rect 16037 18785 16071 18819
rect 17233 18785 17267 18819
rect 18613 18785 18647 18819
rect 22569 18785 22603 18819
rect 23397 18785 23431 18819
rect 27997 18785 28031 18819
rect 28641 18785 28675 18819
rect 1685 18717 1719 18751
rect 3341 18717 3375 18751
rect 3617 18717 3651 18751
rect 8585 18717 8619 18751
rect 11897 18717 11931 18751
rect 14289 18717 14323 18751
rect 14657 18717 14691 18751
rect 14933 18717 14967 18751
rect 15945 18717 15979 18751
rect 17141 18717 17175 18751
rect 17417 18717 17451 18751
rect 17877 18717 17911 18751
rect 18061 18717 18095 18751
rect 19717 18717 19751 18751
rect 20177 18717 20211 18751
rect 23029 18717 23063 18751
rect 23213 18717 23247 18751
rect 23489 18717 23523 18751
rect 24593 18717 24627 18751
rect 27445 18717 27479 18751
rect 27629 18717 27663 18751
rect 28089 18717 28123 18751
rect 28181 18717 28215 18751
rect 28273 18717 28307 18751
rect 28549 18717 28583 18751
rect 28733 18717 28767 18751
rect 4261 18649 4295 18683
rect 5365 18649 5399 18683
rect 14197 18649 14231 18683
rect 20453 18649 20487 18683
rect 28917 18649 28951 18683
rect 29101 18649 29135 18683
rect 1501 18581 1535 18615
rect 3157 18581 3191 18615
rect 3525 18581 3559 18615
rect 3893 18581 3927 18615
rect 4353 18581 4387 18615
rect 24409 18581 24443 18615
rect 27813 18581 27847 18615
rect 4445 18377 4479 18411
rect 6101 18377 6135 18411
rect 12357 18377 12391 18411
rect 12725 18377 12759 18411
rect 25789 18377 25823 18411
rect 26249 18377 26283 18411
rect 28457 18377 28491 18411
rect 29193 18377 29227 18411
rect 2973 18309 3007 18343
rect 10241 18309 10275 18343
rect 24225 18309 24259 18343
rect 28089 18309 28123 18343
rect 28289 18309 28323 18343
rect 2697 18241 2731 18275
rect 6009 18241 6043 18275
rect 7021 18241 7055 18275
rect 8953 18241 8987 18275
rect 9137 18241 9171 18275
rect 9597 18241 9631 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 9899 18241 9933 18275
rect 10149 18241 10183 18275
rect 10333 18241 10367 18275
rect 11897 18241 11931 18275
rect 12817 18241 12851 18275
rect 14013 18241 14047 18275
rect 14197 18241 14231 18275
rect 14565 18241 14599 18275
rect 14933 18241 14967 18275
rect 15209 18241 15243 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 16957 18241 16991 18275
rect 19717 18241 19751 18275
rect 19993 18241 20027 18275
rect 20821 18241 20855 18275
rect 20913 18241 20947 18275
rect 21189 18241 21223 18275
rect 21833 18241 21867 18275
rect 22201 18241 22235 18275
rect 22477 18241 22511 18275
rect 22845 18241 22879 18275
rect 23949 18241 23983 18275
rect 26157 18241 26191 18275
rect 26985 18241 27019 18275
rect 27261 18241 27295 18275
rect 29193 18241 29227 18275
rect 29377 18241 29411 18275
rect 6745 18173 6779 18207
rect 9321 18173 9355 18207
rect 10057 18173 10091 18207
rect 10517 18173 10551 18207
rect 11805 18173 11839 18207
rect 12909 18173 12943 18207
rect 14473 18173 14507 18207
rect 15945 18173 15979 18207
rect 20269 18173 20303 18207
rect 25697 18173 25731 18207
rect 26341 18173 26375 18207
rect 6837 18105 6871 18139
rect 10793 18105 10827 18139
rect 11529 18105 11563 18139
rect 6929 18037 6963 18071
rect 9413 18037 9447 18071
rect 10977 18037 11011 18071
rect 16773 18037 16807 18071
rect 20729 18037 20763 18071
rect 22569 18037 22603 18071
rect 27997 18037 28031 18071
rect 28273 18037 28307 18071
rect 6377 17833 6411 17867
rect 6561 17833 6595 17867
rect 10517 17833 10551 17867
rect 11069 17833 11103 17867
rect 11437 17833 11471 17867
rect 19073 17833 19107 17867
rect 24869 17833 24903 17867
rect 27537 17833 27571 17867
rect 28089 17833 28123 17867
rect 28825 17833 28859 17867
rect 29193 17833 29227 17867
rect 29653 17833 29687 17867
rect 30021 17833 30055 17867
rect 11529 17765 11563 17799
rect 13001 17765 13035 17799
rect 17969 17765 18003 17799
rect 5549 17697 5583 17731
rect 7205 17697 7239 17731
rect 7481 17697 7515 17731
rect 8493 17697 8527 17731
rect 10885 17697 10919 17731
rect 16221 17697 16255 17731
rect 16497 17697 16531 17731
rect 19717 17697 19751 17731
rect 22569 17697 22603 17731
rect 23397 17697 23431 17731
rect 25789 17697 25823 17731
rect 27353 17697 27387 17731
rect 3801 17629 3835 17663
rect 6101 17629 6135 17663
rect 6653 17629 6687 17663
rect 6837 17629 6871 17663
rect 7113 17629 7147 17663
rect 8033 17629 8067 17663
rect 8217 17629 8251 17663
rect 8335 17629 8369 17663
rect 8585 17629 8619 17663
rect 8769 17629 8803 17663
rect 9321 17629 9355 17663
rect 10425 17629 10459 17663
rect 10977 17629 11011 17663
rect 11713 17629 11747 17663
rect 11805 17629 11839 17663
rect 12817 17629 12851 17663
rect 13185 17629 13219 17663
rect 18061 17629 18095 17663
rect 18337 17629 18371 17663
rect 19257 17629 19291 17663
rect 23029 17629 23063 17663
rect 23305 17629 23339 17663
rect 23581 17629 23615 17663
rect 24777 17629 24811 17663
rect 25605 17629 25639 17663
rect 27905 17629 27939 17663
rect 27997 17629 28031 17663
rect 28181 17629 28215 17663
rect 28733 17629 28767 17663
rect 29561 17629 29595 17663
rect 4077 17561 4111 17595
rect 6745 17561 6779 17595
rect 8125 17561 8159 17595
rect 8953 17561 8987 17595
rect 9137 17561 9171 17595
rect 11529 17561 11563 17595
rect 12633 17561 12667 17595
rect 19441 17561 19475 17595
rect 27721 17561 27755 17595
rect 7849 17493 7883 17527
rect 8585 17493 8619 17527
rect 4169 17289 4203 17323
rect 4537 17289 4571 17323
rect 4721 17289 4755 17323
rect 5089 17289 5123 17323
rect 6837 17289 6871 17323
rect 9689 17289 9723 17323
rect 12173 17289 12207 17323
rect 15577 17289 15611 17323
rect 17049 17289 17083 17323
rect 17233 17289 17267 17323
rect 17693 17289 17727 17323
rect 25513 17289 25547 17323
rect 27353 17289 27387 17323
rect 5181 17221 5215 17255
rect 17601 17221 17635 17255
rect 20361 17221 20395 17255
rect 23489 17221 23523 17255
rect 4353 17153 4387 17187
rect 4445 17153 4479 17187
rect 6377 17153 6411 17187
rect 7113 17153 7147 17187
rect 7205 17153 7239 17187
rect 9597 17153 9631 17187
rect 11529 17153 11563 17187
rect 12265 17153 12299 17187
rect 12357 17153 12391 17187
rect 12633 17153 12667 17187
rect 13461 17153 13495 17187
rect 15485 17153 15519 17187
rect 16037 17153 16071 17187
rect 16957 17153 16991 17187
rect 19349 17153 19383 17187
rect 19533 17153 19567 17187
rect 20085 17153 20119 17187
rect 20545 17153 20579 17187
rect 20821 17153 20855 17187
rect 21005 17153 21039 17187
rect 23673 17153 23707 17187
rect 23765 17153 23799 17187
rect 27537 17153 27571 17187
rect 27813 17153 27847 17187
rect 5273 17085 5307 17119
rect 9781 17085 9815 17119
rect 11805 17085 11839 17119
rect 13553 17085 13587 17119
rect 13829 17085 13863 17119
rect 15301 17085 15335 17119
rect 17877 17085 17911 17119
rect 23121 17085 23155 17119
rect 24041 17085 24075 17119
rect 27721 17085 27755 17119
rect 6469 16949 6503 16983
rect 7297 16949 7331 16983
rect 7481 16949 7515 16983
rect 9229 16949 9263 16983
rect 16129 16949 16163 16983
rect 27721 16949 27755 16983
rect 10977 16745 11011 16779
rect 11713 16745 11747 16779
rect 11897 16745 11931 16779
rect 14105 16745 14139 16779
rect 14657 16745 14691 16779
rect 15301 16745 15335 16779
rect 18981 16745 19015 16779
rect 28641 16745 28675 16779
rect 5825 16677 5859 16711
rect 18337 16677 18371 16711
rect 4261 16609 4295 16643
rect 4445 16609 4479 16643
rect 6929 16609 6963 16643
rect 9229 16609 9263 16643
rect 12081 16609 12115 16643
rect 12633 16609 12667 16643
rect 15669 16609 15703 16643
rect 19349 16609 19383 16643
rect 19533 16609 19567 16643
rect 20453 16609 20487 16643
rect 21925 16609 21959 16643
rect 22385 16609 22419 16643
rect 24133 16609 24167 16643
rect 24501 16609 24535 16643
rect 24777 16609 24811 16643
rect 7021 16541 7055 16575
rect 8493 16541 8527 16575
rect 8677 16541 8711 16575
rect 8953 16541 8987 16575
rect 11069 16541 11103 16575
rect 11437 16541 11471 16575
rect 14289 16541 14323 16575
rect 14565 16541 14599 16575
rect 15025 16541 15059 16575
rect 15485 16541 15519 16575
rect 19265 16541 19299 16575
rect 22661 16541 22695 16575
rect 26341 16541 26375 16575
rect 28181 16541 28215 16575
rect 5457 16473 5491 16507
rect 9505 16473 9539 16507
rect 11161 16473 11195 16507
rect 12265 16473 12299 16507
rect 18153 16473 18187 16507
rect 18705 16473 18739 16507
rect 20637 16473 20671 16507
rect 23857 16473 23891 16507
rect 26525 16473 26559 16507
rect 28273 16473 28307 16507
rect 28457 16473 28491 16507
rect 3801 16405 3835 16439
rect 4169 16405 4203 16439
rect 5917 16405 5951 16439
rect 7389 16405 7423 16439
rect 8493 16405 8527 16439
rect 9137 16405 9171 16439
rect 14841 16405 14875 16439
rect 19717 16405 19751 16439
rect 23397 16405 23431 16439
rect 23489 16405 23523 16439
rect 23949 16405 23983 16439
rect 26249 16405 26283 16439
rect 3801 16201 3835 16235
rect 6193 16201 6227 16235
rect 13737 16201 13771 16235
rect 18429 16201 18463 16235
rect 18613 16201 18647 16235
rect 23213 16201 23247 16235
rect 25053 16201 25087 16235
rect 25421 16201 25455 16235
rect 25605 16201 25639 16235
rect 8309 16133 8343 16167
rect 12265 16133 12299 16167
rect 16037 16133 16071 16167
rect 17601 16133 17635 16167
rect 23949 16133 23983 16167
rect 4077 16065 4111 16099
rect 4445 16065 4479 16099
rect 5457 16065 5491 16099
rect 6009 16065 6043 16099
rect 6193 16065 6227 16099
rect 6469 16065 6503 16099
rect 6561 16065 6595 16099
rect 6745 16065 6779 16099
rect 8125 16065 8159 16099
rect 8217 16065 8251 16099
rect 8427 16065 8461 16099
rect 8585 16065 8619 16099
rect 8953 16065 8987 16099
rect 11345 16065 11379 16099
rect 14105 16065 14139 16099
rect 16129 16065 16163 16099
rect 16957 16065 16991 16099
rect 17693 16065 17727 16099
rect 17785 16065 17819 16099
rect 20269 16065 20303 16099
rect 20637 16065 20671 16099
rect 20913 16065 20947 16099
rect 23029 16065 23063 16099
rect 23857 16065 23891 16099
rect 25237 16065 25271 16099
rect 25329 16065 25363 16099
rect 25973 16065 26007 16099
rect 26985 16065 27019 16099
rect 27261 16065 27295 16099
rect 28089 16065 28123 16099
rect 28273 16065 28307 16099
rect 2053 15997 2087 16031
rect 2329 15997 2363 16031
rect 3985 15997 4019 16031
rect 4169 15997 4203 16031
rect 5917 15997 5951 16031
rect 6653 15997 6687 16031
rect 11161 15997 11195 16031
rect 14381 15997 14415 16031
rect 18153 15997 18187 16031
rect 18337 15997 18371 16031
rect 26065 15997 26099 16031
rect 26157 15997 26191 16031
rect 7941 15929 7975 15963
rect 15853 15929 15887 15963
rect 18981 15929 19015 15963
rect 27997 15929 28031 15963
rect 5191 15861 5225 15895
rect 5733 15861 5767 15895
rect 6929 15861 6963 15895
rect 8769 15861 8803 15895
rect 17049 15861 17083 15895
rect 18621 15861 18655 15895
rect 20177 15861 20211 15895
rect 21649 15861 21683 15895
rect 28181 15861 28215 15895
rect 2513 15657 2547 15691
rect 5917 15657 5951 15691
rect 6101 15657 6135 15691
rect 8953 15657 8987 15691
rect 9413 15657 9447 15691
rect 12173 15657 12207 15691
rect 13829 15657 13863 15691
rect 14841 15657 14875 15691
rect 17785 15657 17819 15691
rect 18429 15657 18463 15691
rect 19514 15657 19548 15691
rect 21005 15657 21039 15691
rect 22569 15657 22603 15691
rect 23029 15657 23063 15691
rect 23305 15657 23339 15691
rect 24133 15657 24167 15691
rect 25237 15657 25271 15691
rect 26341 15657 26375 15691
rect 19073 15589 19107 15623
rect 24961 15589 24995 15623
rect 4445 15521 4479 15555
rect 5825 15521 5859 15555
rect 7021 15521 7055 15555
rect 9137 15521 9171 15555
rect 10885 15521 10919 15555
rect 13921 15521 13955 15555
rect 14197 15521 14231 15555
rect 15301 15521 15335 15555
rect 15485 15521 15519 15555
rect 19257 15521 19291 15555
rect 22753 15521 22787 15555
rect 23857 15521 23891 15555
rect 26433 15521 26467 15555
rect 27169 15521 27203 15555
rect 2697 15453 2731 15487
rect 6377 15453 6411 15487
rect 6561 15453 6595 15487
rect 8953 15453 8987 15487
rect 9229 15453 9263 15487
rect 9781 15453 9815 15487
rect 10609 15453 10643 15487
rect 11069 15453 11103 15487
rect 11805 15453 11839 15487
rect 11897 15453 11931 15487
rect 12449 15453 12483 15487
rect 13093 15453 13127 15487
rect 13277 15453 13311 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 16037 15453 16071 15487
rect 18521 15453 18555 15487
rect 18889 15453 18923 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 22293 15453 22327 15487
rect 22477 15453 22511 15487
rect 22845 15453 22879 15487
rect 23673 15453 23707 15487
rect 23765 15453 23799 15487
rect 23949 15453 23983 15487
rect 24593 15453 24627 15487
rect 25145 15453 25179 15487
rect 26157 15453 26191 15487
rect 26249 15453 26283 15487
rect 27353 15453 27387 15487
rect 27537 15453 27571 15487
rect 27629 15453 27663 15487
rect 5641 15385 5675 15419
rect 6745 15385 6779 15419
rect 11529 15385 11563 15419
rect 14473 15385 14507 15419
rect 16313 15385 16347 15419
rect 22569 15385 22603 15419
rect 23121 15385 23155 15419
rect 23321 15385 23355 15419
rect 11161 15317 11195 15351
rect 14381 15317 14415 15351
rect 15577 15317 15611 15351
rect 15945 15317 15979 15351
rect 21465 15317 21499 15351
rect 22477 15317 22511 15351
rect 23489 15317 23523 15351
rect 25053 15317 25087 15351
rect 25605 15317 25639 15351
rect 6009 15113 6043 15147
rect 8493 15113 8527 15147
rect 14933 15113 14967 15147
rect 16037 15113 16071 15147
rect 17969 15113 18003 15147
rect 19717 15113 19751 15147
rect 20085 15113 20119 15147
rect 25697 15113 25731 15147
rect 26525 15113 26559 15147
rect 3617 15045 3651 15079
rect 11989 15045 12023 15079
rect 12081 15045 12115 15079
rect 12219 15045 12253 15079
rect 17693 15045 17727 15079
rect 18245 15045 18279 15079
rect 19441 15045 19475 15079
rect 21281 15045 21315 15079
rect 21419 15045 21453 15079
rect 22477 15045 22511 15079
rect 3525 14977 3559 15011
rect 5917 14977 5951 15011
rect 7757 14977 7791 15011
rect 9505 14977 9539 15011
rect 11713 14977 11747 15011
rect 11897 14977 11931 15011
rect 13553 14977 13587 15011
rect 14105 14977 14139 15011
rect 14749 14977 14783 15011
rect 15117 14977 15151 15011
rect 15853 14977 15887 15011
rect 18797 14977 18831 15011
rect 20177 14977 20211 15011
rect 20913 14977 20947 15011
rect 21097 14977 21131 15011
rect 21189 14977 21223 15011
rect 21557 14977 21591 15011
rect 21833 14977 21867 15011
rect 22015 14977 22049 15011
rect 22293 14977 22327 15011
rect 25605 14977 25639 15011
rect 25881 14977 25915 15011
rect 26065 14977 26099 15011
rect 26157 14977 26191 15011
rect 27261 14977 27295 15011
rect 27813 14977 27847 15011
rect 3801 14909 3835 14943
rect 7481 14909 7515 14943
rect 9689 14909 9723 14943
rect 9965 14909 9999 14943
rect 12357 14909 12391 14943
rect 12449 14909 12483 14943
rect 13001 14909 13035 14943
rect 13369 14909 13403 14943
rect 13461 14909 13495 14943
rect 20269 14909 20303 14943
rect 26249 14909 26283 14943
rect 26341 14909 26375 14943
rect 13921 14841 13955 14875
rect 18981 14841 19015 14875
rect 19257 14841 19291 14875
rect 22201 14841 22235 14875
rect 25881 14841 25915 14875
rect 27629 14841 27663 14875
rect 3157 14773 3191 14807
rect 14197 14773 14231 14807
rect 15301 14773 15335 14807
rect 18521 14773 18555 14807
rect 22661 14773 22695 14807
rect 27721 14773 27755 14807
rect 27905 14773 27939 14807
rect 28273 14773 28307 14807
rect 3617 14569 3651 14603
rect 4537 14569 4571 14603
rect 6653 14569 6687 14603
rect 9781 14569 9815 14603
rect 10780 14569 10814 14603
rect 13001 14569 13035 14603
rect 13369 14569 13403 14603
rect 21465 14569 21499 14603
rect 22937 14569 22971 14603
rect 23673 14569 23707 14603
rect 24409 14569 24443 14603
rect 26065 14569 26099 14603
rect 27445 14569 27479 14603
rect 27721 14569 27755 14603
rect 21833 14501 21867 14535
rect 22569 14501 22603 14535
rect 23489 14501 23523 14535
rect 25789 14501 25823 14535
rect 7389 14433 7423 14467
rect 12265 14433 12299 14467
rect 17233 14433 17267 14467
rect 17417 14433 17451 14467
rect 19993 14433 20027 14467
rect 22293 14433 22327 14467
rect 27169 14433 27203 14467
rect 27261 14433 27295 14467
rect 1869 14365 1903 14399
rect 4077 14365 4111 14399
rect 4445 14365 4479 14399
rect 4813 14365 4847 14399
rect 5089 14365 5123 14399
rect 6009 14365 6043 14399
rect 6285 14365 6319 14399
rect 6561 14365 6595 14399
rect 6929 14365 6963 14399
rect 7481 14365 7515 14399
rect 8309 14365 8343 14399
rect 9321 14365 9355 14399
rect 9689 14365 9723 14399
rect 9965 14365 9999 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 12541 14365 12575 14399
rect 12817 14365 12851 14399
rect 13461 14365 13495 14399
rect 13737 14365 13771 14399
rect 14197 14365 14231 14399
rect 16037 14365 16071 14399
rect 16957 14365 16991 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 18429 14365 18463 14399
rect 19073 14365 19107 14399
rect 19717 14365 19751 14399
rect 19809 14365 19843 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22845 14365 22879 14399
rect 23949 14365 23983 14399
rect 24593 14365 24627 14399
rect 24777 14365 24811 14399
rect 24934 14365 24968 14399
rect 25053 14365 25087 14399
rect 25145 14375 25179 14409
rect 25237 14365 25271 14399
rect 25605 14365 25639 14399
rect 26341 14365 26375 14399
rect 26985 14365 27019 14399
rect 27077 14365 27111 14399
rect 27905 14365 27939 14399
rect 21511 14331 21545 14365
rect 2145 14297 2179 14331
rect 7757 14297 7791 14331
rect 8033 14297 8067 14331
rect 8125 14297 8159 14331
rect 14381 14297 14415 14331
rect 17693 14297 17727 14331
rect 18797 14297 18831 14331
rect 19441 14297 19475 14331
rect 21281 14297 21315 14331
rect 24685 14297 24719 14331
rect 25421 14297 25455 14331
rect 25513 14297 25547 14331
rect 8493 14229 8527 14263
rect 13645 14229 13679 14263
rect 16221 14229 16255 14263
rect 21649 14229 21683 14263
rect 22753 14229 22787 14263
rect 23305 14229 23339 14263
rect 25881 14229 25915 14263
rect 26801 14229 26835 14263
rect 2421 14025 2455 14059
rect 3065 14025 3099 14059
rect 7757 14025 7791 14059
rect 8309 14025 8343 14059
rect 9413 14025 9447 14059
rect 11069 14025 11103 14059
rect 23213 14025 23247 14059
rect 9229 13957 9263 13991
rect 9565 13957 9599 13991
rect 9781 13957 9815 13991
rect 10793 13957 10827 13991
rect 13185 13957 13219 13991
rect 16865 13957 16899 13991
rect 24685 13957 24719 13991
rect 23309 13923 23343 13957
rect 1409 13889 1443 13923
rect 1685 13889 1719 13923
rect 2605 13889 2639 13923
rect 3157 13889 3191 13923
rect 3801 13889 3835 13923
rect 3985 13889 4019 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 6561 13889 6595 13923
rect 7573 13889 7607 13923
rect 7757 13889 7791 13923
rect 7849 13889 7883 13923
rect 8033 13889 8067 13923
rect 8493 13889 8527 13923
rect 9137 13889 9171 13923
rect 9321 13889 9355 13923
rect 9873 13889 9907 13923
rect 10057 13889 10091 13923
rect 12265 13889 12299 13923
rect 13461 13889 13495 13923
rect 14013 13889 14047 13923
rect 15393 13889 15427 13923
rect 16681 13889 16715 13923
rect 18613 13889 18647 13923
rect 19165 13889 19199 13923
rect 19257 13889 19291 13923
rect 19533 13889 19567 13923
rect 19809 13889 19843 13923
rect 20085 13889 20119 13923
rect 22937 13889 22971 13923
rect 23029 13889 23063 13923
rect 26157 13889 26191 13923
rect 3249 13821 3283 13855
rect 4537 13821 4571 13855
rect 4813 13821 4847 13855
rect 6653 13821 6687 13855
rect 7941 13821 7975 13855
rect 8585 13821 8619 13855
rect 8677 13821 8711 13855
rect 8769 13821 8803 13855
rect 11989 13821 12023 13855
rect 14105 13821 14139 13855
rect 15669 13821 15703 13855
rect 17141 13821 17175 13855
rect 19441 13821 19475 13855
rect 23121 13821 23155 13855
rect 26249 13821 26283 13855
rect 3709 13753 3743 13787
rect 6929 13753 6963 13787
rect 14381 13753 14415 13787
rect 20821 13753 20855 13787
rect 24961 13753 24995 13787
rect 9597 13685 9631 13719
rect 10241 13685 10275 13719
rect 14657 13685 14691 13719
rect 25145 13685 25179 13719
rect 26157 13685 26191 13719
rect 26525 13685 26559 13719
rect 6653 13481 6687 13515
rect 10241 13481 10275 13515
rect 17693 13481 17727 13515
rect 23489 13481 23523 13515
rect 24593 13481 24627 13515
rect 25513 13481 25547 13515
rect 26801 13481 26835 13515
rect 26525 13413 26559 13447
rect 10885 13345 10919 13379
rect 12909 13345 12943 13379
rect 13645 13345 13679 13379
rect 15209 13345 15243 13379
rect 17417 13345 17451 13379
rect 19533 13345 19567 13379
rect 21833 13345 21867 13379
rect 22201 13345 22235 13379
rect 22293 13345 22327 13379
rect 22385 13345 22419 13379
rect 23029 13345 23063 13379
rect 23857 13345 23891 13379
rect 24869 13345 24903 13379
rect 4629 13277 4663 13311
rect 5457 13277 5491 13311
rect 5733 13277 5767 13311
rect 6561 13277 6595 13311
rect 7849 13277 7883 13311
rect 8033 13277 8067 13311
rect 10149 13277 10183 13311
rect 10609 13277 10643 13311
rect 11161 13277 11195 13311
rect 13369 13277 13403 13311
rect 15117 13277 15151 13311
rect 16865 13277 16899 13311
rect 17049 13277 17083 13311
rect 17877 13277 17911 13311
rect 18153 13277 18187 13311
rect 18429 13277 18463 13311
rect 19349 13277 19383 13311
rect 21189 13277 21223 13311
rect 22477 13277 22511 13311
rect 22937 13277 22971 13311
rect 23397 13277 23431 13311
rect 24041 13277 24075 13311
rect 24225 13277 24259 13311
rect 24961 13277 24995 13311
rect 25421 13277 25455 13311
rect 25605 13277 25639 13311
rect 26341 13277 26375 13311
rect 26433 13277 26467 13311
rect 26617 13277 26651 13311
rect 11437 13209 11471 13243
rect 13461 13209 13495 13243
rect 21649 13209 21683 13243
rect 24133 13209 24167 13243
rect 7021 13141 7055 13175
rect 7849 13141 7883 13175
rect 13001 13141 13035 13175
rect 15485 13141 15519 13175
rect 16865 13141 16899 13175
rect 21281 13141 21315 13175
rect 21741 13141 21775 13175
rect 22661 13141 22695 13175
rect 23305 13141 23339 13175
rect 9873 12937 9907 12971
rect 11621 12937 11655 12971
rect 13829 12937 13863 12971
rect 16681 12937 16715 12971
rect 20085 12937 20119 12971
rect 25053 12937 25087 12971
rect 25605 12937 25639 12971
rect 5733 12869 5767 12903
rect 8401 12869 8435 12903
rect 8861 12869 8895 12903
rect 8953 12869 8987 12903
rect 10241 12869 10275 12903
rect 11069 12869 11103 12903
rect 12173 12869 12207 12903
rect 14565 12869 14599 12903
rect 17167 12869 17201 12903
rect 17785 12869 17819 12903
rect 18613 12869 18647 12903
rect 2789 12801 2823 12835
rect 4353 12801 4387 12835
rect 4629 12801 4663 12835
rect 4997 12801 5031 12835
rect 5365 12801 5399 12835
rect 8723 12801 8757 12835
rect 9045 12801 9079 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10057 12801 10091 12835
rect 11345 12801 11379 12835
rect 11805 12801 11839 12835
rect 12081 12801 12115 12835
rect 14289 12801 14323 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 17049 12801 17083 12835
rect 17601 12801 17635 12835
rect 21649 12801 21683 12835
rect 23213 12801 23247 12835
rect 23489 12801 23523 12835
rect 24317 12801 24351 12835
rect 24409 12801 24443 12835
rect 24501 12801 24535 12835
rect 24685 12801 24719 12835
rect 24869 12801 24903 12835
rect 25421 12801 25455 12835
rect 25513 12801 25547 12835
rect 25697 12801 25731 12835
rect 25881 12801 25915 12835
rect 26065 12801 26099 12835
rect 6653 12733 6687 12767
rect 8585 12733 8619 12767
rect 9597 12733 9631 12767
rect 15025 12733 15059 12767
rect 15117 12733 15151 12767
rect 17325 12733 17359 12767
rect 24961 12733 24995 12767
rect 25329 12733 25363 12767
rect 25973 12733 26007 12767
rect 6101 12665 6135 12699
rect 14841 12665 14875 12699
rect 17417 12665 17451 12699
rect 2605 12597 2639 12631
rect 5089 12597 5123 12631
rect 6193 12597 6227 12631
rect 9229 12597 9263 12631
rect 9321 12597 9355 12631
rect 9781 12597 9815 12631
rect 14105 12597 14139 12631
rect 15577 12597 15611 12631
rect 21557 12597 21591 12631
rect 25237 12597 25271 12631
rect 3801 12393 3835 12427
rect 8309 12393 8343 12427
rect 9413 12393 9447 12427
rect 21373 12393 21407 12427
rect 13829 12325 13863 12359
rect 18061 12325 18095 12359
rect 1869 12257 1903 12291
rect 2145 12257 2179 12291
rect 4353 12257 4387 12291
rect 4905 12257 4939 12291
rect 5181 12257 5215 12291
rect 7849 12257 7883 12291
rect 8473 12257 8507 12291
rect 13553 12257 13587 12291
rect 14933 12257 14967 12291
rect 19625 12257 19659 12291
rect 4721 12189 4755 12223
rect 7021 12189 7055 12223
rect 7481 12189 7515 12223
rect 7941 12189 7975 12223
rect 8391 12189 8425 12223
rect 8677 12189 8711 12223
rect 9321 12189 9355 12223
rect 9505 12189 9539 12223
rect 9597 12189 9631 12223
rect 9781 12189 9815 12223
rect 13461 12189 13495 12223
rect 14841 12189 14875 12223
rect 15301 12189 15335 12223
rect 15485 12189 15519 12223
rect 16865 12189 16899 12223
rect 17049 12189 17083 12223
rect 17325 12189 17359 12223
rect 17509 12189 17543 12223
rect 18797 12189 18831 12223
rect 19073 12189 19107 12223
rect 21741 12189 21775 12223
rect 23029 12189 23063 12223
rect 4169 12121 4203 12155
rect 7297 12121 7331 12155
rect 17233 12121 17267 12155
rect 19901 12121 19935 12155
rect 3617 12053 3651 12087
rect 4261 12053 4295 12087
rect 8585 12053 8619 12087
rect 9689 12053 9723 12087
rect 15209 12053 15243 12087
rect 15393 12053 15427 12087
rect 17325 12053 17359 12087
rect 21925 12053 21959 12087
rect 23121 12053 23155 12087
rect 3249 11849 3283 11883
rect 6929 11849 6963 11883
rect 9981 11849 10015 11883
rect 17417 11849 17451 11883
rect 20085 11849 20119 11883
rect 21649 11849 21683 11883
rect 9781 11781 9815 11815
rect 16819 11781 16853 11815
rect 16957 11781 16991 11815
rect 17049 11781 17083 11815
rect 22293 11781 22327 11815
rect 3341 11713 3375 11747
rect 5457 11713 5491 11747
rect 6469 11713 6503 11747
rect 11161 11713 11195 11747
rect 11529 11713 11563 11747
rect 13829 11713 13863 11747
rect 16681 11713 16715 11747
rect 17141 11713 17175 11747
rect 17601 11713 17635 11747
rect 17785 11713 17819 11747
rect 20269 11713 20303 11747
rect 21281 11713 21315 11747
rect 22017 11713 22051 11747
rect 24225 11713 24259 11747
rect 5181 11645 5215 11679
rect 11805 11645 11839 11679
rect 13277 11645 13311 11679
rect 18153 11645 18187 11679
rect 18337 11645 18371 11679
rect 18705 11645 18739 11679
rect 21097 11645 21131 11679
rect 21189 11645 21223 11679
rect 23765 11645 23799 11679
rect 6193 11577 6227 11611
rect 11345 11577 11379 11611
rect 6745 11509 6779 11543
rect 9965 11509 9999 11543
rect 10149 11509 10183 11543
rect 13369 11509 13403 11543
rect 13553 11509 13587 11543
rect 17325 11509 17359 11543
rect 24317 11509 24351 11543
rect 6837 11305 6871 11339
rect 11989 11305 12023 11339
rect 15485 11305 15519 11339
rect 15761 11305 15795 11339
rect 19349 11305 19383 11339
rect 22017 11305 22051 11339
rect 25145 11305 25179 11339
rect 25329 11305 25363 11339
rect 7113 11237 7147 11271
rect 10333 11237 10367 11271
rect 12173 11237 12207 11271
rect 13645 11237 13679 11271
rect 15853 11237 15887 11271
rect 19717 11237 19751 11271
rect 1777 11169 1811 11203
rect 3525 11169 3559 11203
rect 4353 11169 4387 11203
rect 9873 11169 9907 11203
rect 12633 11169 12667 11203
rect 12817 11169 12851 11203
rect 13369 11169 13403 11203
rect 19349 11169 19383 11203
rect 19993 11169 20027 11203
rect 23765 11169 23799 11203
rect 25513 11169 25547 11203
rect 4261 11101 4295 11135
rect 4721 11101 4755 11135
rect 6653 11101 6687 11135
rect 7389 11101 7423 11135
rect 7665 11101 7699 11135
rect 8309 11101 8343 11135
rect 8401 11101 8435 11135
rect 9965 11101 9999 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 10885 11101 10919 11135
rect 11897 11101 11931 11135
rect 15577 11101 15611 11135
rect 17141 11101 17175 11135
rect 17877 11101 17911 11135
rect 18429 11101 18463 11135
rect 18521 11101 18555 11135
rect 18889 11101 18923 11135
rect 19257 11101 19291 11135
rect 19533 11101 19567 11135
rect 22201 11101 22235 11135
rect 22293 11101 22327 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 23857 11101 23891 11135
rect 24501 11101 24535 11135
rect 24649 11101 24683 11135
rect 24777 11101 24811 11135
rect 24966 11101 25000 11135
rect 25605 11101 25639 11135
rect 2053 11033 2087 11067
rect 4169 11033 4203 11067
rect 4905 11033 4939 11067
rect 6561 11033 6595 11067
rect 8677 11033 8711 11067
rect 10425 11033 10459 11067
rect 12541 11033 12575 11067
rect 16221 11033 16255 11067
rect 16957 11033 16991 11067
rect 17325 11033 17359 11067
rect 18153 11033 18187 11067
rect 20177 11033 20211 11067
rect 21833 11033 21867 11067
rect 22523 11033 22557 11067
rect 24869 11033 24903 11067
rect 3801 10965 3835 10999
rect 13829 10965 13863 10999
rect 15117 10965 15151 10999
rect 24225 10965 24259 10999
rect 2697 10761 2731 10795
rect 3249 10761 3283 10795
rect 7757 10761 7791 10795
rect 8033 10761 8067 10795
rect 15301 10761 15335 10795
rect 21373 10761 21407 10795
rect 22385 10761 22419 10795
rect 24593 10761 24627 10795
rect 25237 10761 25271 10795
rect 8677 10693 8711 10727
rect 10333 10693 10367 10727
rect 13645 10693 13679 10727
rect 14105 10693 14139 10727
rect 22293 10693 22327 10727
rect 2881 10625 2915 10659
rect 3341 10625 3375 10659
rect 4077 10625 4111 10659
rect 4445 10625 4479 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5457 10625 5491 10659
rect 6653 10625 6687 10659
rect 7665 10625 7699 10659
rect 7941 10625 7975 10659
rect 8217 10625 8251 10659
rect 8309 10625 8343 10659
rect 8493 10625 8527 10659
rect 8585 10625 8619 10659
rect 8861 10625 8895 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 9597 10625 9631 10659
rect 10149 10625 10183 10659
rect 10241 10625 10275 10659
rect 12817 10625 12851 10659
rect 13461 10625 13495 10659
rect 13553 10625 13587 10659
rect 13921 10625 13955 10659
rect 14289 10625 14323 10659
rect 14381 10625 14415 10659
rect 14565 10625 14599 10659
rect 14657 10625 14691 10659
rect 14841 10625 14875 10659
rect 16313 10625 16347 10659
rect 17325 10625 17359 10659
rect 17693 10625 17727 10659
rect 17877 10625 17911 10659
rect 19073 10625 19107 10659
rect 19441 10625 19475 10659
rect 19717 10625 19751 10659
rect 20085 10625 20119 10659
rect 20637 10625 20671 10659
rect 22017 10625 22051 10659
rect 22385 10625 22419 10659
rect 22845 10625 22879 10659
rect 24133 10625 24167 10659
rect 24225 10625 24259 10659
rect 24409 10625 24443 10659
rect 25421 10625 25455 10659
rect 4905 10557 4939 10591
rect 5181 10557 5215 10591
rect 6745 10557 6779 10591
rect 7481 10557 7515 10591
rect 9045 10557 9079 10591
rect 9873 10557 9907 10591
rect 12909 10557 12943 10591
rect 14933 10557 14967 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 19901 10557 19935 10591
rect 20361 10557 20395 10591
rect 22201 10557 22235 10591
rect 22707 10557 22741 10591
rect 25605 10557 25639 10591
rect 6193 10489 6227 10523
rect 9689 10489 9723 10523
rect 13829 10489 13863 10523
rect 15853 10489 15887 10523
rect 17785 10489 17819 10523
rect 7941 10421 7975 10455
rect 9965 10421 9999 10455
rect 10057 10421 10091 10455
rect 13185 10421 13219 10455
rect 16037 10421 16071 10455
rect 17509 10421 17543 10455
rect 21833 10421 21867 10455
rect 22293 10421 22327 10455
rect 22569 10421 22603 10455
rect 13461 10217 13495 10251
rect 13645 10217 13679 10251
rect 14289 10217 14323 10251
rect 14657 10217 14691 10251
rect 17233 10217 17267 10251
rect 24961 10217 24995 10251
rect 25973 10217 26007 10251
rect 14473 10149 14507 10183
rect 20913 10149 20947 10183
rect 24777 10149 24811 10183
rect 10149 10081 10183 10115
rect 14749 10081 14783 10115
rect 15025 10081 15059 10115
rect 15485 10081 15519 10115
rect 16681 10081 16715 10115
rect 17325 10081 17359 10115
rect 19625 10081 19659 10115
rect 20177 10081 20211 10115
rect 21465 10081 21499 10115
rect 6469 10013 6503 10047
rect 6745 10013 6779 10047
rect 8953 10013 8987 10047
rect 9137 10013 9171 10047
rect 10241 10013 10275 10047
rect 12541 10013 12575 10047
rect 12633 10013 12667 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 13185 10013 13219 10047
rect 14197 10013 14231 10047
rect 14841 10013 14875 10047
rect 14933 10013 14967 10047
rect 15117 10013 15151 10047
rect 15577 10013 15611 10047
rect 19441 10013 19475 10047
rect 19717 10013 19751 10047
rect 20453 10013 20487 10047
rect 20636 10013 20670 10047
rect 21281 10013 21315 10047
rect 21373 10013 21407 10047
rect 21557 10013 21591 10047
rect 22569 10013 22603 10047
rect 22753 10013 22787 10047
rect 25697 10013 25731 10047
rect 25973 10013 26007 10047
rect 9045 9945 9079 9979
rect 17601 9945 17635 9979
rect 19349 9945 19383 9979
rect 20315 9945 20349 9979
rect 20545 9945 20579 9979
rect 21097 9945 21131 9979
rect 24501 9945 24535 9979
rect 25881 9945 25915 9979
rect 7481 9877 7515 9911
rect 10609 9877 10643 9911
rect 13001 9877 13035 9911
rect 15945 9877 15979 9911
rect 16773 9877 16807 9911
rect 16865 9877 16899 9911
rect 19073 9877 19107 9911
rect 20085 9877 20119 9911
rect 20821 9877 20855 9911
rect 22661 9877 22695 9911
rect 8769 9673 8803 9707
rect 12633 9673 12667 9707
rect 16957 9673 16991 9707
rect 5917 9605 5951 9639
rect 6561 9605 6595 9639
rect 8217 9605 8251 9639
rect 17443 9605 17477 9639
rect 22477 9605 22511 9639
rect 22845 9605 22879 9639
rect 23857 9605 23891 9639
rect 23949 9605 23983 9639
rect 4537 9537 4571 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 9682 9537 9716 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11529 9537 11563 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12541 9537 12575 9571
rect 12817 9537 12851 9571
rect 13185 9537 13219 9571
rect 13369 9537 13403 9571
rect 17141 9537 17175 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 22339 9537 22373 9571
rect 22569 9537 22603 9571
rect 22661 9537 22695 9571
rect 23121 9537 23155 9571
rect 23719 9537 23753 9571
rect 24041 9537 24075 9571
rect 24869 9537 24903 9571
rect 25053 9537 25087 9571
rect 25145 9537 25179 9571
rect 25329 9537 25363 9571
rect 25421 9537 25455 9571
rect 26065 9537 26099 9571
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 4077 9469 4111 9503
rect 4629 9469 4663 9503
rect 4813 9469 4847 9503
rect 6193 9469 6227 9503
rect 6377 9469 6411 9503
rect 8309 9469 8343 9503
rect 8861 9469 8895 9503
rect 9597 9469 9631 9503
rect 9965 9469 9999 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 10241 9469 10275 9503
rect 10701 9469 10735 9503
rect 13093 9469 13127 9503
rect 17601 9469 17635 9503
rect 22201 9469 22235 9503
rect 23029 9469 23063 9503
rect 23489 9469 23523 9503
rect 23581 9469 23615 9503
rect 26157 9469 26191 9503
rect 8585 9401 8619 9435
rect 8953 9401 8987 9435
rect 12265 9401 12299 9435
rect 25697 9401 25731 9435
rect 4169 9333 4203 9367
rect 9781 9333 9815 9367
rect 13001 9333 13035 9367
rect 13185 9333 13219 9367
rect 24225 9333 24259 9367
rect 2881 9129 2915 9163
rect 3433 9129 3467 9163
rect 9781 9129 9815 9163
rect 12633 9129 12667 9163
rect 14565 9129 14599 9163
rect 14749 9129 14783 9163
rect 22937 9129 22971 9163
rect 25329 9129 25363 9163
rect 26249 9129 26283 9163
rect 13277 9061 13311 9095
rect 25421 9061 25455 9095
rect 5549 8993 5583 9027
rect 7941 8993 7975 9027
rect 13001 8993 13035 9027
rect 20913 8993 20947 9027
rect 21833 8993 21867 9027
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 4629 8925 4663 8959
rect 4813 8925 4847 8959
rect 4997 8925 5031 8959
rect 6929 8925 6963 8959
rect 7205 8925 7239 8959
rect 7389 8925 7423 8959
rect 9413 8925 9447 8959
rect 12455 8925 12489 8959
rect 12633 8925 12667 8959
rect 12909 8925 12943 8959
rect 14289 8925 14323 8959
rect 15209 8925 15243 8959
rect 17969 8925 18003 8959
rect 18245 8925 18279 8959
rect 21741 8925 21775 8959
rect 22569 8925 22603 8959
rect 25789 8925 25823 8959
rect 25973 8925 26007 8959
rect 26065 8925 26099 8959
rect 26341 8925 26375 8959
rect 5273 8857 5307 8891
rect 7665 8857 7699 8891
rect 9597 8857 9631 8891
rect 22753 8857 22787 8891
rect 15393 8789 15427 8823
rect 17233 8789 17267 8823
rect 26433 8789 26467 8823
rect 10333 8585 10367 8619
rect 12541 8585 12575 8619
rect 13553 8585 13587 8619
rect 14933 8585 14967 8619
rect 15301 8585 15335 8619
rect 22293 8585 22327 8619
rect 23397 8585 23431 8619
rect 24593 8585 24627 8619
rect 24961 8585 24995 8619
rect 25881 8585 25915 8619
rect 8447 8517 8481 8551
rect 16247 8517 16281 8551
rect 17325 8517 17359 8551
rect 25237 8517 25271 8551
rect 25329 8517 25363 8551
rect 25697 8517 25731 8551
rect 26157 8517 26191 8551
rect 6653 8449 6687 8483
rect 7665 8449 7699 8483
rect 7849 8449 7883 8483
rect 8125 8449 8159 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 8685 8449 8719 8483
rect 8861 8449 8895 8483
rect 9137 8449 9171 8483
rect 9413 8449 9447 8483
rect 10241 8449 10275 8483
rect 10425 8449 10459 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 12449 8449 12483 8483
rect 12633 8449 12667 8483
rect 14381 8449 14415 8483
rect 15393 8449 15427 8483
rect 15761 8449 15795 8483
rect 15945 8449 15979 8483
rect 16037 8449 16071 8483
rect 16129 8449 16163 8483
rect 16405 8449 16439 8483
rect 16865 8449 16899 8483
rect 19717 8449 19751 8483
rect 21833 8449 21867 8483
rect 22661 8449 22695 8483
rect 23673 8449 23707 8483
rect 25145 8449 25179 8483
rect 25513 8449 25547 8483
rect 25605 8449 25639 8483
rect 25973 8449 26007 8483
rect 26065 8449 26099 8483
rect 7757 8381 7791 8415
rect 8585 8381 8619 8415
rect 9321 8381 9355 8415
rect 14473 8381 14507 8415
rect 15577 8381 15611 8415
rect 17141 8381 17175 8415
rect 18153 8381 18187 8415
rect 19901 8381 19935 8415
rect 20821 8381 20855 8415
rect 22385 8381 22419 8415
rect 23581 8381 23615 8415
rect 24133 8381 24167 8415
rect 7941 8313 7975 8347
rect 8769 8313 8803 8347
rect 10517 8313 10551 8347
rect 24041 8313 24075 8347
rect 24501 8313 24535 8347
rect 25697 8313 25731 8347
rect 6929 8245 6963 8279
rect 7113 8245 7147 8279
rect 8953 8245 8987 8279
rect 9137 8245 9171 8279
rect 16773 8245 16807 8279
rect 22017 8245 22051 8279
rect 7205 8041 7239 8075
rect 7757 8041 7791 8075
rect 8953 8041 8987 8075
rect 10885 8041 10919 8075
rect 11253 8041 11287 8075
rect 17141 8041 17175 8075
rect 17969 8041 18003 8075
rect 19717 8041 19751 8075
rect 21373 8041 21407 8075
rect 25881 8041 25915 8075
rect 10793 7973 10827 8007
rect 25697 7973 25731 8007
rect 4997 7905 5031 7939
rect 5365 7905 5399 7939
rect 5641 7905 5675 7939
rect 7573 7905 7607 7939
rect 10517 7905 10551 7939
rect 10701 7905 10735 7939
rect 13277 7905 13311 7939
rect 15393 7905 15427 7939
rect 17693 7905 17727 7939
rect 19257 7905 19291 7939
rect 20361 7905 20395 7939
rect 22569 7905 22603 7939
rect 3985 7837 4019 7871
rect 4077 7837 4111 7871
rect 5181 7837 5215 7871
rect 7113 7837 7147 7871
rect 7665 7837 7699 7871
rect 7849 7837 7883 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 10425 7837 10459 7871
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 11253 7837 11287 7871
rect 13461 7837 13495 7871
rect 18245 7837 18279 7871
rect 18429 7837 18463 7871
rect 18705 7837 18739 7871
rect 19625 7837 19659 7871
rect 19993 7837 20027 7871
rect 20177 7837 20211 7871
rect 20637 7837 20671 7871
rect 23949 7837 23983 7871
rect 4721 7769 4755 7803
rect 9137 7769 9171 7803
rect 9321 7769 9355 7803
rect 11621 7769 11655 7803
rect 15669 7769 15703 7803
rect 23765 7769 23799 7803
rect 25421 7769 25455 7803
rect 3801 7701 3835 7735
rect 4169 7701 4203 7735
rect 4353 7701 4387 7735
rect 4813 7701 4847 7735
rect 9413 7701 9447 7735
rect 10057 7701 10091 7735
rect 5181 7497 5215 7531
rect 7389 7497 7423 7531
rect 15945 7497 15979 7531
rect 20545 7497 20579 7531
rect 20637 7497 20671 7531
rect 23213 7497 23247 7531
rect 25053 7497 25087 7531
rect 25605 7497 25639 7531
rect 3709 7429 3743 7463
rect 8677 7429 8711 7463
rect 8815 7429 8849 7463
rect 13277 7429 13311 7463
rect 23305 7429 23339 7463
rect 6653 7361 6687 7395
rect 8493 7361 8527 7395
rect 8585 7361 8619 7395
rect 8953 7361 8987 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 13093 7361 13127 7395
rect 13185 7361 13219 7395
rect 13395 7361 13429 7395
rect 13829 7361 13863 7395
rect 14013 7361 14047 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 15393 7361 15427 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 16037 7361 16071 7395
rect 18061 7361 18095 7395
rect 18245 7361 18279 7395
rect 18521 7361 18555 7395
rect 19073 7361 19107 7395
rect 19441 7361 19475 7395
rect 19717 7361 19751 7395
rect 19993 7361 20027 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 24593 7361 24627 7395
rect 25145 7361 25179 7395
rect 3433 7293 3467 7327
rect 6377 7293 6411 7327
rect 13553 7293 13587 7327
rect 14289 7293 14323 7327
rect 17509 7293 17543 7327
rect 19901 7293 19935 7327
rect 20821 7293 20855 7327
rect 23029 7293 23063 7327
rect 22845 7225 22879 7259
rect 24961 7225 24995 7259
rect 8309 7157 8343 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 13645 7157 13679 7191
rect 14381 7157 14415 7191
rect 14565 7157 14599 7191
rect 15761 7157 15795 7191
rect 17969 7157 18003 7191
rect 20177 7157 20211 7191
rect 23673 7157 23707 7191
rect 25237 7157 25271 7191
rect 9137 6953 9171 6987
rect 10517 6953 10551 6987
rect 13093 6953 13127 6987
rect 13277 6953 13311 6987
rect 7665 6817 7699 6851
rect 9505 6817 9539 6851
rect 9873 6817 9907 6851
rect 12081 6817 12115 6851
rect 14473 6817 14507 6851
rect 14749 6817 14783 6851
rect 15853 6817 15887 6851
rect 17417 6817 17451 6851
rect 18061 6817 18095 6851
rect 19257 6817 19291 6851
rect 20085 6817 20119 6851
rect 21373 6817 21407 6851
rect 22385 6817 22419 6851
rect 23213 6817 23247 6851
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 7481 6749 7515 6783
rect 9045 6749 9079 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 11989 6749 12023 6783
rect 13001 6749 13035 6783
rect 13185 6749 13219 6783
rect 13456 6749 13490 6783
rect 13773 6749 13807 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 14841 6749 14875 6783
rect 14933 6749 14967 6783
rect 15091 6749 15125 6783
rect 15301 6749 15335 6783
rect 15393 6749 15427 6783
rect 15577 6749 15611 6783
rect 15945 6749 15979 6783
rect 17233 6749 17267 6783
rect 19625 6749 19659 6783
rect 19993 6749 20027 6783
rect 20177 6749 20211 6783
rect 22569 6749 22603 6783
rect 23121 6749 23155 6783
rect 23489 6749 23523 6783
rect 13553 6681 13587 6715
rect 13645 6681 13679 6715
rect 15209 6681 15243 6715
rect 16037 6681 16071 6715
rect 6285 6613 6319 6647
rect 6745 6613 6779 6647
rect 7021 6613 7055 6647
rect 7389 6613 7423 6647
rect 10149 6613 10183 6647
rect 10241 6613 10275 6647
rect 11529 6613 11563 6647
rect 11897 6613 11931 6647
rect 16405 6613 16439 6647
rect 22661 6613 22695 6647
rect 23029 6613 23063 6647
rect 23673 6613 23707 6647
rect 9413 6409 9447 6443
rect 15577 6409 15611 6443
rect 25421 6409 25455 6443
rect 23949 6341 23983 6375
rect 10149 6273 10183 6307
rect 10517 6273 10551 6307
rect 10701 6273 10735 6307
rect 11253 6273 11287 6307
rect 11713 6273 11747 6307
rect 15485 6273 15519 6307
rect 15669 6273 15703 6307
rect 16037 6273 16071 6307
rect 18061 6273 18095 6307
rect 18337 6273 18371 6307
rect 19165 6273 19199 6307
rect 21373 6273 21407 6307
rect 21833 6273 21867 6307
rect 23673 6273 23707 6307
rect 7481 6205 7515 6239
rect 7665 6205 7699 6239
rect 8401 6205 8435 6239
rect 10425 6205 10459 6239
rect 10885 6205 10919 6239
rect 19441 6205 19475 6239
rect 22109 6205 22143 6239
rect 11253 6137 11287 6171
rect 17325 6137 17359 6171
rect 20913 6137 20947 6171
rect 21557 6137 21591 6171
rect 23581 6137 23615 6171
rect 11529 6069 11563 6103
rect 16221 6069 16255 6103
rect 5996 5865 6030 5899
rect 7481 5865 7515 5899
rect 9321 5865 9355 5899
rect 9505 5865 9539 5899
rect 12817 5865 12851 5899
rect 13829 5865 13863 5899
rect 17785 5865 17819 5899
rect 19441 5865 19475 5899
rect 20269 5865 20303 5899
rect 22477 5865 22511 5899
rect 23581 5865 23615 5899
rect 13645 5797 13679 5831
rect 5733 5729 5767 5763
rect 10517 5729 10551 5763
rect 10793 5729 10827 5763
rect 12633 5729 12667 5763
rect 15301 5729 15335 5763
rect 16037 5729 16071 5763
rect 16313 5729 16347 5763
rect 9045 5661 9079 5695
rect 12541 5661 12575 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 14565 5661 14599 5695
rect 15209 5661 15243 5695
rect 18153 5661 18187 5695
rect 19625 5661 19659 5695
rect 20177 5661 20211 5695
rect 22385 5661 22419 5695
rect 23489 5661 23523 5695
rect 13369 5593 13403 5627
rect 18061 5593 18095 5627
rect 12265 5525 12299 5559
rect 14749 5525 14783 5559
rect 14841 5525 14875 5559
rect 11621 5321 11655 5355
rect 12633 5321 12667 5355
rect 13001 5321 13035 5355
rect 14289 5321 14323 5355
rect 15209 5321 15243 5355
rect 13829 5253 13863 5287
rect 11529 5185 11563 5219
rect 12265 5185 12299 5219
rect 13185 5185 13219 5219
rect 13369 5185 13403 5219
rect 14841 5185 14875 5219
rect 12357 5117 12391 5151
rect 14749 5117 14783 5151
rect 14105 5049 14139 5083
<< metal1 >>
rect 1104 29402 30820 29424
rect 1104 29350 5324 29402
rect 5376 29350 5388 29402
rect 5440 29350 5452 29402
rect 5504 29350 5516 29402
rect 5568 29350 5580 29402
rect 5632 29350 12752 29402
rect 12804 29350 12816 29402
rect 12868 29350 12880 29402
rect 12932 29350 12944 29402
rect 12996 29350 13008 29402
rect 13060 29350 20180 29402
rect 20232 29350 20244 29402
rect 20296 29350 20308 29402
rect 20360 29350 20372 29402
rect 20424 29350 20436 29402
rect 20488 29350 27608 29402
rect 27660 29350 27672 29402
rect 27724 29350 27736 29402
rect 27788 29350 27800 29402
rect 27852 29350 27864 29402
rect 27916 29350 30820 29402
rect 1104 29328 30820 29350
rect 13078 29248 13084 29300
rect 13136 29288 13142 29300
rect 13173 29291 13231 29297
rect 13173 29288 13185 29291
rect 13136 29260 13185 29288
rect 13136 29248 13142 29260
rect 13173 29257 13185 29260
rect 13219 29257 13231 29291
rect 13173 29251 13231 29257
rect 15470 29248 15476 29300
rect 15528 29288 15534 29300
rect 15657 29291 15715 29297
rect 15657 29288 15669 29291
rect 15528 29260 15669 29288
rect 15528 29248 15534 29260
rect 15657 29257 15669 29260
rect 15703 29257 15715 29291
rect 15657 29251 15715 29257
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18233 29291 18291 29297
rect 18233 29288 18245 29291
rect 18196 29260 18245 29288
rect 18196 29248 18202 29260
rect 18233 29257 18245 29260
rect 18279 29257 18291 29291
rect 18233 29251 18291 29257
rect 13081 29155 13139 29161
rect 13081 29121 13093 29155
rect 13127 29152 13139 29155
rect 13354 29152 13360 29164
rect 13127 29124 13360 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13354 29112 13360 29124
rect 13412 29112 13418 29164
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29152 15991 29155
rect 16390 29152 16396 29164
rect 15979 29124 16396 29152
rect 15979 29121 15991 29124
rect 15933 29115 15991 29121
rect 16390 29112 16396 29124
rect 16448 29112 16454 29164
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 18509 29155 18567 29161
rect 18509 29152 18521 29155
rect 18104 29124 18521 29152
rect 18104 29112 18110 29124
rect 18509 29121 18521 29124
rect 18555 29121 18567 29155
rect 18509 29115 18567 29121
rect 1104 28858 30820 28880
rect 1104 28806 4664 28858
rect 4716 28806 4728 28858
rect 4780 28806 4792 28858
rect 4844 28806 4856 28858
rect 4908 28806 4920 28858
rect 4972 28806 12092 28858
rect 12144 28806 12156 28858
rect 12208 28806 12220 28858
rect 12272 28806 12284 28858
rect 12336 28806 12348 28858
rect 12400 28806 19520 28858
rect 19572 28806 19584 28858
rect 19636 28806 19648 28858
rect 19700 28806 19712 28858
rect 19764 28806 19776 28858
rect 19828 28806 26948 28858
rect 27000 28806 27012 28858
rect 27064 28806 27076 28858
rect 27128 28806 27140 28858
rect 27192 28806 27204 28858
rect 27256 28806 30820 28858
rect 1104 28784 30820 28806
rect 1104 28314 30820 28336
rect 1104 28262 5324 28314
rect 5376 28262 5388 28314
rect 5440 28262 5452 28314
rect 5504 28262 5516 28314
rect 5568 28262 5580 28314
rect 5632 28262 12752 28314
rect 12804 28262 12816 28314
rect 12868 28262 12880 28314
rect 12932 28262 12944 28314
rect 12996 28262 13008 28314
rect 13060 28262 20180 28314
rect 20232 28262 20244 28314
rect 20296 28262 20308 28314
rect 20360 28262 20372 28314
rect 20424 28262 20436 28314
rect 20488 28262 27608 28314
rect 27660 28262 27672 28314
rect 27724 28262 27736 28314
rect 27788 28262 27800 28314
rect 27852 28262 27864 28314
rect 27916 28262 30820 28314
rect 1104 28240 30820 28262
rect 1104 27770 30820 27792
rect 1104 27718 4664 27770
rect 4716 27718 4728 27770
rect 4780 27718 4792 27770
rect 4844 27718 4856 27770
rect 4908 27718 4920 27770
rect 4972 27718 12092 27770
rect 12144 27718 12156 27770
rect 12208 27718 12220 27770
rect 12272 27718 12284 27770
rect 12336 27718 12348 27770
rect 12400 27718 19520 27770
rect 19572 27718 19584 27770
rect 19636 27718 19648 27770
rect 19700 27718 19712 27770
rect 19764 27718 19776 27770
rect 19828 27718 26948 27770
rect 27000 27718 27012 27770
rect 27064 27718 27076 27770
rect 27128 27718 27140 27770
rect 27192 27718 27204 27770
rect 27256 27718 30820 27770
rect 1104 27696 30820 27718
rect 1104 27226 30820 27248
rect 1104 27174 5324 27226
rect 5376 27174 5388 27226
rect 5440 27174 5452 27226
rect 5504 27174 5516 27226
rect 5568 27174 5580 27226
rect 5632 27174 12752 27226
rect 12804 27174 12816 27226
rect 12868 27174 12880 27226
rect 12932 27174 12944 27226
rect 12996 27174 13008 27226
rect 13060 27174 20180 27226
rect 20232 27174 20244 27226
rect 20296 27174 20308 27226
rect 20360 27174 20372 27226
rect 20424 27174 20436 27226
rect 20488 27174 27608 27226
rect 27660 27174 27672 27226
rect 27724 27174 27736 27226
rect 27788 27174 27800 27226
rect 27852 27174 27864 27226
rect 27916 27174 30820 27226
rect 1104 27152 30820 27174
rect 14550 26936 14556 26988
rect 14608 26936 14614 26988
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26976 14795 26979
rect 15194 26976 15200 26988
rect 14783 26948 15200 26976
rect 14783 26945 14795 26948
rect 14737 26939 14795 26945
rect 15194 26936 15200 26948
rect 15252 26936 15258 26988
rect 15470 26936 15476 26988
rect 15528 26936 15534 26988
rect 16945 26979 17003 26985
rect 16945 26945 16957 26979
rect 16991 26945 17003 26979
rect 16945 26939 17003 26945
rect 16960 26908 16988 26939
rect 17497 26911 17555 26917
rect 17497 26908 17509 26911
rect 16960 26880 17509 26908
rect 17497 26877 17509 26880
rect 17543 26877 17555 26911
rect 17497 26871 17555 26877
rect 17957 26911 18015 26917
rect 17957 26877 17969 26911
rect 18003 26908 18015 26911
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 18003 26880 18061 26908
rect 18003 26877 18015 26880
rect 17957 26871 18015 26877
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 18690 26868 18696 26920
rect 18748 26868 18754 26920
rect 17681 26843 17739 26849
rect 17681 26809 17693 26843
rect 17727 26840 17739 26843
rect 19886 26840 19892 26852
rect 17727 26812 19892 26840
rect 17727 26809 17739 26812
rect 17681 26803 17739 26809
rect 19886 26800 19892 26812
rect 19944 26800 19950 26852
rect 14642 26732 14648 26784
rect 14700 26732 14706 26784
rect 15289 26775 15347 26781
rect 15289 26741 15301 26775
rect 15335 26772 15347 26775
rect 15378 26772 15384 26784
rect 15335 26744 15384 26772
rect 15335 26741 15347 26744
rect 15289 26735 15347 26741
rect 15378 26732 15384 26744
rect 15436 26732 15442 26784
rect 17126 26732 17132 26784
rect 17184 26732 17190 26784
rect 1104 26682 30820 26704
rect 1104 26630 4664 26682
rect 4716 26630 4728 26682
rect 4780 26630 4792 26682
rect 4844 26630 4856 26682
rect 4908 26630 4920 26682
rect 4972 26630 12092 26682
rect 12144 26630 12156 26682
rect 12208 26630 12220 26682
rect 12272 26630 12284 26682
rect 12336 26630 12348 26682
rect 12400 26630 19520 26682
rect 19572 26630 19584 26682
rect 19636 26630 19648 26682
rect 19700 26630 19712 26682
rect 19764 26630 19776 26682
rect 19828 26630 26948 26682
rect 27000 26630 27012 26682
rect 27064 26630 27076 26682
rect 27128 26630 27140 26682
rect 27192 26630 27204 26682
rect 27256 26630 30820 26682
rect 1104 26608 30820 26630
rect 17126 26528 17132 26580
rect 17184 26528 17190 26580
rect 19886 26528 19892 26580
rect 19944 26528 19950 26580
rect 15381 26435 15439 26441
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 16301 26435 16359 26441
rect 16301 26432 16313 26435
rect 15427 26404 16313 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 16301 26401 16313 26404
rect 16347 26401 16359 26435
rect 17144 26432 17172 26528
rect 18601 26503 18659 26509
rect 18601 26469 18613 26503
rect 18647 26469 18659 26503
rect 18601 26463 18659 26469
rect 18616 26432 18644 26463
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 17144 26404 17356 26432
rect 18616 26404 19257 26432
rect 16301 26395 16359 26401
rect 14090 26324 14096 26376
rect 14148 26324 14154 26376
rect 14366 26324 14372 26376
rect 14424 26364 14430 26376
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14424 26336 15025 26364
rect 14424 26324 14430 26336
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15289 26367 15347 26373
rect 15289 26364 15301 26367
rect 15013 26327 15071 26333
rect 15212 26336 15301 26364
rect 14734 26256 14740 26308
rect 14792 26296 14798 26308
rect 14829 26299 14887 26305
rect 14829 26296 14841 26299
rect 14792 26268 14841 26296
rect 14792 26256 14798 26268
rect 14829 26265 14841 26268
rect 14875 26265 14887 26299
rect 14829 26259 14887 26265
rect 15212 26240 15240 26336
rect 15289 26333 15301 26336
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26364 15531 26367
rect 15519 26336 15608 26364
rect 15519 26333 15531 26336
rect 15473 26327 15531 26333
rect 15580 26240 15608 26336
rect 16206 26324 16212 26376
rect 16264 26324 16270 26376
rect 16758 26324 16764 26376
rect 16816 26364 16822 26376
rect 17221 26367 17279 26373
rect 17221 26364 17233 26367
rect 16816 26336 17233 26364
rect 16816 26324 16822 26336
rect 17221 26333 17233 26336
rect 17267 26333 17279 26367
rect 17328 26364 17356 26404
rect 19245 26401 19257 26404
rect 19291 26401 19303 26435
rect 19245 26395 19303 26401
rect 17477 26367 17535 26373
rect 17477 26364 17489 26367
rect 17328 26336 17489 26364
rect 17221 26327 17279 26333
rect 17477 26333 17489 26336
rect 17523 26333 17535 26367
rect 17477 26327 17535 26333
rect 15194 26188 15200 26240
rect 15252 26188 15258 26240
rect 15562 26188 15568 26240
rect 15620 26188 15626 26240
rect 16942 26188 16948 26240
rect 17000 26188 17006 26240
rect 1104 26138 30820 26160
rect 1104 26086 5324 26138
rect 5376 26086 5388 26138
rect 5440 26086 5452 26138
rect 5504 26086 5516 26138
rect 5568 26086 5580 26138
rect 5632 26086 12752 26138
rect 12804 26086 12816 26138
rect 12868 26086 12880 26138
rect 12932 26086 12944 26138
rect 12996 26086 13008 26138
rect 13060 26086 20180 26138
rect 20232 26086 20244 26138
rect 20296 26086 20308 26138
rect 20360 26086 20372 26138
rect 20424 26086 20436 26138
rect 20488 26086 27608 26138
rect 27660 26086 27672 26138
rect 27724 26086 27736 26138
rect 27788 26086 27800 26138
rect 27852 26086 27864 26138
rect 27916 26086 30820 26138
rect 1104 26064 30820 26086
rect 13081 26027 13139 26033
rect 13081 25993 13093 26027
rect 13127 26024 13139 26027
rect 14090 26024 14096 26036
rect 13127 25996 14096 26024
rect 13127 25993 13139 25996
rect 13081 25987 13139 25993
rect 14090 25984 14096 25996
rect 14148 25984 14154 26036
rect 14550 25984 14556 26036
rect 14608 25984 14614 26036
rect 14734 25984 14740 26036
rect 14792 25984 14798 26036
rect 16206 25984 16212 26036
rect 16264 25984 16270 26036
rect 18049 26027 18107 26033
rect 18049 25993 18061 26027
rect 18095 26024 18107 26027
rect 18690 26024 18696 26036
rect 18095 25996 18696 26024
rect 18095 25993 18107 25996
rect 18049 25987 18107 25993
rect 18690 25984 18696 25996
rect 18748 26024 18754 26036
rect 18748 25996 19748 26024
rect 18748 25984 18754 25996
rect 14216 25959 14274 25965
rect 14216 25925 14228 25959
rect 14262 25956 14274 25959
rect 14642 25956 14648 25968
rect 14262 25928 14648 25956
rect 14262 25925 14274 25928
rect 14216 25919 14274 25925
rect 14642 25916 14648 25928
rect 14700 25916 14706 25968
rect 11876 25891 11934 25897
rect 11876 25857 11888 25891
rect 11922 25888 11934 25891
rect 12802 25888 12808 25900
rect 11922 25860 12808 25888
rect 11922 25857 11934 25860
rect 11876 25851 11934 25857
rect 12802 25848 12808 25860
rect 12860 25848 12866 25900
rect 14366 25848 14372 25900
rect 14424 25888 14430 25900
rect 14752 25897 14780 25984
rect 16942 25965 16948 25968
rect 16936 25956 16948 25965
rect 14844 25928 16712 25956
rect 16903 25928 16948 25956
rect 14844 25897 14872 25928
rect 14553 25891 14611 25897
rect 14553 25888 14565 25891
rect 14424 25860 14565 25888
rect 14424 25848 14430 25860
rect 14553 25857 14565 25860
rect 14599 25857 14611 25891
rect 14553 25851 14611 25857
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 14829 25891 14887 25897
rect 14829 25857 14841 25891
rect 14875 25857 14887 25891
rect 14829 25851 14887 25857
rect 15096 25891 15154 25897
rect 15096 25857 15108 25891
rect 15142 25888 15154 25891
rect 15378 25888 15384 25900
rect 15142 25860 15384 25888
rect 15142 25857 15154 25860
rect 15096 25851 15154 25857
rect 10870 25780 10876 25832
rect 10928 25820 10934 25832
rect 11609 25823 11667 25829
rect 11609 25820 11621 25823
rect 10928 25792 11621 25820
rect 10928 25780 10934 25792
rect 11609 25789 11621 25792
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 14461 25823 14519 25829
rect 14461 25789 14473 25823
rect 14507 25820 14519 25823
rect 14844 25820 14872 25851
rect 15378 25848 15384 25860
rect 15436 25848 15442 25900
rect 16684 25897 16712 25928
rect 16936 25919 16948 25928
rect 16942 25916 16948 25919
rect 17000 25916 17006 25968
rect 16669 25891 16727 25897
rect 16669 25857 16681 25891
rect 16715 25888 16727 25891
rect 16758 25888 16764 25900
rect 16715 25860 16764 25888
rect 16715 25857 16727 25860
rect 16669 25851 16727 25857
rect 16758 25848 16764 25860
rect 16816 25848 16822 25900
rect 19720 25897 19748 25996
rect 19705 25891 19763 25897
rect 19705 25857 19717 25891
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 14507 25792 14872 25820
rect 19153 25823 19211 25829
rect 14507 25789 14519 25792
rect 14461 25783 14519 25789
rect 19153 25789 19165 25823
rect 19199 25820 19211 25823
rect 19245 25823 19303 25829
rect 19245 25820 19257 25823
rect 19199 25792 19257 25820
rect 19199 25789 19211 25792
rect 19153 25783 19211 25789
rect 19245 25789 19257 25792
rect 19291 25789 19303 25823
rect 19245 25783 19303 25789
rect 12986 25644 12992 25696
rect 13044 25644 13050 25696
rect 18506 25644 18512 25696
rect 18564 25644 18570 25696
rect 19613 25687 19671 25693
rect 19613 25653 19625 25687
rect 19659 25684 19671 25687
rect 19886 25684 19892 25696
rect 19659 25656 19892 25684
rect 19659 25653 19671 25656
rect 19613 25647 19671 25653
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 1104 25594 30820 25616
rect 1104 25542 4664 25594
rect 4716 25542 4728 25594
rect 4780 25542 4792 25594
rect 4844 25542 4856 25594
rect 4908 25542 4920 25594
rect 4972 25542 12092 25594
rect 12144 25542 12156 25594
rect 12208 25542 12220 25594
rect 12272 25542 12284 25594
rect 12336 25542 12348 25594
rect 12400 25542 19520 25594
rect 19572 25542 19584 25594
rect 19636 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 26948 25594
rect 27000 25542 27012 25594
rect 27064 25542 27076 25594
rect 27128 25542 27140 25594
rect 27192 25542 27204 25594
rect 27256 25542 30820 25594
rect 1104 25520 30820 25542
rect 12802 25440 12808 25492
rect 12860 25440 12866 25492
rect 12986 25440 12992 25492
rect 13044 25440 13050 25492
rect 13633 25483 13691 25489
rect 13633 25449 13645 25483
rect 13679 25480 13691 25483
rect 14366 25480 14372 25492
rect 13679 25452 14372 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 10597 25347 10655 25353
rect 10597 25313 10609 25347
rect 10643 25344 10655 25347
rect 10870 25344 10876 25356
rect 10643 25316 10876 25344
rect 10643 25313 10655 25316
rect 10597 25307 10655 25313
rect 10870 25304 10876 25316
rect 10928 25304 10934 25356
rect 13004 25353 13032 25440
rect 12989 25347 13047 25353
rect 12989 25313 13001 25347
rect 13035 25313 13047 25347
rect 12989 25307 13047 25313
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 8496 25248 9321 25276
rect 8496 25152 8524 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 12897 25279 12955 25285
rect 12897 25245 12909 25279
rect 12943 25276 12955 25279
rect 13648 25276 13676 25443
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 15289 25483 15347 25489
rect 15289 25449 15301 25483
rect 15335 25480 15347 25483
rect 15470 25480 15476 25492
rect 15335 25452 15476 25480
rect 15335 25449 15347 25452
rect 15289 25443 15347 25449
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 18506 25480 18512 25492
rect 17972 25452 18512 25480
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 17972 25344 18000 25452
rect 18506 25440 18512 25452
rect 18564 25440 18570 25492
rect 18049 25415 18107 25421
rect 18049 25381 18061 25415
rect 18095 25381 18107 25415
rect 18049 25375 18107 25381
rect 19245 25415 19303 25421
rect 19245 25381 19257 25415
rect 19291 25381 19303 25415
rect 19245 25375 19303 25381
rect 17819 25316 18000 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 12943 25248 13676 25276
rect 12943 25245 12955 25248
rect 12897 25239 12955 25245
rect 15194 25236 15200 25288
rect 15252 25276 15258 25288
rect 15473 25279 15531 25285
rect 15473 25276 15485 25279
rect 15252 25248 15485 25276
rect 15252 25236 15258 25248
rect 15473 25245 15485 25248
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 15562 25236 15568 25288
rect 15620 25236 15626 25288
rect 17681 25279 17739 25285
rect 17681 25245 17693 25279
rect 17727 25245 17739 25279
rect 17681 25239 17739 25245
rect 10873 25211 10931 25217
rect 10873 25177 10885 25211
rect 10919 25208 10931 25211
rect 10962 25208 10968 25220
rect 10919 25180 10968 25208
rect 10919 25177 10931 25180
rect 10873 25171 10931 25177
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 11882 25168 11888 25220
rect 11940 25168 11946 25220
rect 8478 25100 8484 25152
rect 8536 25100 8542 25152
rect 9398 25100 9404 25152
rect 9456 25100 9462 25152
rect 12342 25100 12348 25152
rect 12400 25100 12406 25152
rect 17696 25140 17724 25239
rect 18064 25208 18092 25375
rect 18785 25347 18843 25353
rect 18785 25313 18797 25347
rect 18831 25344 18843 25347
rect 19260 25344 19288 25375
rect 18831 25316 19288 25344
rect 18831 25313 18843 25316
rect 18785 25307 18843 25313
rect 20622 25236 20628 25288
rect 20680 25236 20686 25288
rect 20358 25211 20416 25217
rect 20358 25208 20370 25211
rect 18064 25180 20370 25208
rect 20358 25177 20370 25180
rect 20404 25177 20416 25211
rect 20358 25171 20416 25177
rect 17954 25140 17960 25152
rect 17696 25112 17960 25140
rect 17954 25100 17960 25112
rect 18012 25140 18018 25152
rect 18141 25143 18199 25149
rect 18141 25140 18153 25143
rect 18012 25112 18153 25140
rect 18012 25100 18018 25112
rect 18141 25109 18153 25112
rect 18187 25140 18199 25143
rect 18782 25140 18788 25152
rect 18187 25112 18788 25140
rect 18187 25109 18199 25112
rect 18141 25103 18199 25109
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 1104 25050 30820 25072
rect 1104 24998 5324 25050
rect 5376 24998 5388 25050
rect 5440 24998 5452 25050
rect 5504 24998 5516 25050
rect 5568 24998 5580 25050
rect 5632 24998 12752 25050
rect 12804 24998 12816 25050
rect 12868 24998 12880 25050
rect 12932 24998 12944 25050
rect 12996 24998 13008 25050
rect 13060 24998 20180 25050
rect 20232 24998 20244 25050
rect 20296 24998 20308 25050
rect 20360 24998 20372 25050
rect 20424 24998 20436 25050
rect 20488 24998 27608 25050
rect 27660 24998 27672 25050
rect 27724 24998 27736 25050
rect 27788 24998 27800 25050
rect 27852 24998 27864 25050
rect 27916 24998 30820 25050
rect 1104 24976 30820 24998
rect 10870 24936 10876 24948
rect 10336 24908 10876 24936
rect 9398 24828 9404 24880
rect 9456 24828 9462 24880
rect 8386 24800 8392 24812
rect 7774 24772 8392 24800
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 10336 24744 10364 24908
rect 10870 24896 10876 24908
rect 10928 24896 10934 24948
rect 10962 24896 10968 24948
rect 11020 24896 11026 24948
rect 11793 24939 11851 24945
rect 11793 24905 11805 24939
rect 11839 24936 11851 24939
rect 11882 24936 11888 24948
rect 11839 24908 11888 24936
rect 11839 24905 11851 24908
rect 11793 24899 11851 24905
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 16936 24871 16994 24877
rect 10796 24840 11008 24868
rect 10413 24803 10471 24809
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 6365 24735 6423 24741
rect 6365 24701 6377 24735
rect 6411 24732 6423 24735
rect 6411 24704 6500 24732
rect 6411 24701 6423 24704
rect 6365 24695 6423 24701
rect 6472 24608 6500 24704
rect 6638 24692 6644 24744
rect 6696 24692 6702 24744
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24732 8355 24735
rect 9306 24732 9312 24744
rect 8343 24704 9312 24732
rect 8343 24701 8355 24704
rect 8297 24695 8355 24701
rect 9306 24692 9312 24704
rect 9364 24692 9370 24744
rect 10042 24692 10048 24744
rect 10100 24692 10106 24744
rect 10318 24692 10324 24744
rect 10376 24692 10382 24744
rect 10428 24676 10456 24763
rect 10594 24760 10600 24812
rect 10652 24760 10658 24812
rect 10796 24809 10824 24840
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24769 10839 24803
rect 10980 24800 11008 24840
rect 16936 24837 16948 24871
rect 16982 24868 16994 24871
rect 17954 24868 17960 24880
rect 16982 24840 17960 24868
rect 16982 24837 16994 24840
rect 16936 24831 16994 24837
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 11054 24800 11060 24812
rect 10980 24772 11060 24800
rect 10781 24763 10839 24769
rect 10410 24624 10416 24676
rect 10468 24624 10474 24676
rect 6454 24556 6460 24608
rect 6512 24556 6518 24608
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 8113 24599 8171 24605
rect 8113 24596 8125 24599
rect 7984 24568 8125 24596
rect 7984 24556 7990 24568
rect 8113 24565 8125 24568
rect 8159 24565 8171 24599
rect 8113 24559 8171 24565
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 10704 24596 10732 24763
rect 11054 24760 11060 24772
rect 11112 24760 11118 24812
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24769 11943 24803
rect 11885 24763 11943 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12342 24800 12348 24812
rect 12299 24772 12348 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 11900 24732 11928 24763
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14214 24772 14749 24800
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 14829 24803 14887 24809
rect 14829 24769 14841 24803
rect 14875 24800 14887 24803
rect 15470 24800 15476 24812
rect 14875 24772 15476 24800
rect 14875 24769 14887 24772
rect 14829 24763 14887 24769
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24800 16727 24803
rect 16758 24800 16764 24812
rect 16715 24772 16764 24800
rect 16715 24769 16727 24772
rect 16669 24763 16727 24769
rect 16758 24760 16764 24772
rect 16816 24760 16822 24812
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 12805 24735 12863 24741
rect 11900 24704 12434 24732
rect 12406 24608 12434 24704
rect 12805 24701 12817 24735
rect 12851 24701 12863 24735
rect 12805 24695 12863 24701
rect 12069 24599 12127 24605
rect 12069 24596 12081 24599
rect 9732 24568 12081 24596
rect 9732 24556 9738 24568
rect 12069 24565 12081 24568
rect 12115 24565 12127 24599
rect 12406 24568 12440 24608
rect 12069 24559 12127 24565
rect 12434 24556 12440 24568
rect 12492 24556 12498 24608
rect 12820 24596 12848 24695
rect 13078 24692 13084 24744
rect 13136 24692 13142 24744
rect 18693 24735 18751 24741
rect 18693 24701 18705 24735
rect 18739 24701 18751 24735
rect 18693 24695 18751 24701
rect 14182 24624 14188 24676
rect 14240 24664 14246 24676
rect 14553 24667 14611 24673
rect 14553 24664 14565 24667
rect 14240 24636 14565 24664
rect 14240 24624 14246 24636
rect 14553 24633 14565 24636
rect 14599 24633 14611 24667
rect 14553 24627 14611 24633
rect 18049 24667 18107 24673
rect 18049 24633 18061 24667
rect 18095 24664 18107 24667
rect 18506 24664 18512 24676
rect 18095 24636 18512 24664
rect 18095 24633 18107 24636
rect 18049 24627 18107 24633
rect 18506 24624 18512 24636
rect 18564 24664 18570 24676
rect 18708 24664 18736 24695
rect 18564 24636 18736 24664
rect 18564 24624 18570 24636
rect 14366 24596 14372 24608
rect 12820 24568 14372 24596
rect 14366 24556 14372 24568
rect 14424 24556 14430 24608
rect 18138 24556 18144 24608
rect 18196 24556 18202 24608
rect 18874 24556 18880 24608
rect 18932 24556 18938 24608
rect 1104 24506 30820 24528
rect 1104 24454 4664 24506
rect 4716 24454 4728 24506
rect 4780 24454 4792 24506
rect 4844 24454 4856 24506
rect 4908 24454 4920 24506
rect 4972 24454 12092 24506
rect 12144 24454 12156 24506
rect 12208 24454 12220 24506
rect 12272 24454 12284 24506
rect 12336 24454 12348 24506
rect 12400 24454 19520 24506
rect 19572 24454 19584 24506
rect 19636 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 26948 24506
rect 27000 24454 27012 24506
rect 27064 24454 27076 24506
rect 27128 24454 27140 24506
rect 27192 24454 27204 24506
rect 27256 24454 30820 24506
rect 1104 24432 30820 24454
rect 6549 24395 6607 24401
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 6638 24392 6644 24404
rect 6595 24364 6644 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 6638 24352 6644 24364
rect 6696 24352 6702 24404
rect 8386 24352 8392 24404
rect 8444 24352 8450 24404
rect 9493 24395 9551 24401
rect 9493 24361 9505 24395
rect 9539 24392 9551 24395
rect 10042 24392 10048 24404
rect 9539 24364 10048 24392
rect 9539 24361 9551 24364
rect 9493 24355 9551 24361
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 18046 24392 18052 24404
rect 17083 24364 18052 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 8478 24284 8484 24336
rect 8536 24324 8542 24336
rect 12434 24324 12440 24336
rect 8536 24296 10548 24324
rect 8536 24284 8542 24296
rect 6454 24216 6460 24268
rect 6512 24256 6518 24268
rect 8294 24256 8300 24268
rect 6512 24228 8300 24256
rect 6512 24216 6518 24228
rect 8294 24216 8300 24228
rect 8352 24256 8358 24268
rect 10318 24256 10324 24268
rect 8352 24228 10324 24256
rect 8352 24216 8358 24228
rect 10318 24216 10324 24228
rect 10376 24256 10382 24268
rect 10413 24259 10471 24265
rect 10413 24256 10425 24259
rect 10376 24228 10425 24256
rect 10376 24216 10382 24228
rect 10413 24225 10425 24228
rect 10459 24225 10471 24259
rect 10520 24256 10548 24296
rect 12360 24296 12440 24324
rect 12360 24256 12388 24296
rect 12434 24284 12440 24296
rect 12492 24324 12498 24336
rect 16761 24327 16819 24333
rect 12492 24296 14688 24324
rect 12492 24284 12498 24296
rect 10520 24228 12480 24256
rect 10413 24219 10471 24225
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24188 6791 24191
rect 6779 24160 7052 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 4430 24080 4436 24132
rect 4488 24080 4494 24132
rect 5718 24080 5724 24132
rect 5776 24080 5782 24132
rect 6178 24080 6184 24132
rect 6236 24080 6242 24132
rect 6825 24123 6883 24129
rect 6825 24089 6837 24123
rect 6871 24089 6883 24123
rect 6825 24083 6883 24089
rect 6840 24052 6868 24083
rect 6914 24080 6920 24132
rect 6972 24080 6978 24132
rect 7024 24120 7052 24160
rect 7098 24148 7104 24200
rect 7156 24148 7162 24200
rect 7190 24148 7196 24200
rect 7248 24188 7254 24200
rect 7926 24188 7932 24200
rect 7248 24160 7932 24188
rect 7248 24148 7254 24160
rect 7926 24148 7932 24160
rect 7984 24188 7990 24200
rect 8113 24191 8171 24197
rect 8113 24188 8125 24191
rect 7984 24160 8125 24188
rect 7984 24148 7990 24160
rect 8113 24157 8125 24160
rect 8159 24157 8171 24191
rect 8481 24191 8539 24197
rect 8481 24188 8493 24191
rect 8113 24151 8171 24157
rect 8404 24160 8493 24188
rect 8404 24132 8432 24160
rect 8481 24157 8493 24160
rect 8527 24157 8539 24191
rect 8481 24151 8539 24157
rect 8941 24191 8999 24197
rect 8941 24157 8953 24191
rect 8987 24188 8999 24191
rect 8987 24160 9076 24188
rect 8987 24157 8999 24160
rect 8941 24151 8999 24157
rect 9048 24132 9076 24160
rect 9214 24148 9220 24200
rect 9272 24148 9278 24200
rect 12452 24197 12480 24228
rect 14366 24216 14372 24268
rect 14424 24256 14430 24268
rect 14553 24259 14611 24265
rect 14553 24256 14565 24259
rect 14424 24228 14565 24256
rect 14424 24216 14430 24228
rect 14553 24225 14565 24228
rect 14599 24225 14611 24259
rect 14660 24256 14688 24296
rect 16761 24293 16773 24327
rect 16807 24324 16819 24327
rect 17052 24324 17080 24355
rect 18046 24352 18052 24364
rect 18104 24352 18110 24404
rect 18506 24352 18512 24404
rect 18564 24352 18570 24404
rect 18969 24395 19027 24401
rect 18969 24361 18981 24395
rect 19015 24392 19027 24395
rect 19058 24392 19064 24404
rect 19015 24364 19064 24392
rect 19015 24361 19027 24364
rect 18969 24355 19027 24361
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 16807 24296 17080 24324
rect 16807 24293 16819 24296
rect 16761 24287 16819 24293
rect 15470 24256 15476 24268
rect 14660 24228 15476 24256
rect 14553 24219 14611 24225
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16390 24216 16396 24268
rect 16448 24216 16454 24268
rect 18524 24265 18552 24352
rect 18782 24284 18788 24336
rect 18840 24284 18846 24336
rect 18509 24259 18567 24265
rect 18509 24225 18521 24259
rect 18555 24225 18567 24259
rect 18509 24219 18567 24225
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24188 13415 24191
rect 14182 24188 14188 24200
rect 13403 24160 14188 24188
rect 13403 24157 13415 24160
rect 13357 24151 13415 24157
rect 7024 24092 8156 24120
rect 8128 24064 8156 24092
rect 8386 24080 8392 24132
rect 8444 24080 8450 24132
rect 9030 24080 9036 24132
rect 9088 24080 9094 24132
rect 9122 24080 9128 24132
rect 9180 24080 9186 24132
rect 7561 24055 7619 24061
rect 7561 24052 7573 24055
rect 6840 24024 7573 24052
rect 7561 24021 7573 24024
rect 7607 24021 7619 24055
rect 7561 24015 7619 24021
rect 8110 24012 8116 24064
rect 8168 24052 8174 24064
rect 9324 24052 9352 24151
rect 14182 24148 14188 24160
rect 14240 24148 14246 24200
rect 14274 24148 14280 24200
rect 14332 24148 14338 24200
rect 16758 24148 16764 24200
rect 16816 24188 16822 24200
rect 18417 24191 18475 24197
rect 18417 24188 18429 24191
rect 16816 24160 18429 24188
rect 16816 24148 16822 24160
rect 18417 24157 18429 24160
rect 18463 24188 18475 24191
rect 19242 24188 19248 24200
rect 18463 24160 19248 24188
rect 18463 24157 18475 24160
rect 18417 24151 18475 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 10686 24080 10692 24132
rect 10744 24080 10750 24132
rect 12345 24123 12403 24129
rect 12345 24120 12357 24123
rect 11914 24092 12357 24120
rect 12345 24089 12357 24092
rect 12391 24089 12403 24123
rect 12345 24083 12403 24089
rect 14829 24123 14887 24129
rect 14829 24089 14841 24123
rect 14875 24089 14887 24123
rect 14829 24083 14887 24089
rect 11054 24052 11060 24064
rect 8168 24024 11060 24052
rect 8168 24012 8174 24024
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11974 24012 11980 24064
rect 12032 24052 12038 24064
rect 12161 24055 12219 24061
rect 12161 24052 12173 24055
rect 12032 24024 12173 24052
rect 12032 24012 12038 24024
rect 12161 24021 12173 24024
rect 12207 24021 12219 24055
rect 12161 24015 12219 24021
rect 13078 24012 13084 24064
rect 13136 24052 13142 24064
rect 13449 24055 13507 24061
rect 13449 24052 13461 24055
rect 13136 24024 13461 24052
rect 13136 24012 13142 24024
rect 13449 24021 13461 24024
rect 13495 24021 13507 24055
rect 13449 24015 13507 24021
rect 14461 24055 14519 24061
rect 14461 24021 14473 24055
rect 14507 24052 14519 24055
rect 14844 24052 14872 24083
rect 15562 24080 15568 24132
rect 15620 24080 15626 24132
rect 18138 24080 18144 24132
rect 18196 24129 18202 24132
rect 18196 24120 18208 24129
rect 18196 24092 18241 24120
rect 18196 24083 18208 24092
rect 18196 24080 18202 24083
rect 14507 24024 14872 24052
rect 14507 24021 14519 24024
rect 14461 24015 14519 24021
rect 16298 24012 16304 24064
rect 16356 24012 16362 24064
rect 16850 24012 16856 24064
rect 16908 24012 16914 24064
rect 1104 23962 30820 23984
rect 1104 23910 5324 23962
rect 5376 23910 5388 23962
rect 5440 23910 5452 23962
rect 5504 23910 5516 23962
rect 5568 23910 5580 23962
rect 5632 23910 12752 23962
rect 12804 23910 12816 23962
rect 12868 23910 12880 23962
rect 12932 23910 12944 23962
rect 12996 23910 13008 23962
rect 13060 23910 20180 23962
rect 20232 23910 20244 23962
rect 20296 23910 20308 23962
rect 20360 23910 20372 23962
rect 20424 23910 20436 23962
rect 20488 23910 27608 23962
rect 27660 23910 27672 23962
rect 27724 23910 27736 23962
rect 27788 23910 27800 23962
rect 27852 23910 27864 23962
rect 27916 23910 30820 23962
rect 1104 23888 30820 23910
rect 5718 23808 5724 23860
rect 5776 23848 5782 23860
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 5776 23820 5825 23848
rect 5776 23808 5782 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 6178 23808 6184 23860
rect 6236 23848 6242 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 6236 23820 6377 23848
rect 6236 23808 6242 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 7837 23851 7895 23857
rect 7837 23848 7849 23851
rect 6365 23811 6423 23817
rect 6748 23820 7849 23848
rect 6748 23789 6776 23820
rect 7837 23817 7849 23820
rect 7883 23817 7895 23851
rect 10505 23851 10563 23857
rect 7837 23811 7895 23817
rect 7944 23820 9076 23848
rect 6733 23783 6791 23789
rect 6733 23749 6745 23783
rect 6779 23749 6791 23783
rect 7098 23780 7104 23792
rect 6733 23743 6791 23749
rect 6840 23752 7104 23780
rect 5905 23715 5963 23721
rect 5905 23681 5917 23715
rect 5951 23681 5963 23715
rect 5905 23675 5963 23681
rect 5920 23644 5948 23675
rect 6546 23672 6552 23724
rect 6604 23672 6610 23724
rect 6641 23715 6699 23721
rect 6641 23681 6653 23715
rect 6687 23712 6699 23715
rect 6840 23712 6868 23752
rect 7098 23740 7104 23752
rect 7156 23780 7162 23792
rect 7944 23780 7972 23820
rect 8386 23780 8392 23792
rect 7156 23752 7972 23780
rect 8036 23752 8392 23780
rect 7156 23740 7162 23752
rect 6687 23684 6868 23712
rect 6917 23715 6975 23721
rect 6687 23681 6699 23684
rect 6641 23675 6699 23681
rect 6917 23681 6929 23715
rect 6963 23712 6975 23715
rect 7006 23712 7012 23724
rect 6963 23684 7012 23712
rect 6963 23681 6975 23684
rect 6917 23675 6975 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 8036 23644 8064 23752
rect 8386 23740 8392 23752
rect 8444 23740 8450 23792
rect 9048 23724 9076 23820
rect 10505 23817 10517 23851
rect 10551 23848 10563 23851
rect 10686 23848 10692 23860
rect 10551 23820 10692 23848
rect 10551 23817 10563 23820
rect 10505 23811 10563 23817
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 14182 23848 14188 23860
rect 13556 23820 14188 23848
rect 10137 23783 10195 23789
rect 10137 23749 10149 23783
rect 10183 23780 10195 23783
rect 10778 23780 10784 23792
rect 10183 23752 10784 23780
rect 10183 23749 10195 23752
rect 10137 23743 10195 23749
rect 10778 23740 10784 23752
rect 10836 23740 10842 23792
rect 13556 23724 13584 23820
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14274 23808 14280 23860
rect 14332 23848 14338 23860
rect 14553 23851 14611 23857
rect 14553 23848 14565 23851
rect 14332 23820 14565 23848
rect 14332 23808 14338 23820
rect 14553 23817 14565 23820
rect 14599 23817 14611 23851
rect 14553 23811 14611 23817
rect 15562 23808 15568 23860
rect 15620 23808 15626 23860
rect 16850 23808 16856 23860
rect 16908 23808 16914 23860
rect 18874 23808 18880 23860
rect 18932 23808 18938 23860
rect 14200 23780 14228 23808
rect 16298 23780 16304 23792
rect 14200 23752 14694 23780
rect 8110 23672 8116 23724
rect 8168 23672 8174 23724
rect 8205 23715 8263 23721
rect 8205 23681 8217 23715
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 5920 23616 8064 23644
rect 8220 23576 8248 23675
rect 9030 23672 9036 23724
rect 9088 23712 9094 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9088 23684 9965 23712
rect 9088 23672 9094 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23681 10287 23715
rect 10229 23675 10287 23681
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23712 10379 23715
rect 11054 23712 11060 23724
rect 10367 23684 11060 23712
rect 10367 23681 10379 23684
rect 10321 23675 10379 23681
rect 7852 23548 8248 23576
rect 9968 23576 9996 23675
rect 10244 23644 10272 23675
rect 11054 23672 11060 23684
rect 11112 23672 11118 23724
rect 13538 23672 13544 23724
rect 13596 23672 13602 23724
rect 13630 23672 13636 23724
rect 13688 23712 13694 23724
rect 13725 23715 13783 23721
rect 13725 23712 13737 23715
rect 13688 23684 13737 23712
rect 13688 23672 13694 23684
rect 13725 23681 13737 23684
rect 13771 23712 13783 23715
rect 14550 23712 14556 23724
rect 13771 23684 14556 23712
rect 13771 23681 13783 23684
rect 13725 23675 13783 23681
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 14666 23721 14694 23752
rect 14844 23752 16304 23780
rect 14645 23715 14703 23721
rect 14645 23681 14657 23715
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 14734 23672 14740 23724
rect 14792 23712 14798 23724
rect 14844 23721 14872 23752
rect 16298 23740 16304 23752
rect 16356 23740 16362 23792
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 14792 23684 14841 23712
rect 14792 23672 14798 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 15470 23672 15476 23724
rect 15528 23712 15534 23724
rect 15933 23715 15991 23721
rect 15528 23684 15884 23712
rect 15528 23672 15534 23684
rect 10502 23644 10508 23656
rect 10244 23616 10508 23644
rect 10502 23604 10508 23616
rect 10560 23604 10566 23656
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 13740 23616 14105 23644
rect 10410 23576 10416 23588
rect 9968 23548 10416 23576
rect 7852 23520 7880 23548
rect 10410 23536 10416 23548
rect 10468 23576 10474 23588
rect 11146 23576 11152 23588
rect 10468 23548 11152 23576
rect 10468 23536 10474 23548
rect 11146 23536 11152 23548
rect 11204 23536 11210 23588
rect 13740 23520 13768 23616
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 15856 23644 15884 23684
rect 15933 23681 15945 23715
rect 15979 23712 15991 23715
rect 16868 23712 16896 23808
rect 18592 23783 18650 23789
rect 18592 23749 18604 23783
rect 18638 23780 18650 23783
rect 18892 23780 18920 23808
rect 18638 23752 18920 23780
rect 18638 23749 18650 23752
rect 18592 23743 18650 23749
rect 25406 23740 25412 23792
rect 25464 23740 25470 23792
rect 15979 23684 16896 23712
rect 15979 23681 15991 23684
rect 15933 23675 15991 23681
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23712 23535 23715
rect 23523 23684 24440 23712
rect 23523 23681 23535 23684
rect 23477 23675 23535 23681
rect 16022 23644 16028 23656
rect 14424 23616 15792 23644
rect 15856 23616 16028 23644
rect 14424 23604 14430 23616
rect 15764 23585 15792 23616
rect 16022 23604 16028 23616
rect 16080 23604 16086 23656
rect 18325 23647 18383 23653
rect 18325 23613 18337 23647
rect 18371 23613 18383 23647
rect 18325 23607 18383 23613
rect 14461 23579 14519 23585
rect 14461 23545 14473 23579
rect 14507 23576 14519 23579
rect 15749 23579 15807 23585
rect 14507 23548 14780 23576
rect 14507 23545 14519 23548
rect 14461 23539 14519 23545
rect 7834 23468 7840 23520
rect 7892 23468 7898 23520
rect 8202 23468 8208 23520
rect 8260 23468 8266 23520
rect 13541 23511 13599 23517
rect 13541 23477 13553 23511
rect 13587 23508 13599 23511
rect 13722 23508 13728 23520
rect 13587 23480 13728 23508
rect 13587 23477 13599 23480
rect 13541 23471 13599 23477
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 14752 23517 14780 23548
rect 15749 23545 15761 23579
rect 15795 23545 15807 23579
rect 15749 23539 15807 23545
rect 14737 23511 14795 23517
rect 14737 23477 14749 23511
rect 14783 23508 14795 23511
rect 14826 23508 14832 23520
rect 14783 23480 14832 23508
rect 14783 23477 14795 23480
rect 14737 23471 14795 23477
rect 14826 23468 14832 23480
rect 14884 23468 14890 23520
rect 18340 23508 18368 23607
rect 24412 23588 24440 23684
rect 24486 23604 24492 23656
rect 24544 23604 24550 23656
rect 24765 23647 24823 23653
rect 24765 23613 24777 23647
rect 24811 23644 24823 23647
rect 24854 23644 24860 23656
rect 24811 23616 24860 23644
rect 24811 23613 24823 23616
rect 24765 23607 24823 23613
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 24394 23536 24400 23588
rect 24452 23536 24458 23588
rect 19242 23508 19248 23520
rect 18340 23480 19248 23508
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 19705 23511 19763 23517
rect 19705 23508 19717 23511
rect 19484 23480 19717 23508
rect 19484 23468 19490 23480
rect 19705 23477 19717 23480
rect 19751 23477 19763 23511
rect 19705 23471 19763 23477
rect 20530 23468 20536 23520
rect 20588 23508 20594 23520
rect 20625 23511 20683 23517
rect 20625 23508 20637 23511
rect 20588 23480 20637 23508
rect 20588 23468 20594 23480
rect 20625 23477 20637 23480
rect 20671 23477 20683 23511
rect 20625 23471 20683 23477
rect 23474 23468 23480 23520
rect 23532 23508 23538 23520
rect 23569 23511 23627 23517
rect 23569 23508 23581 23511
rect 23532 23480 23581 23508
rect 23532 23468 23538 23480
rect 23569 23477 23581 23480
rect 23615 23477 23627 23511
rect 23569 23471 23627 23477
rect 26237 23511 26295 23517
rect 26237 23477 26249 23511
rect 26283 23508 26295 23511
rect 27430 23508 27436 23520
rect 26283 23480 27436 23508
rect 26283 23477 26295 23480
rect 26237 23471 26295 23477
rect 27430 23468 27436 23480
rect 27488 23468 27494 23520
rect 1104 23418 30820 23440
rect 1104 23366 4664 23418
rect 4716 23366 4728 23418
rect 4780 23366 4792 23418
rect 4844 23366 4856 23418
rect 4908 23366 4920 23418
rect 4972 23366 12092 23418
rect 12144 23366 12156 23418
rect 12208 23366 12220 23418
rect 12272 23366 12284 23418
rect 12336 23366 12348 23418
rect 12400 23366 19520 23418
rect 19572 23366 19584 23418
rect 19636 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 26948 23418
rect 27000 23366 27012 23418
rect 27064 23366 27076 23418
rect 27128 23366 27140 23418
rect 27192 23366 27204 23418
rect 27256 23366 30820 23418
rect 1104 23344 30820 23366
rect 6365 23307 6423 23313
rect 6365 23273 6377 23307
rect 6411 23304 6423 23307
rect 6546 23304 6552 23316
rect 6411 23276 6552 23304
rect 6411 23273 6423 23276
rect 6365 23267 6423 23273
rect 6546 23264 6552 23276
rect 6604 23264 6610 23316
rect 9309 23307 9367 23313
rect 6656 23276 7328 23304
rect 6656 23180 6684 23276
rect 6748 23208 7236 23236
rect 6638 23128 6644 23180
rect 6696 23128 6702 23180
rect 6748 23177 6776 23208
rect 6733 23171 6791 23177
rect 6733 23137 6745 23171
rect 6779 23137 6791 23171
rect 7098 23168 7104 23180
rect 6733 23131 6791 23137
rect 6840 23140 7104 23168
rect 6840 23109 6868 23140
rect 7098 23128 7104 23140
rect 7156 23128 7162 23180
rect 6549 23103 6607 23109
rect 6549 23069 6561 23103
rect 6595 23069 6607 23103
rect 6549 23063 6607 23069
rect 6825 23103 6883 23109
rect 6825 23069 6837 23103
rect 6871 23069 6883 23103
rect 6825 23063 6883 23069
rect 7009 23103 7067 23109
rect 7009 23069 7021 23103
rect 7055 23069 7067 23103
rect 7009 23063 7067 23069
rect 6564 22976 6592 23063
rect 7024 22976 7052 23063
rect 7101 23035 7159 23041
rect 7101 23001 7113 23035
rect 7147 23032 7159 23035
rect 7208 23032 7236 23208
rect 7300 23168 7328 23276
rect 7760 23276 8340 23304
rect 7760 23245 7788 23276
rect 7745 23239 7803 23245
rect 7745 23205 7757 23239
rect 7791 23205 7803 23239
rect 7745 23199 7803 23205
rect 7834 23196 7840 23248
rect 7892 23196 7898 23248
rect 8018 23196 8024 23248
rect 8076 23236 8082 23248
rect 8205 23239 8263 23245
rect 8205 23236 8217 23239
rect 8076 23208 8217 23236
rect 8076 23196 8082 23208
rect 8205 23205 8217 23208
rect 8251 23205 8263 23239
rect 8205 23199 8263 23205
rect 8312 23168 8340 23276
rect 9309 23273 9321 23307
rect 9355 23304 9367 23307
rect 9582 23304 9588 23316
rect 9355 23276 9588 23304
rect 9355 23273 9367 23276
rect 9309 23267 9367 23273
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 11054 23264 11060 23316
rect 11112 23304 11118 23316
rect 12069 23307 12127 23313
rect 12069 23304 12081 23307
rect 11112 23276 12081 23304
rect 11112 23264 11118 23276
rect 12069 23273 12081 23276
rect 12115 23273 12127 23307
rect 12069 23267 12127 23273
rect 12250 23264 12256 23316
rect 12308 23264 12314 23316
rect 13173 23307 13231 23313
rect 13173 23273 13185 23307
rect 13219 23304 13231 23307
rect 13538 23304 13544 23316
rect 13219 23276 13544 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 13538 23264 13544 23276
rect 13596 23264 13602 23316
rect 24854 23264 24860 23316
rect 24912 23304 24918 23316
rect 24949 23307 25007 23313
rect 24949 23304 24961 23307
rect 24912 23276 24961 23304
rect 24912 23264 24918 23276
rect 24949 23273 24961 23276
rect 24995 23273 25007 23307
rect 24949 23267 25007 23273
rect 25406 23264 25412 23316
rect 25464 23264 25470 23316
rect 27430 23264 27436 23316
rect 27488 23304 27494 23316
rect 27709 23307 27767 23313
rect 27709 23304 27721 23307
rect 27488 23276 27721 23304
rect 27488 23264 27494 23276
rect 27709 23273 27721 23276
rect 27755 23273 27767 23307
rect 27709 23267 27767 23273
rect 11146 23196 11152 23248
rect 11204 23236 11210 23248
rect 12268 23236 12296 23264
rect 11204 23208 12296 23236
rect 12989 23239 13047 23245
rect 11204 23196 11210 23208
rect 12989 23205 13001 23239
rect 13035 23236 13047 23239
rect 13262 23236 13268 23248
rect 13035 23208 13268 23236
rect 13035 23205 13047 23208
rect 12989 23199 13047 23205
rect 12434 23177 12440 23180
rect 7300 23140 7880 23168
rect 7650 23060 7656 23112
rect 7708 23060 7714 23112
rect 7852 23032 7880 23140
rect 8220 23140 8340 23168
rect 12391 23171 12440 23177
rect 8220 23112 8248 23140
rect 12391 23137 12403 23171
rect 12437 23137 12440 23171
rect 12391 23131 12440 23137
rect 12434 23128 12440 23131
rect 12492 23168 12498 23180
rect 13004 23168 13032 23199
rect 13262 23196 13268 23208
rect 13320 23196 13326 23248
rect 13630 23196 13636 23248
rect 13688 23196 13694 23248
rect 12492 23140 13032 23168
rect 13541 23171 13599 23177
rect 12492 23128 12498 23140
rect 13541 23137 13553 23171
rect 13587 23168 13599 23171
rect 13648 23168 13676 23196
rect 13587 23140 13676 23168
rect 13587 23137 13599 23140
rect 13541 23131 13599 23137
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19978 23168 19984 23180
rect 19392 23140 19984 23168
rect 19392 23128 19398 23140
rect 19978 23128 19984 23140
rect 20036 23168 20042 23180
rect 20349 23171 20407 23177
rect 20349 23168 20361 23171
rect 20036 23140 20361 23168
rect 20036 23128 20042 23140
rect 20349 23137 20361 23140
rect 20395 23168 20407 23171
rect 20622 23168 20628 23180
rect 20395 23140 20628 23168
rect 20395 23137 20407 23140
rect 20349 23131 20407 23137
rect 20622 23128 20628 23140
rect 20680 23168 20686 23180
rect 22465 23171 22523 23177
rect 22465 23168 22477 23171
rect 20680 23140 22477 23168
rect 20680 23128 20686 23140
rect 22465 23137 22477 23140
rect 22511 23168 22523 23171
rect 23934 23168 23940 23180
rect 22511 23140 23940 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 23934 23128 23940 23140
rect 23992 23168 23998 23180
rect 24486 23168 24492 23180
rect 23992 23140 24492 23168
rect 23992 23128 23998 23140
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 7926 23060 7932 23112
rect 7984 23109 7990 23112
rect 7984 23103 7999 23109
rect 7987 23069 7999 23103
rect 7984 23063 7999 23069
rect 7984 23060 7990 23063
rect 8202 23060 8208 23112
rect 8260 23060 8266 23112
rect 9214 23060 9220 23112
rect 9272 23060 9278 23112
rect 11974 23060 11980 23112
rect 12032 23060 12038 23112
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23069 12311 23103
rect 12253 23063 12311 23069
rect 15105 23103 15163 23109
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15654 23100 15660 23112
rect 15151 23072 15660 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 8573 23035 8631 23041
rect 8573 23032 8585 23035
rect 7147 23004 7788 23032
rect 7852 23004 8585 23032
rect 7147 23001 7159 23004
rect 7101 22995 7159 23001
rect 7760 22976 7788 23004
rect 8573 23001 8585 23004
rect 8619 23032 8631 23035
rect 9232 23032 9260 23060
rect 9493 23035 9551 23041
rect 9493 23032 9505 23035
rect 8619 23004 9168 23032
rect 9232 23004 9505 23032
rect 8619 23001 8631 23004
rect 8573 22995 8631 23001
rect 6546 22924 6552 22976
rect 6604 22924 6610 22976
rect 7006 22924 7012 22976
rect 7064 22924 7070 22976
rect 7466 22924 7472 22976
rect 7524 22924 7530 22976
rect 7742 22924 7748 22976
rect 7800 22924 7806 22976
rect 7834 22924 7840 22976
rect 7892 22964 7898 22976
rect 8113 22967 8171 22973
rect 8113 22964 8125 22967
rect 7892 22936 8125 22964
rect 7892 22924 7898 22936
rect 8113 22933 8125 22936
rect 8159 22964 8171 22967
rect 8478 22964 8484 22976
rect 8159 22936 8484 22964
rect 8159 22933 8171 22936
rect 8113 22927 8171 22933
rect 8478 22924 8484 22936
rect 8536 22924 8542 22976
rect 9140 22973 9168 23004
rect 9493 23001 9505 23004
rect 9539 23001 9551 23035
rect 9493 22995 9551 23001
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 12268 23032 12296 23063
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 22373 23103 22431 23109
rect 22373 23069 22385 23103
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 11940 23004 12296 23032
rect 15764 23032 15792 23063
rect 16022 23032 16028 23044
rect 15764 23004 16028 23032
rect 11940 22992 11946 23004
rect 16022 22992 16028 23004
rect 16080 22992 16086 23044
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 20625 23035 20683 23041
rect 20625 23032 20637 23035
rect 20588 23004 20637 23032
rect 20588 22992 20594 23004
rect 20625 23001 20637 23004
rect 20671 23001 20683 23035
rect 22281 23035 22339 23041
rect 22281 23032 22293 23035
rect 21850 23004 22293 23032
rect 20625 22995 20683 23001
rect 22281 23001 22293 23004
rect 22327 23001 22339 23035
rect 22281 22995 22339 23001
rect 9306 22973 9312 22976
rect 9125 22967 9183 22973
rect 9125 22933 9137 22967
rect 9171 22933 9183 22967
rect 9125 22927 9183 22933
rect 9293 22967 9312 22973
rect 9293 22933 9305 22967
rect 9293 22927 9312 22933
rect 9306 22924 9312 22927
rect 9364 22924 9370 22976
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 11606 22964 11612 22976
rect 10560 22936 11612 22964
rect 10560 22924 10566 22936
rect 11606 22924 11612 22936
rect 11664 22964 11670 22976
rect 11793 22967 11851 22973
rect 11793 22964 11805 22967
rect 11664 22936 11805 22964
rect 11664 22924 11670 22936
rect 11793 22933 11805 22936
rect 11839 22933 11851 22967
rect 11793 22927 11851 22933
rect 12250 22924 12256 22976
rect 12308 22964 12314 22976
rect 12713 22967 12771 22973
rect 12713 22964 12725 22967
rect 12308 22936 12725 22964
rect 12308 22924 12314 22936
rect 12713 22933 12725 22936
rect 12759 22933 12771 22967
rect 12713 22927 12771 22933
rect 13170 22924 13176 22976
rect 13228 22924 13234 22976
rect 14918 22924 14924 22976
rect 14976 22924 14982 22976
rect 15657 22967 15715 22973
rect 15657 22933 15669 22967
rect 15703 22964 15715 22967
rect 15746 22964 15752 22976
rect 15703 22936 15752 22964
rect 15703 22933 15715 22936
rect 15657 22927 15715 22933
rect 15746 22924 15752 22936
rect 15804 22924 15810 22976
rect 21910 22924 21916 22976
rect 21968 22964 21974 22976
rect 22097 22967 22155 22973
rect 22097 22964 22109 22967
rect 21968 22936 22109 22964
rect 21968 22924 21974 22936
rect 22097 22933 22109 22936
rect 22143 22933 22155 22967
rect 22388 22964 22416 23063
rect 25130 23060 25136 23112
rect 25188 23060 25194 23112
rect 25317 23103 25375 23109
rect 25317 23100 25329 23103
rect 25240 23072 25329 23100
rect 25240 23044 25268 23072
rect 25317 23069 25329 23072
rect 25363 23069 25375 23103
rect 25317 23063 25375 23069
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 27982 23100 27988 23112
rect 27663 23072 27988 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 22738 22992 22744 23044
rect 22796 22992 22802 23044
rect 23474 22992 23480 23044
rect 23532 22992 23538 23044
rect 24394 23032 24400 23044
rect 24044 23004 24400 23032
rect 24044 22964 24072 23004
rect 24394 22992 24400 23004
rect 24452 23032 24458 23044
rect 25222 23032 25228 23044
rect 24452 23004 25228 23032
rect 24452 22992 24458 23004
rect 25222 22992 25228 23004
rect 25280 22992 25286 23044
rect 22388 22936 24072 22964
rect 22097 22927 22155 22933
rect 24210 22924 24216 22976
rect 24268 22924 24274 22976
rect 28077 22967 28135 22973
rect 28077 22933 28089 22967
rect 28123 22964 28135 22967
rect 28902 22964 28908 22976
rect 28123 22936 28908 22964
rect 28123 22933 28135 22936
rect 28077 22927 28135 22933
rect 28902 22924 28908 22936
rect 28960 22924 28966 22976
rect 1104 22874 30820 22896
rect 1104 22822 5324 22874
rect 5376 22822 5388 22874
rect 5440 22822 5452 22874
rect 5504 22822 5516 22874
rect 5568 22822 5580 22874
rect 5632 22822 12752 22874
rect 12804 22822 12816 22874
rect 12868 22822 12880 22874
rect 12932 22822 12944 22874
rect 12996 22822 13008 22874
rect 13060 22822 20180 22874
rect 20232 22822 20244 22874
rect 20296 22822 20308 22874
rect 20360 22822 20372 22874
rect 20424 22822 20436 22874
rect 20488 22822 27608 22874
rect 27660 22822 27672 22874
rect 27724 22822 27736 22874
rect 27788 22822 27800 22874
rect 27852 22822 27864 22874
rect 27916 22822 30820 22874
rect 1104 22800 30820 22822
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 6365 22763 6423 22769
rect 4488 22732 5488 22760
rect 4488 22720 4494 22732
rect 5166 22692 5172 22704
rect 4080 22664 5172 22692
rect 4080 22633 4108 22664
rect 5166 22652 5172 22664
rect 5224 22652 5230 22704
rect 5460 22633 5488 22732
rect 6365 22729 6377 22763
rect 6411 22729 6423 22763
rect 6365 22723 6423 22729
rect 6086 22692 6092 22704
rect 5552 22664 6092 22692
rect 4065 22627 4123 22633
rect 4065 22593 4077 22627
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 5445 22627 5503 22633
rect 5031 22596 5396 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 4154 22516 4160 22568
rect 4212 22516 4218 22568
rect 4709 22559 4767 22565
rect 4709 22525 4721 22559
rect 4755 22556 4767 22559
rect 5261 22559 5319 22565
rect 5261 22556 5273 22559
rect 4755 22528 5273 22556
rect 4755 22525 4767 22528
rect 4709 22519 4767 22525
rect 5261 22525 5273 22528
rect 5307 22525 5319 22559
rect 5368 22556 5396 22596
rect 5445 22593 5457 22627
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 5552 22556 5580 22664
rect 6086 22652 6092 22664
rect 6144 22652 6150 22704
rect 6181 22695 6239 22701
rect 6181 22661 6193 22695
rect 6227 22692 6239 22695
rect 6380 22692 6408 22723
rect 6638 22720 6644 22772
rect 6696 22720 6702 22772
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7101 22763 7159 22769
rect 7101 22760 7113 22763
rect 6972 22732 7113 22760
rect 6972 22720 6978 22732
rect 7101 22729 7113 22732
rect 7147 22729 7159 22763
rect 7101 22723 7159 22729
rect 7650 22720 7656 22772
rect 7708 22760 7714 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 7708 22732 7757 22760
rect 7708 22720 7714 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 9033 22763 9091 22769
rect 7745 22723 7803 22729
rect 8036 22732 8984 22760
rect 8036 22692 8064 22732
rect 8956 22692 8984 22732
rect 9033 22729 9045 22763
rect 9079 22760 9091 22763
rect 9122 22760 9128 22772
rect 9079 22732 9128 22760
rect 9079 22729 9091 22732
rect 9033 22723 9091 22729
rect 9122 22720 9128 22732
rect 9180 22720 9186 22772
rect 10502 22720 10508 22772
rect 10560 22720 10566 22772
rect 10689 22763 10747 22769
rect 10689 22729 10701 22763
rect 10735 22729 10747 22763
rect 10689 22723 10747 22729
rect 9585 22695 9643 22701
rect 9585 22692 9597 22695
rect 6227 22664 6408 22692
rect 6656 22664 7328 22692
rect 6227 22661 6239 22664
rect 6181 22655 6239 22661
rect 5902 22584 5908 22636
rect 5960 22584 5966 22636
rect 5997 22627 6055 22633
rect 5997 22593 6009 22627
rect 6043 22593 6055 22627
rect 6656 22624 6684 22664
rect 5997 22587 6055 22593
rect 6104 22596 6684 22624
rect 6733 22627 6791 22633
rect 5368 22528 5580 22556
rect 5629 22559 5687 22565
rect 5261 22519 5319 22525
rect 5629 22525 5641 22559
rect 5675 22556 5687 22559
rect 6012 22556 6040 22587
rect 5675 22528 6040 22556
rect 5675 22525 5687 22528
rect 5629 22519 5687 22525
rect 5644 22488 5672 22519
rect 5092 22460 5672 22488
rect 5092 22432 5120 22460
rect 4801 22423 4859 22429
rect 4801 22389 4813 22423
rect 4847 22420 4859 22423
rect 4982 22420 4988 22432
rect 4847 22392 4988 22420
rect 4847 22389 4859 22392
rect 4801 22383 4859 22389
rect 4982 22380 4988 22392
rect 5040 22380 5046 22432
rect 5074 22380 5080 22432
rect 5132 22380 5138 22432
rect 5169 22423 5227 22429
rect 5169 22389 5181 22423
rect 5215 22420 5227 22423
rect 6104 22420 6132 22596
rect 6733 22593 6745 22627
rect 6779 22624 6791 22627
rect 6914 22624 6920 22636
rect 6779 22596 6920 22624
rect 6779 22593 6791 22596
rect 6733 22587 6791 22593
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22624 7067 22627
rect 7190 22624 7196 22636
rect 7055 22596 7196 22624
rect 7055 22593 7067 22596
rect 7009 22587 7067 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7300 22633 7328 22664
rect 7576 22664 8064 22692
rect 8588 22664 8892 22692
rect 8956 22664 9597 22692
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 6546 22565 6552 22568
rect 6524 22559 6552 22565
rect 6524 22525 6536 22559
rect 6604 22556 6610 22568
rect 7576 22556 7604 22664
rect 8588 22636 8616 22664
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 6604 22528 7604 22556
rect 6524 22519 6552 22525
rect 6546 22516 6552 22519
rect 6604 22516 6610 22528
rect 6181 22491 6239 22497
rect 6181 22457 6193 22491
rect 6227 22488 6239 22491
rect 7668 22488 7696 22587
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7800 22596 7941 22624
rect 7800 22584 7806 22596
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 7929 22587 7987 22593
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 8478 22584 8484 22636
rect 8536 22584 8542 22636
rect 8570 22584 8576 22636
rect 8628 22584 8634 22636
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 8754 22584 8760 22636
rect 8812 22584 8818 22636
rect 8864 22633 8892 22664
rect 9585 22661 9597 22664
rect 9631 22692 9643 22695
rect 10704 22692 10732 22723
rect 10778 22720 10784 22772
rect 10836 22720 10842 22772
rect 11974 22720 11980 22772
rect 12032 22720 12038 22772
rect 12250 22720 12256 22772
rect 12308 22760 12314 22772
rect 12529 22763 12587 22769
rect 12529 22760 12541 22763
rect 12308 22732 12541 22760
rect 12308 22720 12314 22732
rect 12529 22729 12541 22732
rect 12575 22729 12587 22763
rect 14918 22760 14924 22772
rect 12529 22723 12587 22729
rect 14752 22732 14924 22760
rect 9631 22664 10359 22692
rect 10704 22664 11284 22692
rect 9631 22661 9643 22664
rect 9585 22655 9643 22661
rect 8854 22627 8912 22633
rect 8854 22593 8866 22627
rect 8900 22624 8912 22627
rect 9674 22624 9680 22636
rect 8900 22596 9680 22624
rect 8900 22593 8912 22596
rect 8854 22587 8912 22593
rect 9674 22584 9680 22596
rect 9732 22584 9738 22636
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 9815 22596 9904 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 8018 22516 8024 22568
rect 8076 22556 8082 22568
rect 8205 22559 8263 22565
rect 8205 22556 8217 22559
rect 8076 22528 8217 22556
rect 8076 22516 8082 22528
rect 8205 22525 8217 22528
rect 8251 22556 8263 22559
rect 8251 22528 9736 22556
rect 8251 22525 8263 22528
rect 8205 22519 8263 22525
rect 6227 22460 7696 22488
rect 8113 22491 8171 22497
rect 6227 22457 6239 22460
rect 6181 22451 6239 22457
rect 8113 22457 8125 22491
rect 8159 22488 8171 22491
rect 9708 22488 9736 22528
rect 9876 22500 9904 22596
rect 9950 22584 9956 22636
rect 10008 22584 10014 22636
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22624 10103 22627
rect 10331 22624 10359 22664
rect 10965 22627 11023 22633
rect 10965 22624 10977 22627
rect 10091 22596 10272 22624
rect 10331 22596 10977 22624
rect 10091 22593 10103 22596
rect 10045 22587 10103 22593
rect 9968 22556 9996 22584
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 9968 22528 10149 22556
rect 10137 22525 10149 22528
rect 10183 22525 10195 22559
rect 10244 22556 10272 22596
rect 10965 22593 10977 22596
rect 11011 22593 11023 22627
rect 10965 22587 11023 22593
rect 11054 22584 11060 22636
rect 11112 22584 11118 22636
rect 11256 22633 11284 22664
rect 11422 22652 11428 22704
rect 11480 22692 11486 22704
rect 11992 22692 12020 22720
rect 11480 22664 11928 22692
rect 11992 22664 12296 22692
rect 11480 22652 11486 22664
rect 11241 22627 11299 22633
rect 11241 22593 11253 22627
rect 11287 22593 11299 22627
rect 11241 22587 11299 22593
rect 11333 22627 11391 22633
rect 11333 22593 11345 22627
rect 11379 22624 11391 22627
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 11379 22596 11529 22624
rect 11379 22593 11391 22596
rect 11333 22587 11391 22593
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11517 22587 11575 22593
rect 11698 22584 11704 22636
rect 11756 22584 11762 22636
rect 11790 22584 11796 22636
rect 11848 22584 11854 22636
rect 11900 22633 11928 22664
rect 11885 22627 11943 22633
rect 11885 22593 11897 22627
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 11974 22584 11980 22636
rect 12032 22633 12038 22636
rect 12268 22633 12296 22664
rect 12342 22652 12348 22704
rect 12400 22652 12406 22704
rect 14752 22701 14780 22732
rect 14918 22720 14924 22732
rect 14976 22720 14982 22772
rect 17862 22720 17868 22772
rect 17920 22760 17926 22772
rect 20717 22763 20775 22769
rect 17920 22732 20668 22760
rect 17920 22720 17926 22732
rect 14737 22695 14795 22701
rect 12452 22664 12664 22692
rect 12452 22633 12480 22664
rect 12032 22627 12061 22633
rect 12049 22593 12061 22627
rect 12032 22587 12061 22593
rect 12253 22627 12311 22633
rect 12253 22593 12265 22627
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 12430 22627 12488 22633
rect 12430 22593 12442 22627
rect 12476 22593 12488 22627
rect 12430 22587 12488 22593
rect 12032 22584 12038 22587
rect 12161 22559 12219 22565
rect 10244 22528 10548 22556
rect 10137 22519 10195 22525
rect 9858 22488 9864 22500
rect 8159 22460 8294 22488
rect 9708 22460 9864 22488
rect 8159 22457 8171 22460
rect 8113 22451 8171 22457
rect 5215 22392 6132 22420
rect 5215 22389 5227 22392
rect 5169 22383 5227 22389
rect 7466 22380 7472 22432
rect 7524 22380 7530 22432
rect 8266 22420 8294 22460
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 10520 22429 10548 22528
rect 12161 22525 12173 22559
rect 12207 22556 12219 22559
rect 12636 22556 12664 22664
rect 14737 22661 14749 22695
rect 14783 22661 14795 22695
rect 14737 22655 14795 22661
rect 15746 22652 15752 22704
rect 15804 22652 15810 22704
rect 20640 22692 20668 22732
rect 20717 22729 20729 22763
rect 20763 22760 20775 22763
rect 20806 22760 20812 22772
rect 20763 22732 20812 22760
rect 20763 22729 20775 22732
rect 20717 22723 20775 22729
rect 20806 22720 20812 22732
rect 20864 22720 20870 22772
rect 21085 22763 21143 22769
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 21910 22760 21916 22772
rect 21131 22732 21916 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 23017 22763 23075 22769
rect 23017 22760 23029 22763
rect 22796 22732 23029 22760
rect 22796 22720 22802 22732
rect 23017 22729 23029 22732
rect 23063 22729 23075 22763
rect 23017 22723 23075 22729
rect 23569 22763 23627 22769
rect 23569 22729 23581 22763
rect 23615 22729 23627 22763
rect 23569 22723 23627 22729
rect 20640 22664 21312 22692
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22593 12771 22627
rect 12713 22587 12771 22593
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 13262 22624 13268 22636
rect 13035 22596 13268 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 12207 22528 12388 22556
rect 12207 22525 12219 22528
rect 12161 22519 12219 22525
rect 11790 22448 11796 22500
rect 11848 22488 11854 22500
rect 12250 22488 12256 22500
rect 11848 22460 12256 22488
rect 11848 22448 11854 22460
rect 12250 22448 12256 22460
rect 12308 22448 12314 22500
rect 12360 22488 12388 22528
rect 12544 22528 12664 22556
rect 12728 22556 12756 22587
rect 13262 22584 13268 22596
rect 13320 22584 13326 22636
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 14366 22584 14372 22636
rect 14424 22624 14430 22636
rect 14461 22627 14519 22633
rect 14461 22624 14473 22627
rect 14424 22596 14473 22624
rect 14424 22584 14430 22596
rect 14461 22593 14473 22596
rect 14507 22593 14519 22627
rect 14461 22587 14519 22593
rect 18046 22584 18052 22636
rect 18104 22584 18110 22636
rect 19521 22627 19579 22633
rect 19521 22624 19533 22627
rect 19352 22596 19533 22624
rect 13556 22556 13584 22584
rect 12728 22528 13584 22556
rect 12544 22500 12572 22528
rect 15194 22516 15200 22568
rect 15252 22556 15258 22568
rect 16485 22559 16543 22565
rect 16485 22556 16497 22559
rect 15252 22528 16497 22556
rect 15252 22516 15258 22528
rect 16485 22525 16497 22528
rect 16531 22525 16543 22559
rect 16485 22519 16543 22525
rect 16669 22559 16727 22565
rect 16669 22525 16681 22559
rect 16715 22556 16727 22559
rect 16715 22528 16804 22556
rect 16715 22525 16727 22528
rect 16669 22519 16727 22525
rect 12526 22488 12532 22500
rect 12360 22460 12532 22488
rect 12526 22448 12532 22460
rect 12584 22448 12590 22500
rect 16776 22432 16804 22528
rect 16942 22516 16948 22568
rect 17000 22516 17006 22568
rect 19061 22491 19119 22497
rect 19061 22488 19073 22491
rect 18432 22460 19073 22488
rect 10505 22423 10563 22429
rect 10505 22420 10517 22423
rect 8266 22392 10517 22420
rect 10505 22389 10517 22392
rect 10551 22420 10563 22423
rect 10686 22420 10692 22432
rect 10551 22392 10692 22420
rect 10551 22389 10563 22392
rect 10505 22383 10563 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 10962 22380 10968 22432
rect 11020 22420 11026 22432
rect 12897 22423 12955 22429
rect 12897 22420 12909 22423
rect 11020 22392 12909 22420
rect 11020 22380 11026 22392
rect 12897 22389 12909 22392
rect 12943 22420 12955 22423
rect 13262 22420 13268 22432
rect 12943 22392 13268 22420
rect 12943 22389 12955 22392
rect 12897 22383 12955 22389
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 16758 22380 16764 22432
rect 16816 22380 16822 22432
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18432 22429 18460 22460
rect 19061 22457 19073 22460
rect 19107 22457 19119 22491
rect 19061 22451 19119 22457
rect 18417 22423 18475 22429
rect 18417 22420 18429 22423
rect 18012 22392 18429 22420
rect 18012 22380 18018 22392
rect 18417 22389 18429 22392
rect 18463 22389 18475 22423
rect 18417 22383 18475 22389
rect 18966 22380 18972 22432
rect 19024 22380 19030 22432
rect 19076 22420 19104 22451
rect 19352 22420 19380 22596
rect 19521 22593 19533 22596
rect 19567 22593 19579 22627
rect 19521 22587 19579 22593
rect 19429 22559 19487 22565
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 19475 22528 19840 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 19812 22497 19840 22528
rect 21174 22516 21180 22568
rect 21232 22516 21238 22568
rect 21284 22565 21312 22664
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22624 23259 22627
rect 23584 22624 23612 22723
rect 25130 22720 25136 22772
rect 25188 22720 25194 22772
rect 25593 22763 25651 22769
rect 25593 22729 25605 22763
rect 25639 22760 25651 22763
rect 27522 22760 27528 22772
rect 25639 22732 27528 22760
rect 25639 22729 25651 22732
rect 25593 22723 25651 22729
rect 27522 22720 27528 22732
rect 27580 22720 27586 22772
rect 28902 22720 28908 22772
rect 28960 22720 28966 22772
rect 23937 22695 23995 22701
rect 23937 22661 23949 22695
rect 23983 22692 23995 22695
rect 24210 22692 24216 22704
rect 23983 22664 24216 22692
rect 23983 22661 23995 22664
rect 23937 22655 23995 22661
rect 24210 22652 24216 22664
rect 24268 22692 24274 22704
rect 24762 22692 24768 22704
rect 24268 22664 24768 22692
rect 24268 22652 24274 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 28721 22695 28779 22701
rect 28721 22692 28733 22695
rect 28000 22664 28733 22692
rect 23247 22596 23612 22624
rect 24029 22627 24087 22633
rect 23247 22593 23259 22596
rect 23201 22587 23259 22593
rect 24029 22593 24041 22627
rect 24075 22624 24087 22627
rect 25038 22624 25044 22636
rect 24075 22596 25044 22624
rect 24075 22593 24087 22596
rect 24029 22587 24087 22593
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 25498 22584 25504 22636
rect 25556 22584 25562 22636
rect 28000 22633 28028 22664
rect 28721 22661 28733 22664
rect 28767 22661 28779 22695
rect 28920 22692 28948 22720
rect 28920 22664 29408 22692
rect 28721 22655 28779 22661
rect 27985 22627 28043 22633
rect 27985 22624 27997 22627
rect 26804 22596 27997 22624
rect 21269 22559 21327 22565
rect 21269 22525 21281 22559
rect 21315 22556 21327 22559
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 21315 22528 24133 22556
rect 21315 22525 21327 22528
rect 21269 22519 21327 22525
rect 24121 22525 24133 22528
rect 24167 22556 24179 22559
rect 25406 22556 25412 22568
rect 24167 22528 25412 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 25406 22516 25412 22528
rect 25464 22556 25470 22568
rect 26804 22565 26832 22596
rect 27985 22593 27997 22596
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 28166 22584 28172 22636
rect 28224 22584 28230 22636
rect 29380 22633 29408 22664
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22622 28503 22627
rect 28905 22627 28963 22633
rect 28491 22594 28580 22622
rect 28491 22593 28503 22594
rect 28445 22587 28503 22593
rect 25685 22559 25743 22565
rect 25685 22556 25697 22559
rect 25464 22528 25697 22556
rect 25464 22516 25470 22528
rect 25685 22525 25697 22528
rect 25731 22525 25743 22559
rect 25685 22519 25743 22525
rect 26329 22559 26387 22565
rect 26329 22525 26341 22559
rect 26375 22525 26387 22559
rect 26329 22519 26387 22525
rect 26789 22559 26847 22565
rect 26789 22525 26801 22559
rect 26835 22525 26847 22559
rect 26789 22519 26847 22525
rect 26973 22559 27031 22565
rect 26973 22525 26985 22559
rect 27019 22556 27031 22559
rect 28552 22556 28580 22594
rect 28905 22593 28917 22627
rect 28951 22593 28963 22627
rect 28905 22587 28963 22593
rect 29181 22627 29239 22633
rect 29181 22593 29193 22627
rect 29227 22593 29239 22627
rect 29181 22587 29239 22593
rect 29365 22627 29423 22633
rect 29365 22593 29377 22627
rect 29411 22593 29423 22627
rect 29365 22587 29423 22593
rect 28920 22556 28948 22587
rect 27019 22528 27384 22556
rect 27019 22525 27031 22528
rect 26973 22519 27031 22525
rect 19797 22491 19855 22497
rect 19797 22457 19809 22491
rect 19843 22488 19855 22491
rect 20162 22488 20168 22500
rect 19843 22460 20168 22488
rect 19843 22457 19855 22460
rect 19797 22451 19855 22457
rect 20162 22448 20168 22460
rect 20220 22448 20226 22500
rect 24762 22448 24768 22500
rect 24820 22488 24826 22500
rect 26344 22488 26372 22519
rect 24820 22460 26372 22488
rect 24820 22448 24826 22460
rect 19426 22420 19432 22432
rect 19076 22392 19432 22420
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 19886 22380 19892 22432
rect 19944 22420 19950 22432
rect 19981 22423 20039 22429
rect 19981 22420 19993 22423
rect 19944 22392 19993 22420
rect 19944 22380 19950 22392
rect 19981 22389 19993 22392
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 26050 22420 26056 22432
rect 22152 22392 26056 22420
rect 22152 22380 22158 22392
rect 26050 22380 26056 22392
rect 26108 22380 26114 22432
rect 26344 22420 26372 22460
rect 26697 22491 26755 22497
rect 26697 22457 26709 22491
rect 26743 22488 26755 22491
rect 26988 22488 27016 22519
rect 26743 22460 27016 22488
rect 27249 22491 27307 22497
rect 26743 22457 26755 22460
rect 26697 22451 26755 22457
rect 27249 22457 27261 22491
rect 27295 22457 27307 22491
rect 27249 22451 27307 22457
rect 27264 22420 27292 22451
rect 27356 22432 27384 22528
rect 28552 22528 28948 22556
rect 26344 22392 27292 22420
rect 27338 22380 27344 22432
rect 27396 22380 27402 22432
rect 27433 22423 27491 22429
rect 27433 22389 27445 22423
rect 27479 22420 27491 22423
rect 28552 22420 28580 22528
rect 28810 22448 28816 22500
rect 28868 22488 28874 22500
rect 29196 22488 29224 22587
rect 28868 22460 29224 22488
rect 28868 22448 28874 22460
rect 27479 22392 28580 22420
rect 27479 22389 27491 22392
rect 27433 22383 27491 22389
rect 28626 22380 28632 22432
rect 28684 22380 28690 22432
rect 29086 22380 29092 22432
rect 29144 22380 29150 22432
rect 29270 22380 29276 22432
rect 29328 22380 29334 22432
rect 1104 22330 30820 22352
rect 1104 22278 4664 22330
rect 4716 22278 4728 22330
rect 4780 22278 4792 22330
rect 4844 22278 4856 22330
rect 4908 22278 4920 22330
rect 4972 22278 12092 22330
rect 12144 22278 12156 22330
rect 12208 22278 12220 22330
rect 12272 22278 12284 22330
rect 12336 22278 12348 22330
rect 12400 22278 19520 22330
rect 19572 22278 19584 22330
rect 19636 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 26948 22330
rect 27000 22278 27012 22330
rect 27064 22278 27076 22330
rect 27128 22278 27140 22330
rect 27192 22278 27204 22330
rect 27256 22278 30820 22330
rect 1104 22256 30820 22278
rect 4154 22176 4160 22228
rect 4212 22176 4218 22228
rect 4893 22219 4951 22225
rect 4893 22185 4905 22219
rect 4939 22216 4951 22219
rect 4982 22216 4988 22228
rect 4939 22188 4988 22216
rect 4939 22185 4951 22188
rect 4893 22179 4951 22185
rect 4982 22176 4988 22188
rect 5040 22176 5046 22228
rect 5902 22176 5908 22228
rect 5960 22216 5966 22228
rect 6730 22216 6736 22228
rect 5960 22188 6736 22216
rect 5960 22176 5966 22188
rect 6730 22176 6736 22188
rect 6788 22216 6794 22228
rect 8570 22216 8576 22228
rect 6788 22188 8576 22216
rect 6788 22176 6794 22188
rect 8570 22176 8576 22188
rect 8628 22176 8634 22228
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 8941 22219 8999 22225
rect 8941 22216 8953 22219
rect 8720 22188 8953 22216
rect 8720 22176 8726 22188
rect 8941 22185 8953 22188
rect 8987 22185 8999 22219
rect 8941 22179 8999 22185
rect 11609 22219 11667 22225
rect 11609 22185 11621 22219
rect 11655 22216 11667 22219
rect 11698 22216 11704 22228
rect 11655 22188 11704 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 11698 22176 11704 22188
rect 11756 22176 11762 22228
rect 13630 22216 13636 22228
rect 13464 22188 13636 22216
rect 9232 22120 9720 22148
rect 4430 22040 4436 22092
rect 4488 22080 4494 22092
rect 4488 22052 4936 22080
rect 4488 22040 4494 22052
rect 4338 21972 4344 22024
rect 4396 21972 4402 22024
rect 4908 22021 4936 22052
rect 5166 22040 5172 22092
rect 5224 22080 5230 22092
rect 7190 22080 7196 22092
rect 5224 22052 7196 22080
rect 5224 22040 5230 22052
rect 7190 22040 7196 22052
rect 7248 22040 7254 22092
rect 9232 22024 9260 22120
rect 9306 22040 9312 22092
rect 9364 22040 9370 22092
rect 4617 22015 4675 22021
rect 4617 22012 4629 22015
rect 4448 21984 4629 22012
rect 4448 21888 4476 21984
rect 4617 21981 4629 21984
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4709 22015 4767 22021
rect 4709 21981 4721 22015
rect 4755 21981 4767 22015
rect 4709 21975 4767 21981
rect 4893 22015 4951 22021
rect 4893 21981 4905 22015
rect 4939 21981 4951 22015
rect 4893 21975 4951 21981
rect 4724 21944 4752 21975
rect 4982 21972 4988 22024
rect 5040 21972 5046 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9214 22012 9220 22024
rect 9171 21984 9220 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9214 21972 9220 21984
rect 9272 21972 9278 22024
rect 9324 22012 9352 22040
rect 9692 22021 9720 22120
rect 9858 22108 9864 22160
rect 9916 22148 9922 22160
rect 10962 22148 10968 22160
rect 9916 22120 10968 22148
rect 9916 22108 9922 22120
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 10505 22083 10563 22089
rect 9784 22052 10088 22080
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 9324 21984 9413 22012
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9677 22015 9735 22021
rect 9677 21981 9689 22015
rect 9723 21981 9735 22015
rect 9677 21975 9735 21981
rect 5000 21944 5028 21972
rect 4724 21916 5028 21944
rect 9416 21944 9444 21975
rect 9784 21944 9812 22052
rect 10060 22024 10088 22052
rect 10505 22049 10517 22083
rect 10551 22080 10563 22083
rect 11054 22080 11060 22092
rect 10551 22052 11060 22080
rect 10551 22049 10563 22052
rect 10505 22043 10563 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 13464 22089 13492 22188
rect 13630 22176 13636 22188
rect 13688 22176 13694 22228
rect 15654 22176 15660 22228
rect 15712 22176 15718 22228
rect 16942 22176 16948 22228
rect 17000 22176 17006 22228
rect 18046 22176 18052 22228
rect 18104 22216 18110 22228
rect 18141 22219 18199 22225
rect 18141 22216 18153 22219
rect 18104 22188 18153 22216
rect 18104 22176 18110 22188
rect 18141 22185 18153 22188
rect 18187 22185 18199 22219
rect 18141 22179 18199 22185
rect 18969 22219 19027 22225
rect 18969 22185 18981 22219
rect 19015 22216 19027 22219
rect 19245 22219 19303 22225
rect 19245 22216 19257 22219
rect 19015 22188 19257 22216
rect 19015 22185 19027 22188
rect 18969 22179 19027 22185
rect 19245 22185 19257 22188
rect 19291 22185 19303 22219
rect 19245 22179 19303 22185
rect 19536 22188 20024 22216
rect 17221 22151 17279 22157
rect 17221 22117 17233 22151
rect 17267 22117 17279 22151
rect 17221 22111 17279 22117
rect 13449 22083 13507 22089
rect 13449 22080 13461 22083
rect 13004 22052 13461 22080
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 9416 21916 9812 21944
rect 4430 21836 4436 21888
rect 4488 21836 4494 21888
rect 4522 21836 4528 21888
rect 4580 21836 4586 21888
rect 4614 21836 4620 21888
rect 4672 21876 4678 21888
rect 4724 21876 4752 21916
rect 9876 21888 9904 21975
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10413 22015 10471 22021
rect 10413 22012 10425 22015
rect 10100 21984 10425 22012
rect 10100 21972 10106 21984
rect 10413 21981 10425 21984
rect 10459 22012 10471 22015
rect 10459 21984 11744 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 11716 21956 11744 21984
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 13004 22021 13032 22052
rect 13449 22049 13461 22052
rect 13495 22049 13507 22083
rect 13658 22083 13716 22089
rect 13658 22080 13670 22083
rect 13449 22043 13507 22049
rect 13648 22049 13670 22080
rect 13704 22049 13716 22083
rect 13648 22043 13716 22049
rect 14476 22052 15516 22080
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 21981 12863 22015
rect 12805 21975 12863 21981
rect 12989 22015 13047 22021
rect 12989 21981 13001 22015
rect 13035 21981 13047 22015
rect 12989 21975 13047 21981
rect 11422 21904 11428 21956
rect 11480 21904 11486 21956
rect 11698 21904 11704 21956
rect 11756 21944 11762 21956
rect 11793 21947 11851 21953
rect 11793 21944 11805 21947
rect 11756 21916 11805 21944
rect 11756 21904 11762 21916
rect 11793 21913 11805 21916
rect 11839 21913 11851 21947
rect 11793 21907 11851 21913
rect 11977 21947 12035 21953
rect 11977 21913 11989 21947
rect 12023 21944 12035 21947
rect 12544 21944 12572 21972
rect 12023 21916 12572 21944
rect 12023 21913 12035 21916
rect 11977 21907 12035 21913
rect 4672 21848 4752 21876
rect 4672 21836 4678 21848
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9490 21836 9496 21888
rect 9548 21836 9554 21888
rect 9858 21836 9864 21888
rect 9916 21836 9922 21888
rect 11440 21876 11468 21904
rect 11992 21876 12020 21907
rect 11440 21848 12020 21876
rect 12526 21836 12532 21888
rect 12584 21836 12590 21888
rect 12636 21876 12664 21975
rect 12820 21944 12848 21975
rect 13170 21972 13176 22024
rect 13228 21972 13234 22024
rect 13078 21944 13084 21956
rect 12820 21916 13084 21944
rect 13078 21904 13084 21916
rect 13136 21944 13142 21956
rect 13648 21944 13676 22043
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 14476 22021 14504 22052
rect 14461 22015 14519 22021
rect 14461 22012 14473 22015
rect 14056 21984 14473 22012
rect 14056 21972 14062 21984
rect 14461 21981 14473 21984
rect 14507 21981 14519 22015
rect 14461 21975 14519 21981
rect 14737 22015 14795 22021
rect 14737 21981 14749 22015
rect 14783 22012 14795 22015
rect 14826 22012 14832 22024
rect 14783 21984 14832 22012
rect 14783 21981 14795 21984
rect 14737 21975 14795 21981
rect 14826 21972 14832 21984
rect 14884 21972 14890 22024
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 15488 22021 15516 22052
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 21981 15531 22015
rect 15473 21975 15531 21981
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 17236 22012 17264 22111
rect 17862 22108 17868 22160
rect 17920 22108 17926 22160
rect 17770 22080 17776 22092
rect 17731 22052 17776 22080
rect 17770 22040 17776 22052
rect 17828 22080 17834 22092
rect 17880 22080 17908 22108
rect 17828 22052 17908 22080
rect 17828 22040 17834 22052
rect 18690 22040 18696 22092
rect 18748 22080 18754 22092
rect 19536 22080 19564 22188
rect 18748 22052 19564 22080
rect 19705 22083 19763 22089
rect 18748 22040 18754 22052
rect 19705 22049 19717 22083
rect 19751 22080 19763 22083
rect 19996 22080 20024 22188
rect 21174 22176 21180 22228
rect 21232 22216 21238 22228
rect 21453 22219 21511 22225
rect 21453 22216 21465 22219
rect 21232 22188 21465 22216
rect 21232 22176 21238 22188
rect 21453 22185 21465 22188
rect 21499 22185 21511 22219
rect 21453 22179 21511 22185
rect 25038 22176 25044 22228
rect 25096 22216 25102 22228
rect 25961 22219 26019 22225
rect 25961 22216 25973 22219
rect 25096 22188 25973 22216
rect 25096 22176 25102 22188
rect 25961 22185 25973 22188
rect 26007 22185 26019 22219
rect 27430 22216 27436 22228
rect 25961 22179 26019 22185
rect 26068 22188 27436 22216
rect 20530 22108 20536 22160
rect 20588 22108 20594 22160
rect 21910 22108 21916 22160
rect 21968 22148 21974 22160
rect 22281 22151 22339 22157
rect 22281 22148 22293 22151
rect 21968 22120 22293 22148
rect 21968 22108 21974 22120
rect 22281 22117 22293 22120
rect 22327 22117 22339 22151
rect 22281 22111 22339 22117
rect 25409 22151 25467 22157
rect 25409 22117 25421 22151
rect 25455 22117 25467 22151
rect 25409 22111 25467 22117
rect 20548 22080 20576 22108
rect 22833 22083 22891 22089
rect 22833 22080 22845 22083
rect 19751 22052 20576 22080
rect 21652 22052 22845 22080
rect 19751 22049 19763 22052
rect 19705 22043 19763 22049
rect 17175 21984 17264 22012
rect 17589 22015 17647 22021
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 17954 22012 17960 22024
rect 17635 21984 17960 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 21981 18107 22015
rect 18049 21975 18107 21981
rect 13136 21916 13676 21944
rect 13740 21916 14596 21944
rect 13136 21904 13142 21916
rect 13170 21876 13176 21888
rect 12636 21848 13176 21876
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 13740 21876 13768 21916
rect 14568 21888 14596 21916
rect 15286 21904 15292 21956
rect 15344 21904 15350 21956
rect 16758 21904 16764 21956
rect 16816 21944 16822 21956
rect 18064 21944 18092 21975
rect 19058 21972 19064 22024
rect 19116 21972 19122 22024
rect 19242 21972 19248 22024
rect 19300 22012 19306 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19300 21984 19441 22012
rect 19300 21972 19306 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19521 22015 19579 22021
rect 19521 21981 19533 22015
rect 19567 22012 19579 22015
rect 19610 22012 19616 22024
rect 19567 21984 19616 22012
rect 19567 21981 19579 21984
rect 19521 21975 19579 21981
rect 19610 21972 19616 21984
rect 19668 21972 19674 22024
rect 19794 21972 19800 22024
rect 19852 21972 19858 22024
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 21652 22021 21680 22052
rect 22833 22049 22845 22052
rect 22879 22049 22891 22083
rect 25424 22080 25452 22111
rect 25498 22108 25504 22160
rect 25556 22148 25562 22160
rect 26068 22148 26096 22188
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 27890 22176 27896 22228
rect 27948 22176 27954 22228
rect 28000 22188 29592 22216
rect 27448 22148 27476 22176
rect 25556 22120 26096 22148
rect 26160 22120 27292 22148
rect 27448 22120 27660 22148
rect 25556 22108 25562 22120
rect 26160 22080 26188 22120
rect 25424 22052 26188 22080
rect 22833 22043 22891 22049
rect 26234 22040 26240 22092
rect 26292 22080 26298 22092
rect 26292 22052 26464 22080
rect 26292 22040 26298 22052
rect 20533 22015 20591 22021
rect 20533 22012 20545 22015
rect 20220 21984 20545 22012
rect 20220 21972 20226 21984
rect 20533 21981 20545 21984
rect 20579 21981 20591 22015
rect 20533 21975 20591 21981
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 21637 22015 21695 22021
rect 20763 21984 21036 22012
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 16816 21916 18092 21944
rect 16816 21904 16822 21916
rect 18506 21904 18512 21956
rect 18564 21944 18570 21956
rect 20625 21947 20683 21953
rect 20625 21944 20637 21947
rect 18564 21916 20637 21944
rect 18564 21904 18570 21916
rect 20625 21913 20637 21916
rect 20671 21913 20683 21947
rect 20625 21907 20683 21913
rect 13596 21848 13768 21876
rect 13596 21836 13602 21848
rect 13814 21836 13820 21888
rect 13872 21836 13878 21888
rect 14550 21836 14556 21888
rect 14608 21836 14614 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 18598 21836 18604 21888
rect 18656 21836 18662 21888
rect 19794 21836 19800 21888
rect 19852 21876 19858 21888
rect 20806 21876 20812 21888
rect 19852 21848 20812 21876
rect 19852 21836 19858 21848
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 21008 21885 21036 21984
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 22094 21972 22100 22024
rect 22152 21972 22158 22024
rect 22741 22015 22799 22021
rect 22741 21981 22753 22015
rect 22787 21981 22799 22015
rect 22741 21975 22799 21981
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 21174 21904 21180 21956
rect 21232 21904 21238 21956
rect 21361 21947 21419 21953
rect 21361 21913 21373 21947
rect 21407 21944 21419 21947
rect 21542 21944 21548 21956
rect 21407 21916 21548 21944
rect 21407 21913 21419 21916
rect 21361 21907 21419 21913
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 21729 21947 21787 21953
rect 21729 21913 21741 21947
rect 21775 21913 21787 21947
rect 21729 21907 21787 21913
rect 20993 21879 21051 21885
rect 20993 21845 21005 21879
rect 21039 21876 21051 21879
rect 21744 21876 21772 21907
rect 21818 21904 21824 21956
rect 21876 21904 21882 21956
rect 21959 21947 22017 21953
rect 21959 21913 21971 21947
rect 22005 21944 22017 21947
rect 22554 21944 22560 21956
rect 22005 21916 22560 21944
rect 22005 21913 22017 21916
rect 21959 21907 22017 21913
rect 22554 21904 22560 21916
rect 22612 21904 22618 21956
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 22756 21944 22784 21975
rect 22695 21916 22784 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 21039 21848 21772 21876
rect 21039 21845 21051 21848
rect 20993 21839 21051 21845
rect 22186 21836 22192 21888
rect 22244 21836 22250 21888
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 22664 21876 22692 21907
rect 22830 21904 22836 21956
rect 22888 21944 22894 21956
rect 22940 21944 22968 21975
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 24084 21984 24409 22012
rect 24084 21972 24090 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 22012 24731 22015
rect 26145 22015 26203 22021
rect 24719 21984 25360 22012
rect 24719 21981 24731 21984
rect 24673 21975 24731 21981
rect 25332 21956 25360 21984
rect 26145 21981 26157 22015
rect 26191 21981 26203 22015
rect 26145 21975 26203 21981
rect 22888 21916 24440 21944
rect 22888 21904 22894 21916
rect 24412 21888 24440 21916
rect 25314 21904 25320 21956
rect 25372 21904 25378 21956
rect 22336 21848 22692 21876
rect 22336 21836 22342 21848
rect 24394 21836 24400 21888
rect 24452 21836 24458 21888
rect 26160 21876 26188 21975
rect 26326 21972 26332 22024
rect 26384 22021 26390 22024
rect 26384 22015 26400 22021
rect 26388 21981 26400 22015
rect 26436 22012 26464 22052
rect 26712 22021 26740 22120
rect 27264 22024 27292 22120
rect 26559 22015 26617 22021
rect 26559 22012 26571 22015
rect 26436 21984 26571 22012
rect 26384 21975 26400 21981
rect 26559 21981 26571 21984
rect 26605 21981 26617 22015
rect 26559 21975 26617 21981
rect 26697 22015 26755 22021
rect 26697 21981 26709 22015
rect 26743 21981 26755 22015
rect 26697 21975 26755 21981
rect 26384 21972 26390 21975
rect 26878 21972 26884 22024
rect 26936 21972 26942 22024
rect 27246 21972 27252 22024
rect 27304 21972 27310 22024
rect 27632 22021 27660 22120
rect 27617 22015 27675 22021
rect 27617 21981 27629 22015
rect 27663 21981 27675 22015
rect 27617 21975 27675 21981
rect 26234 21904 26240 21956
rect 26292 21904 26298 21956
rect 26467 21947 26525 21953
rect 26467 21913 26479 21947
rect 26513 21944 26525 21947
rect 28000 21944 28028 22188
rect 28077 22151 28135 22157
rect 28077 22117 28089 22151
rect 28123 22148 28135 22151
rect 28166 22148 28172 22160
rect 28123 22120 28172 22148
rect 28123 22117 28135 22120
rect 28077 22111 28135 22117
rect 28166 22108 28172 22120
rect 28224 22148 28230 22160
rect 28810 22148 28816 22160
rect 28224 22120 28816 22148
rect 28224 22108 28230 22120
rect 28810 22108 28816 22120
rect 28868 22108 28874 22160
rect 29564 22157 29592 22188
rect 29549 22151 29607 22157
rect 29549 22117 29561 22151
rect 29595 22117 29607 22151
rect 29549 22111 29607 22117
rect 28721 22083 28779 22089
rect 28721 22049 28733 22083
rect 28767 22080 28779 22083
rect 29825 22083 29883 22089
rect 29825 22080 29837 22083
rect 28767 22052 29837 22080
rect 28767 22049 28779 22052
rect 28721 22043 28779 22049
rect 29825 22049 29837 22052
rect 29871 22049 29883 22083
rect 29825 22043 29883 22049
rect 28626 21972 28632 22024
rect 28684 21972 28690 22024
rect 28810 21972 28816 22024
rect 28868 21972 28874 22024
rect 29086 21972 29092 22024
rect 29144 22012 29150 22024
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29144 21984 29929 22012
rect 29144 21972 29150 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 29917 21975 29975 21981
rect 26513 21916 28028 21944
rect 26513 21913 26525 21916
rect 26467 21907 26525 21913
rect 29270 21904 29276 21956
rect 29328 21904 29334 21956
rect 26697 21879 26755 21885
rect 26697 21876 26709 21879
rect 26160 21848 26709 21876
rect 26697 21845 26709 21848
rect 26743 21845 26755 21879
rect 26697 21839 26755 21845
rect 26878 21836 26884 21888
rect 26936 21876 26942 21888
rect 28074 21876 28080 21888
rect 26936 21848 28080 21876
rect 26936 21836 26942 21848
rect 28074 21836 28080 21848
rect 28132 21836 28138 21888
rect 28905 21879 28963 21885
rect 28905 21845 28917 21879
rect 28951 21876 28963 21879
rect 29362 21876 29368 21888
rect 28951 21848 29368 21876
rect 28951 21845 28963 21848
rect 28905 21839 28963 21845
rect 29362 21836 29368 21848
rect 29420 21836 29426 21888
rect 1104 21786 30820 21808
rect 1104 21734 5324 21786
rect 5376 21734 5388 21786
rect 5440 21734 5452 21786
rect 5504 21734 5516 21786
rect 5568 21734 5580 21786
rect 5632 21734 12752 21786
rect 12804 21734 12816 21786
rect 12868 21734 12880 21786
rect 12932 21734 12944 21786
rect 12996 21734 13008 21786
rect 13060 21734 20180 21786
rect 20232 21734 20244 21786
rect 20296 21734 20308 21786
rect 20360 21734 20372 21786
rect 20424 21734 20436 21786
rect 20488 21734 27608 21786
rect 27660 21734 27672 21786
rect 27724 21734 27736 21786
rect 27788 21734 27800 21786
rect 27852 21734 27864 21786
rect 27916 21734 30820 21786
rect 1104 21712 30820 21734
rect 4338 21632 4344 21684
rect 4396 21672 4402 21684
rect 5261 21675 5319 21681
rect 5261 21672 5273 21675
rect 4396 21644 5273 21672
rect 4396 21632 4402 21644
rect 5261 21641 5273 21644
rect 5307 21641 5319 21675
rect 5261 21635 5319 21641
rect 6822 21632 6828 21684
rect 6880 21632 6886 21684
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7098 21672 7104 21684
rect 6963 21644 7104 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 9214 21672 9220 21684
rect 7708 21644 9220 21672
rect 7708 21632 7714 21644
rect 9214 21632 9220 21644
rect 9272 21672 9278 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9272 21644 9597 21672
rect 9272 21632 9278 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 9677 21675 9735 21681
rect 9677 21641 9689 21675
rect 9723 21641 9735 21675
rect 9677 21635 9735 21641
rect 4522 21564 4528 21616
rect 4580 21604 4586 21616
rect 4982 21604 4988 21616
rect 4580 21576 4988 21604
rect 4580 21564 4586 21576
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 4816 21545 4844 21576
rect 4982 21564 4988 21576
rect 5040 21604 5046 21616
rect 6840 21604 6868 21632
rect 5040 21576 6868 21604
rect 5040 21564 5046 21576
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 5445 21539 5503 21545
rect 5445 21505 5457 21539
rect 5491 21536 5503 21539
rect 5534 21536 5540 21548
rect 5491 21508 5540 21536
rect 5491 21505 5503 21508
rect 5445 21499 5503 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5736 21545 5764 21576
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 9692 21604 9720 21635
rect 9766 21632 9772 21684
rect 9824 21632 9830 21684
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 10594 21672 10600 21684
rect 10183 21644 10600 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 13173 21675 13231 21681
rect 13173 21641 13185 21675
rect 13219 21672 13231 21675
rect 13262 21672 13268 21684
rect 13219 21644 13268 21672
rect 13219 21641 13231 21644
rect 13173 21635 13231 21641
rect 13262 21632 13268 21644
rect 13320 21632 13326 21684
rect 15197 21675 15255 21681
rect 15197 21641 15209 21675
rect 15243 21672 15255 21675
rect 15286 21672 15292 21684
rect 15243 21644 15292 21672
rect 15243 21641 15255 21644
rect 15197 21635 15255 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 17678 21672 17684 21684
rect 17543 21644 17684 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 18506 21672 18512 21684
rect 17788 21644 18512 21672
rect 8260 21576 9720 21604
rect 9784 21604 9812 21632
rect 11974 21604 11980 21616
rect 9784 21576 11980 21604
rect 8260 21564 8266 21576
rect 5721 21539 5779 21545
rect 5721 21505 5733 21539
rect 5767 21505 5779 21539
rect 5721 21499 5779 21505
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 6144 21508 6377 21536
rect 6144 21496 6150 21508
rect 6365 21505 6377 21508
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6546 21496 6552 21548
rect 6604 21496 6610 21548
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 4448 21440 4905 21468
rect 4448 21344 4476 21440
rect 4893 21437 4905 21440
rect 4939 21468 4951 21471
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 4939 21440 5641 21468
rect 4939 21437 4951 21440
rect 4893 21431 4951 21437
rect 5629 21437 5641 21440
rect 5675 21468 5687 21471
rect 6656 21468 6684 21499
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 9398 21496 9404 21548
rect 9456 21496 9462 21548
rect 10331 21545 10359 21576
rect 11974 21564 11980 21576
rect 12032 21564 12038 21616
rect 16758 21564 16764 21616
rect 16816 21564 16822 21616
rect 17788 21604 17816 21644
rect 18506 21632 18512 21644
rect 18564 21632 18570 21684
rect 18598 21632 18604 21684
rect 18656 21632 18662 21684
rect 19058 21632 19064 21684
rect 19116 21632 19122 21684
rect 19705 21675 19763 21681
rect 19705 21641 19717 21675
rect 19751 21672 19763 21675
rect 19978 21672 19984 21684
rect 19751 21644 19984 21672
rect 19751 21641 19763 21644
rect 19705 21635 19763 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 20073 21675 20131 21681
rect 20073 21641 20085 21675
rect 20119 21641 20131 21675
rect 20073 21635 20131 21641
rect 17696 21576 17816 21604
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 10316 21539 10374 21545
rect 9539 21508 9904 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 9876 21480 9904 21508
rect 10316 21505 10328 21539
rect 10362 21505 10374 21539
rect 10316 21499 10374 21505
rect 10410 21496 10416 21548
rect 10468 21496 10474 21548
rect 10502 21496 10508 21548
rect 10560 21496 10566 21548
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 10778 21496 10784 21548
rect 10836 21496 10842 21548
rect 12618 21496 12624 21548
rect 12676 21496 12682 21548
rect 13722 21536 13728 21548
rect 13372 21508 13728 21536
rect 5675 21440 6684 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 9858 21428 9864 21480
rect 9916 21428 9922 21480
rect 9953 21471 10011 21477
rect 9953 21437 9965 21471
rect 9999 21468 10011 21471
rect 10704 21468 10732 21496
rect 12636 21468 12664 21496
rect 9999 21440 12664 21468
rect 9999 21437 10011 21440
rect 9953 21431 10011 21437
rect 11054 21400 11060 21412
rect 6840 21372 11060 21400
rect 6840 21344 6868 21372
rect 11054 21360 11060 21372
rect 11112 21360 11118 21412
rect 13372 21409 13400 21508
rect 13722 21496 13728 21508
rect 13780 21536 13786 21548
rect 14001 21539 14059 21545
rect 14001 21536 14013 21539
rect 13780 21508 14013 21536
rect 13780 21496 13786 21508
rect 14001 21505 14013 21508
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 14884 21508 15393 21536
rect 14884 21496 14890 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16776 21536 16804 21564
rect 17696 21545 17724 21576
rect 17862 21564 17868 21616
rect 17920 21564 17926 21616
rect 18003 21607 18061 21613
rect 18003 21573 18015 21607
rect 18049 21604 18061 21607
rect 18616 21604 18644 21632
rect 18049 21576 18644 21604
rect 19076 21604 19104 21632
rect 20088 21604 20116 21635
rect 21174 21632 21180 21684
rect 21232 21632 21238 21684
rect 22554 21632 22560 21684
rect 22612 21672 22618 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22612 21644 23029 21672
rect 22612 21632 22618 21644
rect 23017 21641 23029 21644
rect 23063 21641 23075 21675
rect 23017 21635 23075 21641
rect 24394 21632 24400 21684
rect 24452 21672 24458 21684
rect 26142 21672 26148 21684
rect 24452 21644 26148 21672
rect 24452 21632 24458 21644
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 19076 21576 20116 21604
rect 18049 21573 18061 21576
rect 18003 21567 18061 21573
rect 20162 21564 20168 21616
rect 20220 21604 20226 21616
rect 20220 21576 21128 21604
rect 20220 21564 20226 21576
rect 16715 21508 16804 21536
rect 17681 21539 17739 21545
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21505 17831 21539
rect 17773 21502 17831 21505
rect 17773 21499 17908 21502
rect 13633 21471 13691 21477
rect 13633 21437 13645 21471
rect 13679 21468 13691 21471
rect 14185 21471 14243 21477
rect 14185 21468 14197 21471
rect 13679 21440 14197 21468
rect 13679 21437 13691 21440
rect 13633 21431 13691 21437
rect 14185 21437 14197 21440
rect 14231 21437 14243 21471
rect 14185 21431 14243 21437
rect 13357 21403 13415 21409
rect 13357 21369 13369 21403
rect 13403 21369 13415 21403
rect 13357 21363 13415 21369
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1489 21335 1547 21341
rect 1489 21332 1501 21335
rect 992 21304 1501 21332
rect 992 21292 998 21304
rect 1489 21301 1501 21304
rect 1535 21301 1547 21335
rect 1489 21295 1547 21301
rect 4430 21292 4436 21344
rect 4488 21292 4494 21344
rect 5074 21292 5080 21344
rect 5132 21292 5138 21344
rect 6822 21292 6828 21344
rect 6880 21292 6886 21344
rect 8113 21335 8171 21341
rect 8113 21301 8125 21335
rect 8159 21332 8171 21335
rect 8478 21332 8484 21344
rect 8159 21304 8484 21332
rect 8159 21301 8171 21304
rect 8113 21295 8171 21301
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 9674 21292 9680 21344
rect 9732 21332 9738 21344
rect 10042 21332 10048 21344
rect 9732 21304 10048 21332
rect 9732 21292 9738 21304
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 13170 21292 13176 21344
rect 13228 21332 13234 21344
rect 13648 21332 13676 21431
rect 14200 21400 14228 21431
rect 15010 21428 15016 21480
rect 15068 21428 15074 21480
rect 15194 21428 15200 21480
rect 15252 21468 15258 21480
rect 15565 21471 15623 21477
rect 17788 21474 17908 21499
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18782 21496 18788 21548
rect 18840 21496 18846 21548
rect 19886 21496 19892 21548
rect 19944 21536 19950 21548
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 19944 21508 20269 21536
rect 19944 21496 19950 21508
rect 20257 21505 20269 21508
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 20346 21496 20352 21548
rect 20404 21496 20410 21548
rect 20533 21539 20591 21545
rect 20533 21536 20545 21539
rect 20456 21508 20545 21536
rect 15565 21468 15577 21471
rect 15252 21440 15577 21468
rect 15252 21428 15258 21440
rect 15565 21437 15577 21440
rect 15611 21437 15623 21471
rect 15565 21431 15623 21437
rect 15212 21400 15240 21428
rect 14200 21372 15240 21400
rect 13228 21304 13676 21332
rect 13817 21335 13875 21341
rect 13228 21292 13234 21304
rect 13817 21301 13829 21335
rect 13863 21332 13875 21335
rect 14274 21332 14280 21344
rect 13863 21304 14280 21332
rect 13863 21301 13875 21304
rect 13817 21295 13875 21301
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 14458 21292 14464 21344
rect 14516 21292 14522 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 16761 21335 16819 21341
rect 16761 21332 16773 21335
rect 16632 21304 16773 21332
rect 16632 21292 16638 21304
rect 16761 21301 16773 21304
rect 16807 21301 16819 21335
rect 17880 21332 17908 21474
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18141 21471 18199 21477
rect 18141 21468 18153 21471
rect 18104 21440 18153 21468
rect 18104 21428 18110 21440
rect 18141 21437 18153 21440
rect 18187 21437 18199 21471
rect 18800 21468 18828 21496
rect 20456 21468 20484 21508
rect 20533 21505 20545 21508
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 20806 21468 20812 21480
rect 18800 21440 20484 21468
rect 20548 21440 20812 21468
rect 18141 21431 18199 21437
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 19334 21400 19340 21412
rect 18380 21372 19340 21400
rect 18380 21360 18386 21372
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 18598 21332 18604 21344
rect 17880 21304 18604 21332
rect 16761 21295 16819 21301
rect 18598 21292 18604 21304
rect 18656 21332 18662 21344
rect 20438 21332 20444 21344
rect 18656 21304 20444 21332
rect 18656 21292 18662 21304
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 20548 21341 20576 21440
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21100 21400 21128 21576
rect 21192 21468 21220 21632
rect 24210 21604 24216 21616
rect 23676 21576 24216 21604
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 22830 21536 22836 21548
rect 21600 21508 22836 21536
rect 21600 21496 21606 21508
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21536 22983 21539
rect 23014 21536 23020 21548
rect 22971 21508 23020 21536
rect 22971 21505 22983 21508
rect 22925 21499 22983 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23676 21545 23704 21576
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 26786 21564 26792 21616
rect 26844 21604 26850 21616
rect 27801 21607 27859 21613
rect 27801 21604 27813 21607
rect 26844 21576 27813 21604
rect 26844 21564 26850 21576
rect 27801 21573 27813 21576
rect 27847 21573 27859 21607
rect 27801 21567 27859 21573
rect 27982 21564 27988 21616
rect 28040 21564 28046 21616
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21505 23719 21539
rect 23661 21499 23719 21505
rect 25056 21508 25636 21536
rect 21453 21471 21511 21477
rect 21453 21468 21465 21471
rect 21192 21440 21465 21468
rect 21453 21437 21465 21440
rect 21499 21468 21511 21471
rect 22278 21468 22284 21480
rect 21499 21440 22284 21468
rect 21499 21437 21511 21440
rect 21453 21431 21511 21437
rect 22278 21428 22284 21440
rect 22336 21428 22342 21480
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 24026 21428 24032 21480
rect 24084 21468 24090 21480
rect 25056 21468 25084 21508
rect 24084 21440 25084 21468
rect 24084 21428 24090 21440
rect 25314 21428 25320 21480
rect 25372 21468 25378 21480
rect 25608 21477 25636 21508
rect 25866 21496 25872 21548
rect 25924 21496 25930 21548
rect 26418 21496 26424 21548
rect 26476 21536 26482 21548
rect 26970 21536 26976 21548
rect 26476 21508 26976 21536
rect 26476 21496 26482 21508
rect 26970 21496 26976 21508
rect 27028 21496 27034 21548
rect 27338 21496 27344 21548
rect 27396 21536 27402 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 27396 21508 27445 21536
rect 27396 21496 27402 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21536 27675 21539
rect 28000 21536 28028 21564
rect 27663 21508 28028 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 25501 21471 25559 21477
rect 25501 21468 25513 21471
rect 25372 21440 25513 21468
rect 25372 21428 25378 21440
rect 25501 21437 25513 21440
rect 25547 21437 25559 21471
rect 25501 21431 25559 21437
rect 25593 21471 25651 21477
rect 25593 21437 25605 21471
rect 25639 21437 25651 21471
rect 26878 21468 26884 21480
rect 25593 21431 25651 21437
rect 26252 21440 26884 21468
rect 21100 21372 21404 21400
rect 20533 21335 20591 21341
rect 20533 21301 20545 21335
rect 20579 21301 20591 21335
rect 20533 21295 20591 21301
rect 20622 21292 20628 21344
rect 20680 21332 20686 21344
rect 21376 21341 21404 21372
rect 21177 21335 21235 21341
rect 21177 21332 21189 21335
rect 20680 21304 21189 21332
rect 20680 21292 20686 21304
rect 21177 21301 21189 21304
rect 21223 21301 21235 21335
rect 21177 21295 21235 21301
rect 21361 21335 21419 21341
rect 21361 21301 21373 21335
rect 21407 21301 21419 21335
rect 25516 21332 25544 21431
rect 26252 21332 26280 21440
rect 26878 21428 26884 21440
rect 26936 21428 26942 21480
rect 27249 21471 27307 21477
rect 27249 21437 27261 21471
rect 27295 21468 27307 21471
rect 27632 21468 27660 21499
rect 27295 21440 27660 21468
rect 27295 21437 27307 21440
rect 27249 21431 27307 21437
rect 26602 21360 26608 21412
rect 26660 21400 26666 21412
rect 27264 21400 27292 21431
rect 26660 21372 27292 21400
rect 26660 21360 26666 21372
rect 25516 21304 26280 21332
rect 21361 21295 21419 21301
rect 26970 21292 26976 21344
rect 27028 21292 27034 21344
rect 27246 21292 27252 21344
rect 27304 21292 27310 21344
rect 1104 21242 30820 21264
rect 1104 21190 4664 21242
rect 4716 21190 4728 21242
rect 4780 21190 4792 21242
rect 4844 21190 4856 21242
rect 4908 21190 4920 21242
rect 4972 21190 12092 21242
rect 12144 21190 12156 21242
rect 12208 21190 12220 21242
rect 12272 21190 12284 21242
rect 12336 21190 12348 21242
rect 12400 21190 19520 21242
rect 19572 21190 19584 21242
rect 19636 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 26948 21242
rect 27000 21190 27012 21242
rect 27064 21190 27076 21242
rect 27128 21190 27140 21242
rect 27192 21190 27204 21242
rect 27256 21190 30820 21242
rect 1104 21168 30820 21190
rect 5074 21088 5080 21140
rect 5132 21088 5138 21140
rect 5721 21131 5779 21137
rect 5721 21097 5733 21131
rect 5767 21128 5779 21131
rect 6546 21128 6552 21140
rect 5767 21100 6552 21128
rect 5767 21097 5779 21100
rect 5721 21091 5779 21097
rect 6546 21088 6552 21100
rect 6604 21088 6610 21140
rect 8021 21131 8079 21137
rect 8021 21097 8033 21131
rect 8067 21128 8079 21131
rect 8570 21128 8576 21140
rect 8067 21100 8576 21128
rect 8067 21097 8079 21100
rect 8021 21091 8079 21097
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 9490 21088 9496 21140
rect 9548 21088 9554 21140
rect 9674 21088 9680 21140
rect 9732 21088 9738 21140
rect 9950 21128 9956 21140
rect 9784 21100 9956 21128
rect 5092 20992 5120 21088
rect 6086 21020 6092 21072
rect 6144 21060 6150 21072
rect 6822 21060 6828 21072
rect 6144 21032 6828 21060
rect 6144 21020 6150 21032
rect 6822 21020 6828 21032
rect 6880 21020 6886 21072
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21029 6975 21063
rect 9217 21063 9275 21069
rect 9217 21060 9229 21063
rect 6917 21023 6975 21029
rect 7484 21032 9229 21060
rect 5353 20995 5411 21001
rect 5353 20992 5365 20995
rect 5092 20964 5365 20992
rect 5353 20961 5365 20964
rect 5399 20961 5411 20995
rect 6932 20992 6960 21023
rect 5353 20955 5411 20961
rect 6012 20964 6960 20992
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 4154 20924 4160 20936
rect 1719 20896 4160 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 4246 20884 4252 20936
rect 4304 20924 4310 20936
rect 5074 20924 5080 20936
rect 4304 20896 5080 20924
rect 4304 20884 4310 20896
rect 5074 20884 5080 20896
rect 5132 20884 5138 20936
rect 5534 20933 5540 20936
rect 5523 20927 5540 20933
rect 5523 20893 5535 20927
rect 5592 20924 5598 20936
rect 6012 20924 6040 20964
rect 7006 20952 7012 21004
rect 7064 20952 7070 21004
rect 5592 20896 6040 20924
rect 5523 20887 5540 20893
rect 5534 20884 5540 20887
rect 5592 20884 5598 20896
rect 6454 20884 6460 20936
rect 6512 20884 6518 20936
rect 6641 20927 6699 20933
rect 6641 20893 6653 20927
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 6650 20856 6678 20887
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 7484 20933 7512 21032
rect 9217 21029 9229 21032
rect 9263 21029 9275 21063
rect 9217 21023 9275 21029
rect 7558 20952 7564 21004
rect 7616 20952 7622 21004
rect 7837 20995 7895 21001
rect 7837 20961 7849 20995
rect 7883 20961 7895 20995
rect 9508 20992 9536 21088
rect 7837 20955 7895 20961
rect 8404 20964 9536 20992
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7469 20927 7527 20933
rect 7469 20924 7481 20927
rect 6871 20896 7481 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 7469 20893 7481 20896
rect 7515 20893 7527 20927
rect 7852 20924 7880 20955
rect 8404 20933 8432 20964
rect 9674 20952 9680 21004
rect 9732 20992 9738 21004
rect 9784 20992 9812 21100
rect 9950 21088 9956 21100
rect 10008 21128 10014 21140
rect 10008 21100 10456 21128
rect 10008 21088 10014 21100
rect 10428 21072 10456 21100
rect 10502 21088 10508 21140
rect 10560 21088 10566 21140
rect 10689 21131 10747 21137
rect 10689 21097 10701 21131
rect 10735 21128 10747 21131
rect 10778 21128 10784 21140
rect 10735 21100 10784 21128
rect 10735 21097 10747 21100
rect 10689 21091 10747 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11974 21088 11980 21140
rect 12032 21088 12038 21140
rect 12161 21131 12219 21137
rect 12161 21097 12173 21131
rect 12207 21128 12219 21131
rect 12434 21128 12440 21140
rect 12207 21100 12440 21128
rect 12207 21097 12219 21100
rect 12161 21091 12219 21097
rect 12434 21088 12440 21100
rect 12492 21128 12498 21140
rect 12805 21131 12863 21137
rect 12805 21128 12817 21131
rect 12492 21100 12817 21128
rect 12492 21088 12498 21100
rect 12805 21097 12817 21100
rect 12851 21097 12863 21131
rect 12805 21091 12863 21097
rect 14829 21131 14887 21137
rect 14829 21097 14841 21131
rect 14875 21128 14887 21131
rect 15010 21128 15016 21140
rect 14875 21100 15016 21128
rect 14875 21097 14887 21100
rect 14829 21091 14887 21097
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 16390 21128 16396 21140
rect 15580 21100 16396 21128
rect 9858 21020 9864 21072
rect 9916 21060 9922 21072
rect 10229 21063 10287 21069
rect 9916 21032 10180 21060
rect 9916 21020 9922 21032
rect 9732 20964 9996 20992
rect 9732 20952 9738 20964
rect 9968 20933 9996 20964
rect 8205 20927 8263 20933
rect 8205 20924 8217 20927
rect 7852 20896 8217 20924
rect 7469 20887 7527 20893
rect 8205 20893 8217 20896
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 8389 20927 8447 20933
rect 8389 20893 8401 20927
rect 8435 20893 8447 20927
rect 8573 20927 8631 20933
rect 8573 20924 8585 20927
rect 8389 20887 8447 20893
rect 8496 20896 8585 20924
rect 6650 20828 6776 20856
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 4522 20748 4528 20800
rect 4580 20748 4586 20800
rect 6549 20791 6607 20797
rect 6549 20757 6561 20791
rect 6595 20788 6607 20791
rect 6638 20788 6644 20800
rect 6595 20760 6644 20788
rect 6595 20757 6607 20760
rect 6549 20751 6607 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 6748 20788 6776 20828
rect 6914 20816 6920 20868
rect 6972 20856 6978 20868
rect 8297 20859 8355 20865
rect 8297 20856 8309 20859
rect 6972 20828 8309 20856
rect 6972 20816 6978 20828
rect 8297 20825 8309 20828
rect 8343 20825 8355 20859
rect 8297 20819 8355 20825
rect 7650 20788 7656 20800
rect 6748 20760 7656 20788
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 8496 20788 8524 20896
rect 8573 20893 8585 20896
rect 8619 20893 8631 20927
rect 8573 20887 8631 20893
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 9953 20927 10011 20933
rect 9447 20896 9904 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 8260 20760 8524 20788
rect 8956 20788 8984 20887
rect 9876 20868 9904 20896
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 10042 20884 10048 20936
rect 10100 20884 10106 20936
rect 10152 20924 10180 21032
rect 10229 21029 10241 21063
rect 10275 21029 10287 21063
rect 10229 21023 10287 21029
rect 10244 20992 10272 21023
rect 10410 21020 10416 21072
rect 10468 21020 10474 21072
rect 12618 21020 12624 21072
rect 12676 21020 12682 21072
rect 15580 21004 15608 21100
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 19426 21088 19432 21140
rect 19484 21088 19490 21140
rect 20346 21088 20352 21140
rect 20404 21128 20410 21140
rect 20404 21100 23060 21128
rect 20404 21088 20410 21100
rect 23032 21072 23060 21100
rect 23106 21088 23112 21140
rect 23164 21128 23170 21140
rect 23569 21131 23627 21137
rect 23569 21128 23581 21131
rect 23164 21100 23581 21128
rect 23164 21088 23170 21100
rect 23569 21097 23581 21100
rect 23615 21097 23627 21131
rect 23569 21091 23627 21097
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 26694 21128 26700 21140
rect 23799 21100 26700 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 18690 21020 18696 21072
rect 18748 21020 18754 21072
rect 19536 21032 20852 21060
rect 10244 20964 10548 20992
rect 10520 20933 10548 20964
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 11333 20995 11391 21001
rect 11333 20992 11345 20995
rect 11020 20964 11345 20992
rect 11020 20952 11026 20964
rect 11333 20961 11345 20964
rect 11379 20961 11391 20995
rect 11333 20955 11391 20961
rect 14185 20995 14243 21001
rect 14185 20961 14197 20995
rect 14231 20992 14243 20995
rect 14231 20964 15332 20992
rect 14231 20961 14243 20964
rect 14185 20955 14243 20961
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 10152 20896 10333 20924
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 10505 20927 10563 20933
rect 10505 20893 10517 20927
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20924 10931 20927
rect 11514 20924 11520 20936
rect 10919 20896 11520 20924
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11514 20884 11520 20896
rect 11572 20884 11578 20936
rect 11790 20884 11796 20936
rect 11848 20884 11854 20936
rect 12529 20927 12587 20933
rect 12529 20893 12541 20927
rect 12575 20924 12587 20927
rect 13078 20924 13084 20936
rect 12575 20896 13084 20924
rect 12575 20893 12587 20896
rect 12529 20887 12587 20893
rect 13078 20884 13084 20896
rect 13136 20924 13142 20936
rect 13173 20927 13231 20933
rect 13173 20924 13185 20927
rect 13136 20896 13185 20924
rect 13136 20884 13142 20896
rect 13173 20893 13185 20896
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 9033 20859 9091 20865
rect 9033 20825 9045 20859
rect 9079 20856 9091 20859
rect 9306 20856 9312 20868
rect 9079 20828 9312 20856
rect 9079 20825 9091 20828
rect 9033 20819 9091 20825
rect 9306 20816 9312 20828
rect 9364 20856 9370 20868
rect 9493 20859 9551 20865
rect 9493 20856 9505 20859
rect 9364 20828 9505 20856
rect 9364 20816 9370 20828
rect 9493 20825 9505 20828
rect 9539 20856 9551 20859
rect 9539 20828 9812 20856
rect 9539 20825 9551 20828
rect 9493 20819 9551 20825
rect 9582 20788 9588 20800
rect 8956 20760 9588 20788
rect 8260 20748 8266 20760
rect 9582 20748 9588 20760
rect 9640 20748 9646 20800
rect 9674 20748 9680 20800
rect 9732 20797 9738 20800
rect 9732 20791 9751 20797
rect 9739 20757 9751 20791
rect 9784 20788 9812 20828
rect 9858 20816 9864 20868
rect 9916 20816 9922 20868
rect 10134 20856 10140 20868
rect 9968 20828 10140 20856
rect 9968 20788 9996 20828
rect 10134 20816 10140 20828
rect 10192 20856 10198 20868
rect 10229 20859 10287 20865
rect 10229 20856 10241 20859
rect 10192 20828 10241 20856
rect 10192 20816 10198 20828
rect 10229 20825 10241 20828
rect 10275 20825 10287 20859
rect 10229 20819 10287 20825
rect 10962 20816 10968 20868
rect 11020 20816 11026 20868
rect 11054 20816 11060 20868
rect 11112 20816 11118 20868
rect 11146 20816 11152 20868
rect 11204 20865 11210 20868
rect 11204 20859 11233 20865
rect 11221 20825 11233 20859
rect 11204 20819 11233 20825
rect 11204 20816 11210 20819
rect 11606 20816 11612 20868
rect 11664 20816 11670 20868
rect 12434 20816 12440 20868
rect 12492 20856 12498 20868
rect 12805 20859 12863 20865
rect 12805 20856 12817 20859
rect 12492 20828 12817 20856
rect 12492 20816 12498 20828
rect 12805 20825 12817 20828
rect 12851 20856 12863 20859
rect 14200 20856 14228 20955
rect 15304 20936 15332 20964
rect 15562 20952 15568 21004
rect 15620 20952 15626 21004
rect 15654 20952 15660 21004
rect 15712 20992 15718 21004
rect 16666 20992 16672 21004
rect 15712 20964 16672 20992
rect 15712 20952 15718 20964
rect 16666 20952 16672 20964
rect 16724 20952 16730 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 18892 20964 19257 20992
rect 18892 20936 18920 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20924 14703 20927
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14691 20896 14933 20924
rect 14691 20893 14703 20896
rect 14645 20887 14703 20893
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 15286 20884 15292 20936
rect 15344 20884 15350 20936
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 12851 20828 14228 20856
rect 12851 20825 12863 20828
rect 12805 20819 12863 20825
rect 14274 20816 14280 20868
rect 14332 20856 14338 20868
rect 14332 20828 15056 20856
rect 14332 20816 14338 20828
rect 9784 20760 9996 20788
rect 10980 20788 11008 20816
rect 15028 20800 15056 20828
rect 15930 20816 15936 20868
rect 15988 20816 15994 20868
rect 16574 20816 16580 20868
rect 16632 20816 16638 20868
rect 17681 20859 17739 20865
rect 17681 20825 17693 20859
rect 17727 20825 17739 20859
rect 18616 20856 18644 20887
rect 18782 20884 18788 20936
rect 18840 20884 18846 20936
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 19061 20927 19119 20933
rect 19061 20893 19073 20927
rect 19107 20924 19119 20927
rect 19334 20924 19340 20936
rect 19107 20896 19340 20924
rect 19107 20893 19119 20896
rect 19061 20887 19119 20893
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 18966 20856 18972 20868
rect 18616 20828 18972 20856
rect 17681 20819 17739 20825
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 10980 20760 11437 20788
rect 9732 20751 9751 20757
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 9732 20748 9738 20751
rect 12066 20748 12072 20800
rect 12124 20788 12130 20800
rect 12161 20791 12219 20797
rect 12161 20788 12173 20791
rect 12124 20760 12173 20788
rect 12124 20748 12130 20760
rect 12161 20757 12173 20760
rect 12207 20757 12219 20791
rect 12161 20751 12219 20757
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 14182 20788 14188 20800
rect 13780 20760 14188 20788
rect 13780 20748 13786 20760
rect 14182 20748 14188 20760
rect 14240 20788 14246 20800
rect 14369 20791 14427 20797
rect 14369 20788 14381 20791
rect 14240 20760 14381 20788
rect 14240 20748 14246 20760
rect 14369 20757 14381 20760
rect 14415 20757 14427 20791
rect 14369 20751 14427 20757
rect 15010 20748 15016 20800
rect 15068 20748 15074 20800
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 17696 20788 17724 20819
rect 18966 20816 18972 20828
rect 19024 20856 19030 20868
rect 19536 20856 19564 21032
rect 20824 21004 20852 21032
rect 22278 21020 22284 21072
rect 22336 21060 22342 21072
rect 22830 21060 22836 21072
rect 22336 21032 22836 21060
rect 22336 21020 22342 21032
rect 22830 21020 22836 21032
rect 22888 21020 22894 21072
rect 23014 21020 23020 21072
rect 23072 21020 23078 21072
rect 23768 21060 23796 21091
rect 26694 21088 26700 21100
rect 26752 21088 26758 21140
rect 26786 21088 26792 21140
rect 26844 21128 26850 21140
rect 27249 21131 27307 21137
rect 27249 21128 27261 21131
rect 26844 21100 27261 21128
rect 26844 21088 26850 21100
rect 27249 21097 27261 21100
rect 27295 21097 27307 21131
rect 27249 21091 27307 21097
rect 27522 21088 27528 21140
rect 27580 21128 27586 21140
rect 28077 21131 28135 21137
rect 28077 21128 28089 21131
rect 27580 21100 28089 21128
rect 27580 21088 27586 21100
rect 28077 21097 28089 21100
rect 28123 21097 28135 21131
rect 28077 21091 28135 21097
rect 27433 21063 27491 21069
rect 23308 21032 23796 21060
rect 23860 21032 27384 21060
rect 19610 20952 19616 21004
rect 19668 20992 19674 21004
rect 19797 20995 19855 21001
rect 19797 20992 19809 20995
rect 19668 20964 19809 20992
rect 19668 20952 19674 20964
rect 19797 20961 19809 20964
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 20714 20952 20720 21004
rect 20772 20952 20778 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 20864 20964 22232 20992
rect 20864 20952 20870 20964
rect 22204 20936 22232 20964
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19024 20828 19564 20856
rect 19720 20856 19748 20887
rect 22186 20884 22192 20936
rect 22244 20924 22250 20936
rect 23308 20933 23336 21032
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20992 23535 20995
rect 23860 20992 23888 21032
rect 24857 20995 24915 21001
rect 23523 20964 24072 20992
rect 23523 20961 23535 20964
rect 23477 20955 23535 20961
rect 22649 20927 22707 20933
rect 22649 20924 22661 20927
rect 22244 20896 22661 20924
rect 22244 20884 22250 20896
rect 22649 20893 22661 20896
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 22925 20927 22983 20933
rect 22925 20893 22937 20927
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23293 20927 23351 20933
rect 23293 20893 23305 20927
rect 23339 20893 23351 20927
rect 23293 20887 23351 20893
rect 19981 20859 20039 20865
rect 19720 20828 19932 20856
rect 19024 20816 19030 20828
rect 19904 20800 19932 20828
rect 19981 20825 19993 20859
rect 20027 20825 20039 20859
rect 19981 20819 20039 20825
rect 16816 20760 17724 20788
rect 16816 20748 16822 20760
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 18417 20791 18475 20797
rect 18417 20788 18429 20791
rect 18012 20760 18429 20788
rect 18012 20748 18018 20760
rect 18417 20757 18429 20760
rect 18463 20757 18475 20791
rect 18417 20751 18475 20757
rect 19886 20748 19892 20800
rect 19944 20748 19950 20800
rect 19996 20788 20024 20819
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 21910 20856 21916 20868
rect 21048 20828 21916 20856
rect 21048 20816 21054 20828
rect 21910 20816 21916 20828
rect 21968 20816 21974 20868
rect 22465 20859 22523 20865
rect 22465 20825 22477 20859
rect 22511 20825 22523 20859
rect 22465 20819 22523 20825
rect 22833 20859 22891 20865
rect 22833 20825 22845 20859
rect 22879 20856 22891 20859
rect 22940 20856 22968 20887
rect 23937 20859 23995 20865
rect 23937 20856 23949 20859
rect 22879 20828 23949 20856
rect 22879 20825 22891 20828
rect 22833 20819 22891 20825
rect 23937 20825 23949 20828
rect 23983 20825 23995 20859
rect 23937 20819 23995 20825
rect 20070 20788 20076 20800
rect 19996 20760 20076 20788
rect 20070 20748 20076 20760
rect 20128 20748 20134 20800
rect 22373 20791 22431 20797
rect 22373 20757 22385 20791
rect 22419 20788 22431 20791
rect 22480 20788 22508 20819
rect 22419 20760 22508 20788
rect 23737 20791 23795 20797
rect 22419 20757 22431 20760
rect 22373 20751 22431 20757
rect 23737 20757 23749 20791
rect 23783 20788 23795 20791
rect 24044 20788 24072 20964
rect 24857 20961 24869 20995
rect 24903 20992 24915 20995
rect 25498 20992 25504 21004
rect 24903 20964 25504 20992
rect 24903 20961 24915 20964
rect 24857 20955 24915 20961
rect 25498 20952 25504 20964
rect 25556 20952 25562 21004
rect 26602 20952 26608 21004
rect 26660 20952 26666 21004
rect 26697 20995 26755 21001
rect 26697 20961 26709 20995
rect 26743 20992 26755 20995
rect 27154 20992 27160 21004
rect 26743 20964 27160 20992
rect 26743 20961 26755 20964
rect 26697 20955 26755 20961
rect 27154 20952 27160 20964
rect 27212 20952 27218 21004
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 25041 20859 25099 20865
rect 25041 20856 25053 20859
rect 24176 20828 25053 20856
rect 24176 20816 24182 20828
rect 25041 20825 25053 20828
rect 25087 20825 25099 20859
rect 26620 20856 26648 20952
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 26973 20927 27031 20933
rect 26973 20893 26985 20927
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 26988 20856 27016 20887
rect 26620 20828 27016 20856
rect 27065 20859 27123 20865
rect 25041 20819 25099 20825
rect 27065 20825 27077 20859
rect 27111 20856 27123 20859
rect 27154 20856 27160 20868
rect 27111 20828 27160 20856
rect 27111 20825 27123 20828
rect 27065 20819 27123 20825
rect 27154 20816 27160 20828
rect 27212 20816 27218 20868
rect 27356 20856 27384 21032
rect 27433 21029 27445 21063
rect 27479 21060 27491 21063
rect 27982 21060 27988 21072
rect 27479 21032 27660 21060
rect 27479 21029 27491 21032
rect 27433 21023 27491 21029
rect 27632 21001 27660 21032
rect 27724 21032 27988 21060
rect 27724 21001 27752 21032
rect 27982 21020 27988 21032
rect 28040 21020 28046 21072
rect 28626 21020 28632 21072
rect 28684 21020 28690 21072
rect 27617 20995 27675 21001
rect 27617 20961 27629 20995
rect 27663 20961 27675 20995
rect 27617 20955 27675 20961
rect 27709 20995 27767 21001
rect 27709 20961 27721 20995
rect 27755 20961 27767 20995
rect 27709 20955 27767 20961
rect 27801 20995 27859 21001
rect 27801 20961 27813 20995
rect 27847 20992 27859 20995
rect 28644 20992 28672 21020
rect 27847 20964 28672 20992
rect 27847 20961 27859 20964
rect 27801 20955 27859 20961
rect 27893 20927 27951 20933
rect 27893 20893 27905 20927
rect 27939 20924 27951 20927
rect 28353 20927 28411 20933
rect 27939 20896 28304 20924
rect 27939 20893 27951 20896
rect 27893 20887 27951 20893
rect 28169 20859 28227 20865
rect 28169 20856 28181 20859
rect 27356 20828 28181 20856
rect 28169 20825 28181 20828
rect 28215 20825 28227 20859
rect 28169 20819 28227 20825
rect 23783 20760 24072 20788
rect 26973 20791 27031 20797
rect 23783 20757 23795 20760
rect 23737 20751 23795 20757
rect 26973 20757 26985 20791
rect 27019 20788 27031 20791
rect 27265 20791 27323 20797
rect 27265 20788 27277 20791
rect 27019 20760 27277 20788
rect 27019 20757 27031 20760
rect 26973 20751 27031 20757
rect 27265 20757 27277 20760
rect 27311 20757 27323 20791
rect 28276 20788 28304 20896
rect 28353 20893 28365 20927
rect 28399 20924 28411 20927
rect 28442 20924 28448 20936
rect 28399 20896 28448 20924
rect 28399 20893 28411 20896
rect 28353 20887 28411 20893
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28534 20884 28540 20936
rect 28592 20884 28598 20936
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20924 28687 20927
rect 29362 20924 29368 20936
rect 28675 20896 29368 20924
rect 28675 20893 28687 20896
rect 28629 20887 28687 20893
rect 29362 20884 29368 20896
rect 29420 20884 29426 20936
rect 29638 20788 29644 20800
rect 28276 20760 29644 20788
rect 27265 20751 27323 20757
rect 29638 20748 29644 20760
rect 29696 20748 29702 20800
rect 1104 20698 30820 20720
rect 1104 20646 5324 20698
rect 5376 20646 5388 20698
rect 5440 20646 5452 20698
rect 5504 20646 5516 20698
rect 5568 20646 5580 20698
rect 5632 20646 12752 20698
rect 12804 20646 12816 20698
rect 12868 20646 12880 20698
rect 12932 20646 12944 20698
rect 12996 20646 13008 20698
rect 13060 20646 20180 20698
rect 20232 20646 20244 20698
rect 20296 20646 20308 20698
rect 20360 20646 20372 20698
rect 20424 20646 20436 20698
rect 20488 20646 27608 20698
rect 27660 20646 27672 20698
rect 27724 20646 27736 20698
rect 27788 20646 27800 20698
rect 27852 20646 27864 20698
rect 27916 20646 30820 20698
rect 1104 20624 30820 20646
rect 4246 20544 4252 20596
rect 4304 20544 4310 20596
rect 4522 20544 4528 20596
rect 4580 20584 4586 20596
rect 4709 20587 4767 20593
rect 4709 20584 4721 20587
rect 4580 20556 4721 20584
rect 4580 20544 4586 20556
rect 4709 20553 4721 20556
rect 4755 20553 4767 20587
rect 4709 20547 4767 20553
rect 5074 20544 5080 20596
rect 5132 20584 5138 20596
rect 5132 20556 5764 20584
rect 5132 20544 5138 20556
rect 4614 20516 4620 20528
rect 4264 20488 4620 20516
rect 4264 20460 4292 20488
rect 4614 20476 4620 20488
rect 4672 20516 4678 20528
rect 4801 20519 4859 20525
rect 4801 20516 4813 20519
rect 4672 20488 4813 20516
rect 4672 20476 4678 20488
rect 4801 20485 4813 20488
rect 4847 20485 4859 20519
rect 4801 20479 4859 20485
rect 5166 20476 5172 20528
rect 5224 20516 5230 20528
rect 5445 20519 5503 20525
rect 5445 20516 5457 20519
rect 5224 20488 5457 20516
rect 5224 20476 5230 20488
rect 5445 20485 5457 20488
rect 5491 20485 5503 20519
rect 5445 20479 5503 20485
rect 3878 20408 3884 20460
rect 3936 20408 3942 20460
rect 4246 20408 4252 20460
rect 4304 20408 4310 20460
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 2498 20340 2504 20392
rect 2556 20340 2562 20392
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 4154 20340 4160 20392
rect 4212 20340 4218 20392
rect 4985 20383 5043 20389
rect 4985 20349 4997 20383
rect 5031 20380 5043 20383
rect 5074 20380 5080 20392
rect 5031 20352 5080 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 4172 20312 4200 20340
rect 5169 20315 5227 20321
rect 5169 20312 5181 20315
rect 4172 20284 5181 20312
rect 5169 20281 5181 20284
rect 5215 20281 5227 20315
rect 5169 20275 5227 20281
rect 5368 20256 5396 20411
rect 5534 20408 5540 20460
rect 5592 20408 5598 20460
rect 5736 20457 5764 20556
rect 7006 20544 7012 20596
rect 7064 20544 7070 20596
rect 7558 20544 7564 20596
rect 7616 20544 7622 20596
rect 9858 20544 9864 20596
rect 9916 20584 9922 20596
rect 10962 20584 10968 20596
rect 9916 20556 10968 20584
rect 9916 20544 9922 20556
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 11514 20544 11520 20596
rect 11572 20544 11578 20596
rect 11790 20544 11796 20596
rect 11848 20544 11854 20596
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 12069 20587 12127 20593
rect 12069 20584 12081 20587
rect 11940 20556 12081 20584
rect 11940 20544 11946 20556
rect 12069 20553 12081 20556
rect 12115 20553 12127 20587
rect 12434 20584 12440 20596
rect 12069 20547 12127 20553
rect 12176 20556 12440 20584
rect 7024 20516 7052 20544
rect 7745 20519 7803 20525
rect 7745 20516 7757 20519
rect 7024 20488 7757 20516
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20417 5779 20451
rect 5721 20411 5779 20417
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 7576 20457 7604 20488
rect 7745 20485 7757 20488
rect 7791 20485 7803 20519
rect 8754 20516 8760 20528
rect 7745 20479 7803 20485
rect 7852 20488 8760 20516
rect 6917 20451 6975 20457
rect 6917 20448 6929 20451
rect 6512 20420 6929 20448
rect 6512 20408 6518 20420
rect 6917 20417 6929 20420
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7285 20451 7343 20457
rect 7285 20417 7297 20451
rect 7331 20448 7343 20451
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 7331 20420 7389 20448
rect 7331 20417 7343 20420
rect 7285 20411 7343 20417
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20417 7619 20451
rect 7561 20411 7619 20417
rect 6932 20312 6960 20411
rect 7116 20380 7144 20411
rect 7650 20408 7656 20460
rect 7708 20408 7714 20460
rect 7852 20457 7880 20488
rect 8754 20476 8760 20488
rect 8812 20476 8818 20528
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20417 7895 20451
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 7837 20411 7895 20417
rect 11072 20420 11529 20448
rect 7668 20380 7696 20408
rect 7116 20352 7696 20380
rect 7852 20312 7880 20411
rect 11072 20324 11100 20420
rect 11517 20417 11529 20420
rect 11563 20448 11575 20451
rect 11606 20448 11612 20460
rect 11563 20420 11612 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 11808 20448 11836 20544
rect 11747 20420 11836 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11238 20340 11244 20392
rect 11296 20340 11302 20392
rect 6932 20284 7880 20312
rect 11054 20272 11060 20324
rect 11112 20272 11118 20324
rect 4338 20204 4344 20256
rect 4396 20204 4402 20256
rect 5350 20204 5356 20256
rect 5408 20244 5414 20256
rect 8018 20244 8024 20256
rect 5408 20216 8024 20244
rect 5408 20204 5414 20216
rect 8018 20204 8024 20216
rect 8076 20204 8082 20256
rect 11256 20244 11284 20340
rect 11900 20312 11928 20544
rect 11977 20451 12035 20457
rect 11977 20417 11989 20451
rect 12023 20448 12035 20451
rect 12066 20448 12072 20460
rect 12023 20420 12072 20448
rect 12023 20417 12035 20420
rect 11977 20411 12035 20417
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12176 20457 12204 20556
rect 12434 20544 12440 20556
rect 12492 20544 12498 20596
rect 13078 20584 13084 20596
rect 12636 20556 13084 20584
rect 12636 20525 12664 20556
rect 13078 20544 13084 20556
rect 13136 20584 13142 20596
rect 13722 20584 13728 20596
rect 13136 20556 13728 20584
rect 13136 20544 13142 20556
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 15654 20584 15660 20596
rect 13924 20556 15660 20584
rect 12621 20519 12679 20525
rect 12391 20485 12449 20491
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12391 20451 12403 20485
rect 12437 20460 12449 20485
rect 12621 20485 12633 20519
rect 12667 20485 12679 20519
rect 12621 20479 12679 20485
rect 12989 20519 13047 20525
rect 12989 20485 13001 20519
rect 13035 20516 13047 20519
rect 13035 20488 13768 20516
rect 13035 20485 13047 20488
rect 12989 20479 13047 20485
rect 12437 20451 12440 20460
rect 12391 20448 12440 20451
rect 12161 20411 12219 20417
rect 12268 20420 12440 20448
rect 12084 20380 12112 20408
rect 12268 20380 12296 20420
rect 12434 20408 12440 20420
rect 12492 20448 12498 20460
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12492 20420 12909 20448
rect 12492 20408 12498 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20417 13139 20451
rect 13081 20411 13139 20417
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13096 20380 13124 20411
rect 12084 20352 12296 20380
rect 12406 20352 13124 20380
rect 12406 20312 12434 20352
rect 11900 20284 12434 20312
rect 13280 20312 13308 20411
rect 13740 20380 13768 20488
rect 13814 20408 13820 20460
rect 13872 20408 13878 20460
rect 13924 20457 13952 20556
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 15930 20544 15936 20596
rect 15988 20584 15994 20596
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 15988 20556 16221 20584
rect 15988 20544 15994 20556
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 16209 20547 16267 20553
rect 16669 20587 16727 20593
rect 16669 20553 16681 20587
rect 16715 20553 16727 20587
rect 16669 20547 16727 20553
rect 14185 20519 14243 20525
rect 14185 20485 14197 20519
rect 14231 20516 14243 20519
rect 14458 20516 14464 20528
rect 14231 20488 14464 20516
rect 14231 20485 14243 20488
rect 14185 20479 14243 20485
rect 14458 20476 14464 20488
rect 14516 20476 14522 20528
rect 15841 20519 15899 20525
rect 15841 20516 15853 20519
rect 15410 20488 15853 20516
rect 15841 20485 15853 20488
rect 15887 20485 15899 20519
rect 15841 20479 15899 20485
rect 16022 20476 16028 20528
rect 16080 20476 16086 20528
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 15562 20408 15568 20460
rect 15620 20408 15626 20460
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 16040 20448 16068 20476
rect 15795 20420 16068 20448
rect 16393 20451 16451 20457
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 16393 20417 16405 20451
rect 16439 20448 16451 20451
rect 16684 20448 16712 20547
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 20036 20556 20085 20584
rect 20036 20544 20042 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20073 20547 20131 20553
rect 20714 20544 20720 20596
rect 20772 20544 20778 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22094 20584 22100 20596
rect 21876 20556 22100 20584
rect 21876 20544 21882 20556
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 22830 20544 22836 20596
rect 22888 20544 22894 20596
rect 26786 20544 26792 20596
rect 26844 20584 26850 20596
rect 27338 20584 27344 20596
rect 26844 20556 27344 20584
rect 26844 20544 26850 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 28537 20587 28595 20593
rect 28537 20553 28549 20587
rect 28583 20584 28595 20587
rect 28626 20584 28632 20596
rect 28583 20556 28632 20584
rect 28583 20553 28595 20556
rect 28537 20547 28595 20553
rect 28626 20544 28632 20556
rect 28684 20544 28690 20596
rect 28810 20544 28816 20596
rect 28868 20544 28874 20596
rect 28920 20556 29316 20584
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 19392 20488 19441 20516
rect 19392 20476 19398 20488
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 19429 20479 19487 20485
rect 16439 20420 16712 20448
rect 16439 20417 16451 20420
rect 16393 20411 16451 20417
rect 14274 20380 14280 20392
rect 13740 20352 14280 20380
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 15580 20380 15608 20408
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15580 20352 15669 20380
rect 15657 20349 15669 20352
rect 15703 20349 15715 20383
rect 15657 20343 15715 20349
rect 13280 20284 14044 20312
rect 14016 20256 14044 20284
rect 15194 20272 15200 20324
rect 15252 20312 15258 20324
rect 15764 20312 15792 20411
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 16816 20420 17049 20448
rect 16816 20408 16822 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18874 20448 18880 20460
rect 18739 20420 18880 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 18966 20408 18972 20460
rect 19024 20408 19030 20460
rect 19153 20451 19211 20457
rect 19153 20417 19165 20451
rect 19199 20448 19211 20451
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 19199 20420 19257 20448
rect 19199 20417 19211 20420
rect 19153 20411 19211 20417
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 20732 20448 20760 20544
rect 25038 20516 25044 20528
rect 24872 20488 25044 20516
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20732 20420 20821 20448
rect 19245 20411 19303 20417
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20448 22155 20451
rect 22143 20420 22876 20448
rect 22143 20417 22155 20420
rect 22097 20411 22155 20417
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17770 20380 17776 20392
rect 17359 20352 17776 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 15252 20284 15792 20312
rect 17144 20312 17172 20343
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 18782 20340 18788 20392
rect 18840 20340 18846 20392
rect 21082 20340 21088 20392
rect 21140 20340 21146 20392
rect 21450 20340 21456 20392
rect 21508 20380 21514 20392
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 21508 20352 21833 20380
rect 21508 20340 21514 20352
rect 21821 20349 21833 20352
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 17402 20312 17408 20324
rect 17144 20284 17408 20312
rect 15252 20272 15258 20284
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 18690 20272 18696 20324
rect 18748 20312 18754 20324
rect 18877 20315 18935 20321
rect 18877 20312 18889 20315
rect 18748 20284 18889 20312
rect 18748 20272 18754 20284
rect 18877 20281 18889 20284
rect 18923 20281 18935 20315
rect 18877 20275 18935 20281
rect 22848 20256 22876 20420
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23293 20451 23351 20457
rect 23293 20448 23305 20451
rect 23072 20420 23305 20448
rect 23072 20408 23078 20420
rect 23293 20417 23305 20420
rect 23339 20417 23351 20451
rect 23293 20411 23351 20417
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 24872 20457 24900 20488
rect 25038 20476 25044 20488
rect 25096 20516 25102 20528
rect 25222 20516 25228 20528
rect 25096 20488 25228 20516
rect 25096 20476 25102 20488
rect 25222 20476 25228 20488
rect 25280 20476 25286 20528
rect 26694 20476 26700 20528
rect 26752 20516 26758 20528
rect 28828 20516 28856 20544
rect 28920 20525 28948 20556
rect 26752 20488 28856 20516
rect 28905 20519 28963 20525
rect 26752 20476 26758 20488
rect 28905 20485 28917 20519
rect 28951 20485 28963 20519
rect 28905 20479 28963 20485
rect 28994 20476 29000 20528
rect 29052 20476 29058 20528
rect 29288 20516 29316 20556
rect 29641 20519 29699 20525
rect 29641 20516 29653 20519
rect 29288 20488 29653 20516
rect 29641 20485 29653 20488
rect 29687 20516 29699 20519
rect 29687 20488 30144 20516
rect 29687 20485 29699 20488
rect 29641 20479 29699 20485
rect 23569 20451 23627 20457
rect 23569 20448 23581 20451
rect 23440 20420 23581 20448
rect 23440 20408 23446 20420
rect 23569 20417 23581 20420
rect 23615 20417 23627 20451
rect 23569 20411 23627 20417
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 24857 20451 24915 20457
rect 24857 20417 24869 20451
rect 24903 20417 24915 20451
rect 28721 20451 28779 20457
rect 28721 20448 28733 20451
rect 24857 20411 24915 20417
rect 28184 20420 28733 20448
rect 22922 20340 22928 20392
rect 22980 20340 22986 20392
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 23860 20380 23888 20411
rect 23532 20352 23888 20380
rect 23532 20340 23538 20352
rect 23385 20315 23443 20321
rect 23385 20281 23397 20315
rect 23431 20312 23443 20315
rect 23842 20312 23848 20324
rect 23431 20284 23848 20312
rect 23431 20281 23443 20284
rect 23385 20275 23443 20281
rect 23842 20272 23848 20284
rect 23900 20272 23906 20324
rect 28184 20256 28212 20420
rect 28721 20417 28733 20420
rect 28767 20417 28779 20451
rect 28721 20411 28779 20417
rect 28813 20451 28871 20457
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 29012 20446 29040 20476
rect 30116 20460 30144 20488
rect 29089 20451 29147 20457
rect 29089 20446 29101 20451
rect 29012 20418 29101 20446
rect 28813 20411 28871 20417
rect 29089 20417 29101 20418
rect 29135 20417 29147 20451
rect 29454 20448 29460 20460
rect 29089 20411 29147 20417
rect 29181 20441 29239 20447
rect 28534 20340 28540 20392
rect 28592 20340 28598 20392
rect 12253 20247 12311 20253
rect 12253 20244 12265 20247
rect 11256 20216 12265 20244
rect 12253 20213 12265 20216
rect 12299 20213 12311 20247
rect 12253 20207 12311 20213
rect 12342 20204 12348 20256
rect 12400 20244 12406 20256
rect 12437 20247 12495 20253
rect 12437 20244 12449 20247
rect 12400 20216 12449 20244
rect 12400 20204 12406 20216
rect 12437 20213 12449 20216
rect 12483 20213 12495 20247
rect 12437 20207 12495 20213
rect 12710 20204 12716 20256
rect 12768 20204 12774 20256
rect 13630 20204 13636 20256
rect 13688 20204 13694 20256
rect 13998 20204 14004 20256
rect 14056 20204 14062 20256
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19484 20216 19625 20244
rect 19484 20204 19490 20216
rect 19613 20213 19625 20216
rect 19659 20213 19671 20247
rect 19613 20207 19671 20213
rect 22830 20204 22836 20256
rect 22888 20204 22894 20256
rect 24946 20204 24952 20256
rect 25004 20204 25010 20256
rect 28166 20204 28172 20256
rect 28224 20204 28230 20256
rect 28552 20244 28580 20340
rect 28736 20312 28764 20411
rect 28828 20380 28856 20411
rect 29181 20407 29193 20441
rect 29227 20438 29239 20441
rect 29288 20438 29460 20448
rect 29227 20420 29460 20438
rect 29227 20410 29316 20420
rect 29227 20407 29239 20410
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 29733 20451 29791 20457
rect 29733 20448 29745 20451
rect 29564 20420 29745 20448
rect 29181 20401 29239 20407
rect 28828 20352 29132 20380
rect 29104 20324 29132 20352
rect 28994 20312 29000 20324
rect 28736 20284 29000 20312
rect 28994 20272 29000 20284
rect 29052 20272 29058 20324
rect 29086 20272 29092 20324
rect 29144 20272 29150 20324
rect 28902 20244 28908 20256
rect 28552 20216 28908 20244
rect 28902 20204 28908 20216
rect 28960 20244 28966 20256
rect 29273 20247 29331 20253
rect 29273 20244 29285 20247
rect 28960 20216 29285 20244
rect 28960 20204 28966 20216
rect 29273 20213 29285 20216
rect 29319 20213 29331 20247
rect 29472 20244 29500 20408
rect 29564 20392 29592 20420
rect 29733 20417 29745 20420
rect 29779 20448 29791 20451
rect 29825 20451 29883 20457
rect 29825 20448 29837 20451
rect 29779 20420 29837 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 29825 20417 29837 20420
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 29546 20340 29552 20392
rect 29604 20340 29610 20392
rect 29917 20247 29975 20253
rect 29917 20244 29929 20247
rect 29472 20216 29929 20244
rect 29273 20207 29331 20213
rect 29917 20213 29929 20216
rect 29963 20213 29975 20247
rect 29917 20207 29975 20213
rect 30282 20204 30288 20256
rect 30340 20204 30346 20256
rect 1104 20154 30820 20176
rect 1104 20102 4664 20154
rect 4716 20102 4728 20154
rect 4780 20102 4792 20154
rect 4844 20102 4856 20154
rect 4908 20102 4920 20154
rect 4972 20102 12092 20154
rect 12144 20102 12156 20154
rect 12208 20102 12220 20154
rect 12272 20102 12284 20154
rect 12336 20102 12348 20154
rect 12400 20102 19520 20154
rect 19572 20102 19584 20154
rect 19636 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 26948 20154
rect 27000 20102 27012 20154
rect 27064 20102 27076 20154
rect 27128 20102 27140 20154
rect 27192 20102 27204 20154
rect 27256 20102 30820 20154
rect 1104 20080 30820 20102
rect 2774 20000 2780 20052
rect 2832 20040 2838 20052
rect 3053 20043 3111 20049
rect 3053 20040 3065 20043
rect 2832 20012 3065 20040
rect 2832 20000 2838 20012
rect 3053 20009 3065 20012
rect 3099 20009 3111 20043
rect 3053 20003 3111 20009
rect 3878 20000 3884 20052
rect 3936 20000 3942 20052
rect 4338 20000 4344 20052
rect 4396 20000 4402 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 8205 20043 8263 20049
rect 8205 20040 8217 20043
rect 7984 20012 8217 20040
rect 7984 20000 7990 20012
rect 8205 20009 8217 20012
rect 8251 20009 8263 20043
rect 8205 20003 8263 20009
rect 9140 20012 10824 20040
rect 4356 19904 4384 20000
rect 8941 19975 8999 19981
rect 8941 19972 8953 19975
rect 3252 19876 4384 19904
rect 4816 19944 8953 19972
rect 3252 19845 3280 19876
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 1688 19768 1716 19799
rect 3694 19796 3700 19848
rect 3752 19836 3758 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3752 19808 3985 19836
rect 3752 19796 3758 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4816 19768 4844 19944
rect 8941 19941 8953 19944
rect 8987 19941 8999 19975
rect 8941 19935 8999 19941
rect 4982 19864 4988 19916
rect 5040 19904 5046 19916
rect 5040 19876 5304 19904
rect 5040 19864 5046 19876
rect 5276 19845 5304 19876
rect 5350 19864 5356 19916
rect 5408 19864 5414 19916
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 7469 19907 7527 19913
rect 7469 19904 7481 19907
rect 7432 19876 7481 19904
rect 7432 19864 7438 19876
rect 7469 19873 7481 19876
rect 7515 19904 7527 19907
rect 9140 19904 9168 20012
rect 7515 19876 8156 19904
rect 7515 19873 7527 19876
rect 7469 19867 7527 19873
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 5261 19839 5319 19845
rect 4939 19808 5212 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 1688 19740 4844 19768
rect 4985 19771 5043 19777
rect 4985 19737 4997 19771
rect 5031 19737 5043 19771
rect 4985 19731 5043 19737
rect 5077 19771 5135 19777
rect 5077 19737 5089 19771
rect 5123 19737 5135 19771
rect 5184 19768 5212 19808
rect 5261 19805 5273 19839
rect 5307 19805 5319 19839
rect 5261 19799 5319 19805
rect 5368 19768 5396 19864
rect 5534 19836 5540 19848
rect 5184 19740 5396 19768
rect 5460 19808 5540 19836
rect 5077 19731 5135 19737
rect 934 19660 940 19712
rect 992 19700 998 19712
rect 1489 19703 1547 19709
rect 1489 19700 1501 19703
rect 992 19672 1501 19700
rect 992 19660 998 19672
rect 1489 19669 1501 19672
rect 1535 19669 1547 19703
rect 1489 19663 1547 19669
rect 4706 19660 4712 19712
rect 4764 19660 4770 19712
rect 4890 19660 4896 19712
rect 4948 19700 4954 19712
rect 5000 19700 5028 19731
rect 4948 19672 5028 19700
rect 5092 19700 5120 19731
rect 5460 19700 5488 19808
rect 5534 19796 5540 19808
rect 5592 19836 5598 19848
rect 7745 19839 7803 19845
rect 5592 19808 7696 19836
rect 5592 19796 5598 19808
rect 5092 19672 5488 19700
rect 4948 19660 4954 19672
rect 6822 19660 6828 19712
rect 6880 19660 6886 19712
rect 7466 19660 7472 19712
rect 7524 19700 7530 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 7524 19672 7573 19700
rect 7524 19660 7530 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 7668 19700 7696 19808
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8018 19836 8024 19848
rect 7791 19808 8024 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 8018 19796 8024 19808
rect 8076 19796 8082 19848
rect 8128 19845 8156 19876
rect 8220 19876 9168 19904
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 7834 19728 7840 19780
rect 7892 19728 7898 19780
rect 7929 19771 7987 19777
rect 7929 19737 7941 19771
rect 7975 19737 7987 19771
rect 8036 19768 8064 19796
rect 8220 19768 8248 19876
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19836 8447 19839
rect 9030 19836 9036 19848
rect 8435 19808 9036 19836
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9140 19845 9168 19876
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 9585 19907 9643 19913
rect 9585 19904 9597 19907
rect 9364 19876 9597 19904
rect 9364 19864 9370 19876
rect 9508 19845 9536 19876
rect 9585 19873 9597 19876
rect 9631 19873 9643 19907
rect 9585 19867 9643 19873
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 10318 19904 10324 19916
rect 9824 19876 10324 19904
rect 9824 19864 9830 19876
rect 10318 19864 10324 19876
rect 10376 19904 10382 19916
rect 10597 19907 10655 19913
rect 10597 19904 10609 19907
rect 10376 19876 10609 19904
rect 10376 19864 10382 19876
rect 10597 19873 10609 19876
rect 10643 19873 10655 19907
rect 10796 19904 10824 20012
rect 11146 20000 11152 20052
rect 11204 20000 11210 20052
rect 12526 20040 12532 20052
rect 12406 20012 12532 20040
rect 11054 19932 11060 19984
rect 11112 19932 11118 19984
rect 12406 19972 12434 20012
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 13081 20043 13139 20049
rect 13081 20009 13093 20043
rect 13127 20040 13139 20043
rect 13354 20040 13360 20052
rect 13127 20012 13360 20040
rect 13127 20009 13139 20012
rect 13081 20003 13139 20009
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 17221 20043 17279 20049
rect 17221 20009 17233 20043
rect 17267 20040 17279 20043
rect 17310 20040 17316 20052
rect 17267 20012 17316 20040
rect 17267 20009 17279 20012
rect 17221 20003 17279 20009
rect 13906 19972 13912 19984
rect 11164 19944 12434 19972
rect 12544 19944 13912 19972
rect 11164 19904 11192 19944
rect 10796 19876 11192 19904
rect 10597 19867 10655 19873
rect 11606 19864 11612 19916
rect 11664 19864 11670 19916
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19805 9183 19839
rect 9493 19839 9551 19845
rect 9125 19799 9183 19805
rect 9232 19808 9444 19836
rect 9232 19777 9260 19808
rect 8036 19740 8248 19768
rect 9217 19771 9275 19777
rect 7929 19731 7987 19737
rect 9217 19737 9229 19771
rect 9263 19737 9275 19771
rect 9217 19731 9275 19737
rect 9309 19771 9367 19777
rect 9309 19737 9321 19771
rect 9355 19737 9367 19771
rect 9416 19768 9444 19808
rect 9493 19805 9505 19839
rect 9539 19836 9551 19839
rect 9539 19808 9573 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 10226 19796 10232 19848
rect 10284 19796 10290 19848
rect 12544 19845 12572 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 17144 19972 17172 20003
rect 17310 20000 17316 20012
rect 17368 20040 17374 20052
rect 17862 20040 17868 20052
rect 17368 20012 17868 20040
rect 17368 20000 17374 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 19334 20000 19340 20052
rect 19392 20000 19398 20052
rect 20070 20000 20076 20052
rect 20128 20040 20134 20052
rect 20165 20043 20223 20049
rect 20165 20040 20177 20043
rect 20128 20012 20177 20040
rect 20128 20000 20134 20012
rect 20165 20009 20177 20012
rect 20211 20009 20223 20043
rect 20165 20003 20223 20009
rect 23385 20043 23443 20049
rect 23385 20009 23397 20043
rect 23431 20040 23443 20043
rect 24118 20040 24124 20052
rect 23431 20012 24124 20040
rect 23431 20009 23443 20012
rect 23385 20003 23443 20009
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 27614 20040 27620 20052
rect 24688 20012 27620 20040
rect 17678 19972 17684 19984
rect 17144 19944 17684 19972
rect 17678 19932 17684 19944
rect 17736 19932 17742 19984
rect 16393 19907 16451 19913
rect 12636 19876 12940 19904
rect 12636 19848 12664 19876
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19836 10747 19839
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 10735 19808 11529 19836
rect 10735 19805 10747 19808
rect 10689 19799 10747 19805
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19805 12587 19839
rect 12529 19799 12587 19805
rect 10134 19768 10140 19780
rect 9416 19740 10140 19768
rect 9309 19731 9367 19737
rect 7944 19700 7972 19731
rect 9324 19700 9352 19731
rect 10134 19728 10140 19740
rect 10192 19768 10198 19780
rect 10704 19768 10732 19799
rect 12618 19796 12624 19848
rect 12676 19796 12682 19848
rect 12710 19796 12716 19848
rect 12768 19796 12774 19848
rect 12912 19845 12940 19876
rect 16393 19873 16405 19907
rect 16439 19904 16451 19907
rect 17034 19904 17040 19916
rect 16439 19876 17040 19904
rect 16439 19873 16451 19876
rect 16393 19867 16451 19873
rect 17034 19864 17040 19876
rect 17092 19904 17098 19916
rect 17129 19907 17187 19913
rect 17129 19904 17141 19907
rect 17092 19876 17141 19904
rect 17092 19864 17098 19876
rect 17129 19873 17141 19876
rect 17175 19873 17187 19907
rect 19150 19904 19156 19916
rect 17129 19867 17187 19873
rect 17512 19876 19156 19904
rect 17512 19848 17540 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 20990 19864 20996 19916
rect 21048 19864 21054 19916
rect 21174 19864 21180 19916
rect 21232 19864 21238 19916
rect 22922 19864 22928 19916
rect 22980 19864 22986 19916
rect 24688 19904 24716 20012
rect 27614 20000 27620 20012
rect 27672 20000 27678 20052
rect 27985 20043 28043 20049
rect 27985 20009 27997 20043
rect 28031 20009 28043 20043
rect 27985 20003 28043 20009
rect 24765 19975 24823 19981
rect 24765 19941 24777 19975
rect 24811 19941 24823 19975
rect 25406 19972 25412 19984
rect 24765 19935 24823 19941
rect 25332 19944 25412 19972
rect 23216 19876 24716 19904
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 12728 19768 12756 19796
rect 10192 19740 10732 19768
rect 11256 19740 12756 19768
rect 12805 19771 12863 19777
rect 10192 19728 10198 19740
rect 11256 19700 11284 19740
rect 12805 19737 12817 19771
rect 12851 19737 12863 19771
rect 12805 19731 12863 19737
rect 7668 19672 11284 19700
rect 7561 19663 7619 19669
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12820 19700 12848 19731
rect 16040 19712 16068 19799
rect 16206 19796 16212 19848
rect 16264 19796 16270 19848
rect 17313 19839 17371 19845
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 17494 19836 17500 19848
rect 17359 19808 17500 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 18598 19796 18604 19848
rect 18656 19796 18662 19848
rect 18785 19839 18843 19845
rect 18785 19805 18797 19839
rect 18831 19836 18843 19839
rect 18831 19808 18920 19836
rect 18831 19805 18843 19808
rect 18785 19799 18843 19805
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19768 17003 19771
rect 17218 19768 17224 19780
rect 16991 19740 17224 19768
rect 16991 19737 17003 19740
rect 16945 19731 17003 19737
rect 17218 19728 17224 19740
rect 17276 19728 17282 19780
rect 18892 19712 18920 19808
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20070 19836 20076 19848
rect 19935 19808 20076 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19836 20499 19839
rect 20530 19836 20536 19848
rect 20487 19808 20536 19836
rect 20487 19805 20499 19808
rect 20441 19799 20499 19805
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 20714 19836 20720 19848
rect 20671 19808 20720 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 20864 19808 21036 19836
rect 20864 19796 20870 19808
rect 21008 19768 21036 19808
rect 22830 19796 22836 19848
rect 22888 19836 22894 19848
rect 23216 19836 23244 19876
rect 22888 19808 23244 19836
rect 23293 19839 23351 19845
rect 22888 19796 22894 19808
rect 23293 19805 23305 19839
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 21008 19740 22094 19768
rect 11664 19672 12848 19700
rect 11664 19660 11670 19672
rect 16022 19660 16028 19712
rect 16080 19660 16086 19712
rect 18690 19660 18696 19712
rect 18748 19660 18754 19712
rect 18874 19660 18880 19712
rect 18932 19660 18938 19712
rect 22066 19700 22094 19740
rect 23014 19728 23020 19780
rect 23072 19768 23078 19780
rect 23308 19768 23336 19799
rect 23382 19796 23388 19848
rect 23440 19836 23446 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23440 19808 23581 19836
rect 23440 19796 23446 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19836 24731 19839
rect 24780 19836 24808 19935
rect 25332 19913 25360 19944
rect 25406 19932 25412 19944
rect 25464 19932 25470 19984
rect 28000 19972 28028 20003
rect 28166 20000 28172 20052
rect 28224 20000 28230 20052
rect 28258 20000 28264 20052
rect 28316 20000 28322 20052
rect 28721 20043 28779 20049
rect 28721 20009 28733 20043
rect 28767 20040 28779 20043
rect 29454 20040 29460 20052
rect 28767 20012 29460 20040
rect 28767 20009 28779 20012
rect 28721 20003 28779 20009
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 30282 20000 30288 20052
rect 30340 20000 30346 20052
rect 28276 19972 28304 20000
rect 28537 19975 28595 19981
rect 28537 19972 28549 19975
rect 28000 19944 28549 19972
rect 28537 19941 28549 19944
rect 28583 19941 28595 19975
rect 28537 19935 28595 19941
rect 29086 19932 29092 19984
rect 29144 19932 29150 19984
rect 29181 19975 29239 19981
rect 29181 19941 29193 19975
rect 29227 19972 29239 19975
rect 30300 19972 30328 20000
rect 29227 19944 30328 19972
rect 29227 19941 29239 19944
rect 29181 19935 29239 19941
rect 25317 19907 25375 19913
rect 25317 19873 25329 19907
rect 25363 19873 25375 19907
rect 25593 19907 25651 19913
rect 25593 19904 25605 19907
rect 25317 19867 25375 19873
rect 25424 19876 25605 19904
rect 24719 19808 24808 19836
rect 25133 19839 25191 19845
rect 24719 19805 24731 19808
rect 24673 19799 24731 19805
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25424 19836 25452 19876
rect 25593 19873 25605 19876
rect 25639 19904 25651 19907
rect 25774 19904 25780 19916
rect 25639 19876 25780 19904
rect 25639 19873 25651 19876
rect 25593 19867 25651 19873
rect 25774 19864 25780 19876
rect 25832 19904 25838 19916
rect 27433 19907 27491 19913
rect 25832 19876 27016 19904
rect 25832 19864 25838 19876
rect 25179 19808 25452 19836
rect 26988 19836 27016 19876
rect 27433 19873 27445 19907
rect 27479 19904 27491 19907
rect 27982 19904 27988 19916
rect 27479 19876 27988 19904
rect 27479 19873 27491 19876
rect 27433 19867 27491 19873
rect 27982 19864 27988 19876
rect 28040 19904 28046 19916
rect 28040 19876 28672 19904
rect 28040 19864 28046 19876
rect 27709 19839 27767 19845
rect 27709 19836 27721 19839
rect 26988 19808 27721 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 27709 19805 27721 19808
rect 27755 19836 27767 19839
rect 28261 19839 28319 19845
rect 28261 19836 28273 19839
rect 27755 19808 28273 19836
rect 27755 19805 27767 19808
rect 27709 19799 27767 19805
rect 28261 19805 28273 19808
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 23860 19768 23888 19799
rect 28644 19780 28672 19876
rect 28902 19864 28908 19916
rect 28960 19864 28966 19916
rect 28997 19907 29055 19913
rect 28997 19873 29009 19907
rect 29043 19904 29055 19907
rect 29270 19904 29276 19916
rect 29043 19876 29276 19904
rect 29043 19873 29055 19876
rect 28997 19867 29055 19873
rect 29270 19864 29276 19876
rect 29328 19864 29334 19916
rect 29271 19817 29329 19823
rect 29271 19783 29283 19817
rect 29317 19783 29329 19817
rect 29271 19780 29329 19783
rect 23072 19740 23336 19768
rect 23492 19740 23888 19768
rect 23072 19728 23078 19740
rect 23492 19712 23520 19740
rect 24210 19728 24216 19780
rect 24268 19768 24274 19780
rect 25777 19771 25835 19777
rect 25777 19768 25789 19771
rect 24268 19740 25789 19768
rect 24268 19728 24274 19740
rect 25777 19737 25789 19740
rect 25823 19737 25835 19771
rect 25777 19731 25835 19737
rect 28626 19728 28632 19780
rect 28684 19728 28690 19780
rect 29270 19728 29276 19780
rect 29328 19728 29334 19780
rect 23474 19700 23480 19712
rect 22066 19672 23480 19700
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 24486 19660 24492 19712
rect 24544 19660 24550 19712
rect 25222 19660 25228 19712
rect 25280 19660 25286 19712
rect 29086 19660 29092 19712
rect 29144 19700 29150 19712
rect 29638 19700 29644 19712
rect 29144 19672 29644 19700
rect 29144 19660 29150 19672
rect 29638 19660 29644 19672
rect 29696 19660 29702 19712
rect 1104 19610 30820 19632
rect 1104 19558 5324 19610
rect 5376 19558 5388 19610
rect 5440 19558 5452 19610
rect 5504 19558 5516 19610
rect 5568 19558 5580 19610
rect 5632 19558 12752 19610
rect 12804 19558 12816 19610
rect 12868 19558 12880 19610
rect 12932 19558 12944 19610
rect 12996 19558 13008 19610
rect 13060 19558 20180 19610
rect 20232 19558 20244 19610
rect 20296 19558 20308 19610
rect 20360 19558 20372 19610
rect 20424 19558 20436 19610
rect 20488 19558 27608 19610
rect 27660 19558 27672 19610
rect 27724 19558 27736 19610
rect 27788 19558 27800 19610
rect 27852 19558 27864 19610
rect 27916 19558 30820 19610
rect 1104 19536 30820 19558
rect 4706 19496 4712 19508
rect 2746 19468 4712 19496
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 2746 19360 2774 19468
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 6365 19499 6423 19505
rect 6365 19465 6377 19499
rect 6411 19465 6423 19499
rect 6365 19459 6423 19465
rect 1719 19332 2774 19360
rect 5721 19363 5779 19369
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 5721 19329 5733 19363
rect 5767 19360 5779 19363
rect 6380 19360 6408 19459
rect 6454 19456 6460 19508
rect 6512 19456 6518 19508
rect 6733 19499 6791 19505
rect 6733 19465 6745 19499
rect 6779 19496 6791 19499
rect 6822 19496 6828 19508
rect 6779 19468 6828 19496
rect 6779 19465 6791 19468
rect 6733 19459 6791 19465
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 8478 19496 8484 19508
rect 7576 19468 8484 19496
rect 5767 19332 6408 19360
rect 6472 19360 6500 19456
rect 7576 19372 7604 19468
rect 8478 19456 8484 19468
rect 8536 19496 8542 19508
rect 9490 19496 9496 19508
rect 8536 19468 9496 19496
rect 8536 19456 8542 19468
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 9769 19499 9827 19505
rect 9769 19465 9781 19499
rect 9815 19496 9827 19499
rect 10226 19496 10232 19508
rect 9815 19468 10232 19496
rect 9815 19465 9827 19468
rect 9769 19459 9827 19465
rect 10226 19456 10232 19468
rect 10284 19456 10290 19508
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 16022 19496 16028 19508
rect 10468 19468 16028 19496
rect 10468 19456 10474 19468
rect 7837 19431 7895 19437
rect 7837 19397 7849 19431
rect 7883 19428 7895 19431
rect 7926 19428 7932 19440
rect 7883 19400 7932 19428
rect 7883 19397 7895 19400
rect 7837 19391 7895 19397
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 8570 19388 8576 19440
rect 8628 19388 8634 19440
rect 9122 19388 9128 19440
rect 9180 19388 9186 19440
rect 12452 19400 14228 19428
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6472 19332 6837 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 7558 19320 7564 19372
rect 7616 19320 7622 19372
rect 9140 19360 9168 19388
rect 12452 19369 12480 19400
rect 12437 19363 12495 19369
rect 9140 19332 9444 19360
rect 4982 19252 4988 19304
rect 5040 19252 5046 19304
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 4522 19184 4528 19236
rect 4580 19224 4586 19236
rect 5074 19224 5080 19236
rect 4580 19196 5080 19224
rect 4580 19184 4586 19196
rect 5074 19184 5080 19196
rect 5132 19224 5138 19236
rect 7024 19224 7052 19255
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 9416 19233 9444 19332
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12526 19320 12532 19372
rect 12584 19320 12590 19372
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19360 12679 19363
rect 12667 19332 13860 19360
rect 12667 19329 12679 19332
rect 12621 19323 12679 19329
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 9824 19264 9873 19292
rect 9824 19252 9830 19264
rect 9861 19261 9873 19264
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 5132 19196 7052 19224
rect 5132 19184 5138 19196
rect 1486 19116 1492 19168
rect 1544 19116 1550 19168
rect 4430 19116 4436 19168
rect 4488 19116 4494 19168
rect 5534 19116 5540 19168
rect 5592 19116 5598 19168
rect 7024 19156 7052 19196
rect 9401 19227 9459 19233
rect 9401 19193 9413 19227
rect 9447 19193 9459 19227
rect 9968 19224 9996 19255
rect 12618 19224 12624 19236
rect 9401 19187 9459 19193
rect 9646 19196 12624 19224
rect 9646 19156 9674 19196
rect 12618 19184 12624 19196
rect 12676 19224 12682 19236
rect 13630 19224 13636 19236
rect 12676 19196 13636 19224
rect 12676 19184 12682 19196
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 13832 19224 13860 19332
rect 13906 19320 13912 19372
rect 13964 19320 13970 19372
rect 13924 19292 13952 19320
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 13924 19264 14013 19292
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14001 19255 14059 19261
rect 14090 19224 14096 19236
rect 13832 19196 14096 19224
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 14200 19224 14228 19400
rect 14292 19369 14320 19468
rect 16022 19456 16028 19468
rect 16080 19496 16086 19508
rect 16758 19496 16764 19508
rect 16080 19468 16764 19496
rect 16080 19456 16086 19468
rect 14458 19388 14464 19440
rect 14516 19388 14522 19440
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 16206 19320 16212 19372
rect 16264 19320 16270 19372
rect 16408 19369 16436 19468
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 17402 19456 17408 19508
rect 17460 19456 17466 19508
rect 18414 19496 18420 19508
rect 17972 19468 18420 19496
rect 17037 19431 17095 19437
rect 17037 19397 17049 19431
rect 17083 19428 17095 19431
rect 17972 19428 18000 19468
rect 18414 19456 18420 19468
rect 18472 19456 18478 19508
rect 18690 19456 18696 19508
rect 18748 19456 18754 19508
rect 18782 19456 18788 19508
rect 18840 19456 18846 19508
rect 19426 19456 19432 19508
rect 19484 19456 19490 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 21910 19496 21916 19508
rect 20128 19468 21916 19496
rect 20128 19456 20134 19468
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 24486 19496 24492 19508
rect 24320 19468 24492 19496
rect 18708 19428 18736 19456
rect 17083 19400 18000 19428
rect 18064 19400 18736 19428
rect 18800 19428 18828 19456
rect 18969 19431 19027 19437
rect 18969 19428 18981 19431
rect 18800 19400 18981 19428
rect 17083 19397 17095 19400
rect 17037 19391 17095 19397
rect 16942 19369 16948 19372
rect 16393 19363 16451 19369
rect 16393 19329 16405 19363
rect 16439 19329 16451 19363
rect 16393 19323 16451 19329
rect 16919 19363 16948 19369
rect 16919 19329 16931 19363
rect 16919 19323 16948 19329
rect 16942 19320 16948 19323
rect 17000 19320 17006 19372
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17678 19360 17684 19372
rect 17267 19332 17684 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 15102 19252 15108 19304
rect 15160 19252 15166 19304
rect 16758 19252 16764 19304
rect 16816 19252 16822 19304
rect 17144 19292 17172 19323
rect 17678 19320 17684 19332
rect 17736 19320 17742 19372
rect 17862 19320 17868 19372
rect 17920 19320 17926 19372
rect 18064 19369 18092 19400
rect 18969 19397 18981 19400
rect 19015 19397 19027 19431
rect 18969 19391 19027 19397
rect 20530 19388 20536 19440
rect 20588 19428 20594 19440
rect 20588 19400 23060 19428
rect 20588 19388 20594 19400
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 18233 19363 18291 19369
rect 18233 19329 18245 19363
rect 18279 19334 18291 19363
rect 18351 19363 18409 19369
rect 18279 19329 18313 19334
rect 18233 19323 18313 19329
rect 18351 19329 18363 19363
rect 18397 19360 18409 19363
rect 18598 19360 18604 19372
rect 18397 19332 18604 19360
rect 18397 19329 18409 19332
rect 18351 19323 18409 19329
rect 18248 19306 18313 19323
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19360 18843 19363
rect 18874 19360 18880 19372
rect 18831 19332 18880 19360
rect 18831 19329 18843 19332
rect 18785 19323 18843 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19208 19332 19257 19360
rect 19208 19320 19214 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 19334 19320 19340 19372
rect 19392 19320 19398 19372
rect 20073 19363 20131 19369
rect 20073 19360 20085 19363
rect 19444 19332 20085 19360
rect 17586 19292 17592 19304
rect 17144 19264 17592 19292
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17770 19252 17776 19304
rect 17828 19292 17834 19304
rect 18248 19292 18276 19306
rect 17828 19264 18276 19292
rect 18509 19295 18567 19301
rect 17828 19252 17834 19264
rect 14826 19224 14832 19236
rect 14200 19196 14832 19224
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 16209 19227 16267 19233
rect 16209 19193 16221 19227
rect 16255 19224 16267 19227
rect 17218 19224 17224 19236
rect 16255 19196 17224 19224
rect 16255 19193 16267 19196
rect 16209 19187 16267 19193
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 7024 19128 9674 19156
rect 13354 19116 13360 19168
rect 13412 19116 13418 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 17880 19156 17908 19264
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 19352 19292 19380 19320
rect 18555 19264 19380 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 18601 19227 18659 19233
rect 18601 19193 18613 19227
rect 18647 19193 18659 19227
rect 19444 19224 19472 19332
rect 20073 19329 20085 19332
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19360 20407 19363
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20395 19332 20637 19360
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 20625 19329 20637 19332
rect 20671 19360 20683 19363
rect 20806 19360 20812 19372
rect 20671 19332 20812 19360
rect 20671 19329 20683 19332
rect 20625 19323 20683 19329
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 21100 19369 21128 19400
rect 23032 19372 23060 19400
rect 23382 19388 23388 19440
rect 23440 19388 23446 19440
rect 24210 19428 24216 19440
rect 23860 19400 24216 19428
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 20993 19323 21051 19329
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19329 21143 19363
rect 21910 19360 21916 19372
rect 21085 19323 21143 19329
rect 21652 19332 21916 19360
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21008 19292 21036 19323
rect 20772 19264 21036 19292
rect 20772 19252 20778 19264
rect 18601 19187 18659 19193
rect 19306 19196 19472 19224
rect 13872 19128 17908 19156
rect 13872 19116 13878 19128
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18616 19156 18644 19187
rect 18196 19128 18644 19156
rect 18196 19116 18202 19128
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19306 19156 19334 19196
rect 20916 19168 20944 19264
rect 21174 19252 21180 19304
rect 21232 19252 21238 19304
rect 21652 19301 21680 19332
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22553 19363 22611 19369
rect 22553 19329 22565 19363
rect 22599 19329 22611 19363
rect 22553 19323 22611 19329
rect 21637 19295 21695 19301
rect 21637 19261 21649 19295
rect 21683 19261 21695 19295
rect 21928 19292 21956 19320
rect 22572 19292 22600 19323
rect 23014 19320 23020 19372
rect 23072 19320 23078 19372
rect 23293 19363 23351 19369
rect 23293 19329 23305 19363
rect 23339 19360 23351 19363
rect 23400 19360 23428 19388
rect 23339 19332 23428 19360
rect 23339 19329 23351 19332
rect 23293 19323 23351 19329
rect 23474 19320 23480 19372
rect 23532 19320 23538 19372
rect 22922 19292 22928 19304
rect 21928 19264 22928 19292
rect 21637 19255 21695 19261
rect 22922 19252 22928 19264
rect 22980 19252 22986 19304
rect 23385 19295 23443 19301
rect 23385 19261 23397 19295
rect 23431 19292 23443 19295
rect 23860 19292 23888 19400
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 24320 19437 24348 19468
rect 24486 19456 24492 19468
rect 24544 19456 24550 19508
rect 25222 19456 25228 19508
rect 25280 19496 25286 19508
rect 26145 19499 26203 19505
rect 26145 19496 26157 19499
rect 25280 19468 26157 19496
rect 25280 19456 25286 19468
rect 26145 19465 26157 19468
rect 26191 19465 26203 19499
rect 26786 19496 26792 19508
rect 26145 19459 26203 19465
rect 26436 19468 26792 19496
rect 24305 19431 24363 19437
rect 24305 19397 24317 19431
rect 24351 19397 24363 19431
rect 24305 19391 24363 19397
rect 24946 19388 24952 19440
rect 25004 19388 25010 19440
rect 25774 19388 25780 19440
rect 25832 19388 25838 19440
rect 23934 19320 23940 19372
rect 23992 19360 23998 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23992 19332 24041 19360
rect 23992 19320 23998 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 25792 19301 25820 19388
rect 26436 19372 26464 19468
rect 26786 19456 26792 19468
rect 26844 19456 26850 19508
rect 29457 19499 29515 19505
rect 29457 19496 29469 19499
rect 28092 19468 29469 19496
rect 26510 19388 26516 19440
rect 26568 19388 26574 19440
rect 26651 19431 26709 19437
rect 26651 19397 26663 19431
rect 26697 19428 26709 19431
rect 28092 19428 28120 19468
rect 29457 19465 29469 19468
rect 29503 19465 29515 19499
rect 29457 19459 29515 19465
rect 30282 19456 30288 19508
rect 30340 19456 30346 19508
rect 30300 19428 30328 19456
rect 26697 19400 28120 19428
rect 29196 19400 30328 19428
rect 26697 19397 26709 19400
rect 26651 19391 26709 19397
rect 26326 19320 26332 19372
rect 26384 19320 26390 19372
rect 26418 19320 26424 19372
rect 26476 19320 26482 19372
rect 27249 19363 27307 19369
rect 27249 19329 27261 19363
rect 27295 19360 27307 19363
rect 27982 19360 27988 19372
rect 27295 19332 27988 19360
rect 27295 19329 27307 19332
rect 27249 19323 27307 19329
rect 27982 19320 27988 19332
rect 28040 19320 28046 19372
rect 29196 19369 29224 19400
rect 29089 19363 29147 19369
rect 29089 19329 29101 19363
rect 29135 19329 29147 19363
rect 29089 19323 29147 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19329 29239 19363
rect 29181 19323 29239 19329
rect 23431 19264 23888 19292
rect 25777 19295 25835 19301
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 25777 19261 25789 19295
rect 25823 19261 25835 19295
rect 25777 19255 25835 19261
rect 26234 19252 26240 19304
rect 26292 19292 26298 19304
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 26292 19264 26801 19292
rect 26292 19252 26298 19264
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 26878 19252 26884 19304
rect 26936 19292 26942 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26936 19264 26985 19292
rect 26936 19252 26942 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 26973 19255 27031 19261
rect 29104 19224 29132 19323
rect 29362 19320 29368 19372
rect 29420 19320 29426 19372
rect 29840 19369 29868 19400
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19329 29883 19363
rect 29825 19323 29883 19329
rect 30098 19320 30104 19372
rect 30156 19320 30162 19372
rect 30285 19363 30343 19369
rect 30285 19329 30297 19363
rect 30331 19329 30343 19363
rect 30285 19323 30343 19329
rect 29917 19295 29975 19301
rect 29917 19261 29929 19295
rect 29963 19292 29975 19295
rect 30193 19295 30251 19301
rect 30193 19292 30205 19295
rect 29963 19264 30205 19292
rect 29963 19261 29975 19264
rect 29917 19255 29975 19261
rect 30193 19261 30205 19264
rect 30239 19261 30251 19295
rect 30193 19255 30251 19261
rect 28828 19196 29040 19224
rect 29104 19196 29224 19224
rect 28828 19168 28856 19196
rect 18932 19128 19334 19156
rect 18932 19116 18938 19128
rect 20898 19116 20904 19168
rect 20956 19116 20962 19168
rect 23290 19116 23296 19168
rect 23348 19156 23354 19168
rect 27338 19156 27344 19168
rect 23348 19128 27344 19156
rect 23348 19116 23354 19128
rect 27338 19116 27344 19128
rect 27396 19156 27402 19168
rect 27890 19156 27896 19168
rect 27396 19128 27896 19156
rect 27396 19116 27402 19128
rect 27890 19116 27896 19128
rect 27948 19116 27954 19168
rect 27985 19159 28043 19165
rect 27985 19125 27997 19159
rect 28031 19156 28043 19159
rect 28258 19156 28264 19168
rect 28031 19128 28264 19156
rect 28031 19125 28043 19128
rect 27985 19119 28043 19125
rect 28258 19116 28264 19128
rect 28316 19116 28322 19168
rect 28810 19116 28816 19168
rect 28868 19116 28874 19168
rect 28902 19116 28908 19168
rect 28960 19116 28966 19168
rect 29012 19156 29040 19196
rect 29196 19168 29224 19196
rect 29270 19184 29276 19236
rect 29328 19224 29334 19236
rect 30300 19224 30328 19323
rect 29328 19196 30328 19224
rect 29328 19184 29334 19196
rect 29089 19159 29147 19165
rect 29089 19156 29101 19159
rect 29012 19128 29101 19156
rect 29089 19125 29101 19128
rect 29135 19125 29147 19159
rect 29089 19119 29147 19125
rect 29178 19116 29184 19168
rect 29236 19116 29242 19168
rect 1104 19066 30820 19088
rect 1104 19014 4664 19066
rect 4716 19014 4728 19066
rect 4780 19014 4792 19066
rect 4844 19014 4856 19066
rect 4908 19014 4920 19066
rect 4972 19014 12092 19066
rect 12144 19014 12156 19066
rect 12208 19014 12220 19066
rect 12272 19014 12284 19066
rect 12336 19014 12348 19066
rect 12400 19014 19520 19066
rect 19572 19014 19584 19066
rect 19636 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 26948 19066
rect 27000 19014 27012 19066
rect 27064 19014 27076 19066
rect 27128 19014 27140 19066
rect 27192 19014 27204 19066
rect 27256 19014 30820 19066
rect 1104 18992 30820 19014
rect 6825 18955 6883 18961
rect 1688 18924 6408 18952
rect 1688 18757 1716 18924
rect 6380 18884 6408 18924
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 7374 18952 7380 18964
rect 6871 18924 7380 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 7374 18912 7380 18924
rect 7432 18912 7438 18964
rect 7466 18912 7472 18964
rect 7524 18912 7530 18964
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 8665 18955 8723 18961
rect 8665 18952 8677 18955
rect 8628 18924 8677 18952
rect 8628 18912 8634 18924
rect 8665 18921 8677 18924
rect 8711 18921 8723 18955
rect 8665 18915 8723 18921
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 13814 18952 13820 18964
rect 9916 18924 13820 18952
rect 9916 18912 9922 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 13906 18912 13912 18964
rect 13964 18912 13970 18964
rect 16301 18955 16359 18961
rect 16301 18921 16313 18955
rect 16347 18952 16359 18955
rect 16758 18952 16764 18964
rect 16347 18924 16764 18952
rect 16347 18921 16359 18924
rect 16301 18915 16359 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 17310 18912 17316 18964
rect 17368 18912 17374 18964
rect 17586 18912 17592 18964
rect 17644 18912 17650 18964
rect 18049 18955 18107 18961
rect 18049 18921 18061 18955
rect 18095 18952 18107 18955
rect 18322 18952 18328 18964
rect 18095 18924 18328 18952
rect 18095 18921 18107 18924
rect 18049 18915 18107 18921
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 19058 18912 19064 18964
rect 19116 18912 19122 18964
rect 19150 18912 19156 18964
rect 19208 18952 19214 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 19208 18924 19257 18952
rect 19208 18912 19214 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 19245 18915 19303 18921
rect 26326 18912 26332 18964
rect 26384 18952 26390 18964
rect 27525 18955 27583 18961
rect 27525 18952 27537 18955
rect 26384 18924 27537 18952
rect 26384 18912 26390 18924
rect 27525 18921 27537 18924
rect 27571 18921 27583 18955
rect 28074 18952 28080 18964
rect 27525 18915 27583 18921
rect 27632 18924 28080 18952
rect 7484 18884 7512 18912
rect 6380 18856 7512 18884
rect 12069 18887 12127 18893
rect 12069 18853 12081 18887
rect 12115 18884 12127 18887
rect 15657 18887 15715 18893
rect 12115 18856 12296 18884
rect 12115 18853 12127 18856
rect 12069 18847 12127 18853
rect 4522 18776 4528 18828
rect 4580 18776 4586 18828
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18816 5135 18819
rect 7558 18816 7564 18828
rect 5123 18788 7564 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 3329 18751 3387 18757
rect 3329 18717 3341 18751
rect 3375 18717 3387 18751
rect 3329 18711 3387 18717
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 3694 18748 3700 18760
rect 3651 18720 3700 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 3344 18680 3372 18711
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 5092 18748 5120 18779
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 9548 18788 12173 18816
rect 9548 18776 9554 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12268 18816 12296 18856
rect 15657 18853 15669 18887
rect 15703 18884 15715 18887
rect 18138 18884 18144 18896
rect 15703 18856 15976 18884
rect 15703 18853 15715 18856
rect 15657 18847 15715 18853
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 12268 18788 12449 18816
rect 12161 18779 12219 18785
rect 12437 18785 12449 18788
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 3844 18720 5120 18748
rect 3844 18708 3850 18720
rect 7650 18708 7656 18760
rect 7708 18748 7714 18760
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 7708 18720 8585 18748
rect 7708 18708 7714 18720
rect 8573 18717 8585 18720
rect 8619 18748 8631 18751
rect 8619 18720 11744 18748
rect 8619 18717 8631 18720
rect 8573 18711 8631 18717
rect 4249 18683 4307 18689
rect 3344 18652 3924 18680
rect 934 18572 940 18624
rect 992 18612 998 18624
rect 1489 18615 1547 18621
rect 1489 18612 1501 18615
rect 992 18584 1501 18612
rect 992 18572 998 18584
rect 1489 18581 1501 18584
rect 1535 18581 1547 18615
rect 1489 18575 1547 18581
rect 3142 18572 3148 18624
rect 3200 18572 3206 18624
rect 3510 18572 3516 18624
rect 3568 18572 3574 18624
rect 3896 18621 3924 18652
rect 4249 18649 4261 18683
rect 4295 18680 4307 18683
rect 4430 18680 4436 18692
rect 4295 18652 4436 18680
rect 4295 18649 4307 18652
rect 4249 18643 4307 18649
rect 4430 18640 4436 18652
rect 4488 18640 4494 18692
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18649 5411 18683
rect 5353 18643 5411 18649
rect 3881 18615 3939 18621
rect 3881 18581 3893 18615
rect 3927 18581 3939 18615
rect 3881 18575 3939 18581
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 4890 18612 4896 18624
rect 4396 18584 4896 18612
rect 4396 18572 4402 18584
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 5368 18612 5396 18643
rect 6086 18640 6092 18692
rect 6144 18640 6150 18692
rect 11716 18624 11744 18720
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 14645 18751 14703 18757
rect 14332 18720 14596 18748
rect 14332 18708 14338 18720
rect 14185 18683 14243 18689
rect 14185 18680 14197 18683
rect 13662 18652 14197 18680
rect 14185 18649 14197 18652
rect 14231 18649 14243 18683
rect 14185 18643 14243 18649
rect 5534 18612 5540 18624
rect 5368 18584 5540 18612
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 14568 18612 14596 18720
rect 14645 18717 14657 18751
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14921 18751 14979 18757
rect 14921 18717 14933 18751
rect 14967 18748 14979 18751
rect 15102 18748 15108 18760
rect 14967 18720 15108 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 14660 18680 14688 18711
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15378 18708 15384 18760
rect 15436 18708 15442 18760
rect 15948 18757 15976 18856
rect 16040 18856 18144 18884
rect 16040 18825 16068 18856
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 18966 18844 18972 18896
rect 19024 18844 19030 18896
rect 19337 18887 19395 18893
rect 19337 18853 19349 18887
rect 19383 18853 19395 18887
rect 19337 18847 19395 18853
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 17218 18776 17224 18828
rect 17276 18776 17282 18828
rect 18601 18819 18659 18825
rect 17328 18788 18092 18816
rect 17328 18760 17356 18788
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16206 18748 16212 18760
rect 15979 18720 16212 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 17092 18720 17141 18748
rect 17092 18708 17098 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17494 18748 17500 18760
rect 17451 18720 17500 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 18064 18757 18092 18788
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 19242 18816 19248 18828
rect 18647 18788 19248 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 19242 18776 19248 18788
rect 19300 18816 19306 18828
rect 19352 18816 19380 18847
rect 23842 18844 23848 18896
rect 23900 18884 23906 18896
rect 27632 18884 27660 18924
rect 28074 18912 28080 18924
rect 28132 18912 28138 18964
rect 29270 18884 29276 18896
rect 23900 18856 27660 18884
rect 27908 18856 29276 18884
rect 23900 18844 23906 18856
rect 19300 18788 19380 18816
rect 22557 18819 22615 18825
rect 19300 18776 19306 18788
rect 22557 18785 22569 18819
rect 22603 18816 22615 18819
rect 22922 18816 22928 18828
rect 22603 18788 22928 18816
rect 22603 18785 22615 18788
rect 22557 18779 22615 18785
rect 22922 18776 22928 18788
rect 22980 18776 22986 18828
rect 23385 18819 23443 18825
rect 23385 18785 23397 18819
rect 23431 18816 23443 18819
rect 26510 18816 26516 18828
rect 23431 18788 26516 18816
rect 23431 18785 23443 18788
rect 23385 18779 23443 18785
rect 26510 18776 26516 18788
rect 26568 18776 26574 18828
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17644 18720 17877 18748
rect 17644 18708 17650 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 15396 18680 15424 18708
rect 14660 18652 15424 18680
rect 16850 18612 16856 18624
rect 14568 18584 16856 18612
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 17880 18612 17908 18711
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19024 18720 19717 18748
rect 19024 18708 19030 18720
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19886 18708 19892 18760
rect 19944 18748 19950 18760
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19944 18720 20177 18748
rect 19944 18708 19950 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 23014 18708 23020 18760
rect 23072 18708 23078 18760
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 20441 18683 20499 18689
rect 20441 18649 20453 18683
rect 20487 18680 20499 18683
rect 20898 18680 20904 18692
rect 20487 18652 20904 18680
rect 20487 18649 20499 18652
rect 20441 18643 20499 18649
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 23216 18680 23244 18711
rect 23474 18708 23480 18760
rect 23532 18708 23538 18760
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 27430 18708 27436 18760
rect 27488 18708 27494 18760
rect 27617 18751 27675 18757
rect 27617 18717 27629 18751
rect 27663 18717 27675 18751
rect 27908 18748 27936 18856
rect 29270 18844 29276 18856
rect 29328 18844 29334 18896
rect 27985 18819 28043 18825
rect 27985 18785 27997 18819
rect 28031 18816 28043 18819
rect 28629 18819 28687 18825
rect 28629 18816 28641 18819
rect 28031 18788 28641 18816
rect 28031 18785 28043 18788
rect 27985 18779 28043 18785
rect 28629 18785 28641 18788
rect 28675 18785 28687 18819
rect 28629 18779 28687 18785
rect 28077 18751 28135 18757
rect 28077 18748 28089 18751
rect 27908 18720 28089 18748
rect 27617 18711 27675 18717
rect 28077 18717 28089 18720
rect 28123 18717 28135 18751
rect 28077 18711 28135 18717
rect 23382 18680 23388 18692
rect 23216 18652 23388 18680
rect 23382 18640 23388 18652
rect 23440 18640 23446 18692
rect 27632 18680 27660 18711
rect 28166 18708 28172 18760
rect 28224 18708 28230 18760
rect 28261 18751 28319 18757
rect 28261 18717 28273 18751
rect 28307 18748 28319 18751
rect 28442 18748 28448 18760
rect 28307 18720 28448 18748
rect 28307 18717 28319 18720
rect 28261 18711 28319 18717
rect 28442 18708 28448 18720
rect 28500 18708 28506 18760
rect 28537 18751 28595 18757
rect 28537 18717 28549 18751
rect 28583 18717 28595 18751
rect 28537 18711 28595 18717
rect 28721 18751 28779 18757
rect 28721 18717 28733 18751
rect 28767 18748 28779 18751
rect 28767 18720 29132 18748
rect 28767 18717 28779 18720
rect 28721 18711 28779 18717
rect 28552 18680 28580 18711
rect 28810 18680 28816 18692
rect 23492 18652 26004 18680
rect 27632 18652 28304 18680
rect 23492 18612 23520 18652
rect 25976 18624 26004 18652
rect 28276 18624 28304 18652
rect 28368 18652 28816 18680
rect 28368 18624 28396 18652
rect 28810 18640 28816 18652
rect 28868 18680 28874 18692
rect 29104 18689 29132 18720
rect 28905 18683 28963 18689
rect 28905 18680 28917 18683
rect 28868 18652 28917 18680
rect 28868 18640 28874 18652
rect 28905 18649 28917 18652
rect 28951 18649 28963 18683
rect 28905 18643 28963 18649
rect 29089 18683 29147 18689
rect 29089 18649 29101 18683
rect 29135 18680 29147 18683
rect 29178 18680 29184 18692
rect 29135 18652 29184 18680
rect 29135 18649 29147 18652
rect 29089 18643 29147 18649
rect 29178 18640 29184 18652
rect 29236 18640 29242 18692
rect 17880 18584 23520 18612
rect 24394 18572 24400 18624
rect 24452 18572 24458 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26234 18572 26240 18624
rect 26292 18612 26298 18624
rect 27801 18615 27859 18621
rect 27801 18612 27813 18615
rect 26292 18584 27813 18612
rect 26292 18572 26298 18584
rect 27801 18581 27813 18584
rect 27847 18581 27859 18615
rect 27801 18575 27859 18581
rect 28258 18572 28264 18624
rect 28316 18572 28322 18624
rect 28350 18572 28356 18624
rect 28408 18572 28414 18624
rect 1104 18522 30820 18544
rect 1104 18470 5324 18522
rect 5376 18470 5388 18522
rect 5440 18470 5452 18522
rect 5504 18470 5516 18522
rect 5568 18470 5580 18522
rect 5632 18470 12752 18522
rect 12804 18470 12816 18522
rect 12868 18470 12880 18522
rect 12932 18470 12944 18522
rect 12996 18470 13008 18522
rect 13060 18470 20180 18522
rect 20232 18470 20244 18522
rect 20296 18470 20308 18522
rect 20360 18470 20372 18522
rect 20424 18470 20436 18522
rect 20488 18470 27608 18522
rect 27660 18470 27672 18522
rect 27724 18470 27736 18522
rect 27788 18470 27800 18522
rect 27852 18470 27864 18522
rect 27916 18470 30820 18522
rect 1104 18448 30820 18470
rect 3142 18368 3148 18420
rect 3200 18368 3206 18420
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 4433 18411 4491 18417
rect 3752 18380 4292 18408
rect 3752 18368 3758 18380
rect 2961 18343 3019 18349
rect 2961 18309 2973 18343
rect 3007 18340 3019 18343
rect 3160 18340 3188 18368
rect 3007 18312 3188 18340
rect 3007 18309 3019 18312
rect 2961 18303 3019 18309
rect 3510 18300 3516 18352
rect 3568 18300 3574 18352
rect 4264 18340 4292 18380
rect 4433 18377 4445 18411
rect 4479 18408 4491 18411
rect 4982 18408 4988 18420
rect 4479 18380 4988 18408
rect 4479 18377 4491 18380
rect 4433 18371 4491 18377
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 6086 18368 6092 18420
rect 6144 18368 6150 18420
rect 7650 18368 7656 18420
rect 7708 18368 7714 18420
rect 8956 18380 10364 18408
rect 7668 18340 7696 18368
rect 4264 18312 7696 18340
rect 2498 18232 2504 18284
rect 2556 18272 2562 18284
rect 6012 18281 6040 18312
rect 8956 18284 8984 18380
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 9600 18312 10241 18340
rect 2685 18275 2743 18281
rect 2685 18272 2697 18275
rect 2556 18244 2697 18272
rect 2556 18232 2562 18244
rect 2685 18241 2697 18244
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7190 18272 7196 18284
rect 7055 18244 7196 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 2700 18204 2728 18235
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 9600 18281 9628 18312
rect 10229 18309 10241 18312
rect 10275 18309 10287 18343
rect 10229 18303 10287 18309
rect 10336 18340 10364 18380
rect 11422 18368 11428 18420
rect 11480 18368 11486 18420
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 12345 18411 12403 18417
rect 12345 18408 12357 18411
rect 11940 18380 12357 18408
rect 11940 18368 11946 18380
rect 12345 18377 12357 18380
rect 12391 18377 12403 18411
rect 12345 18371 12403 18377
rect 12713 18411 12771 18417
rect 12713 18377 12725 18411
rect 12759 18408 12771 18411
rect 13354 18408 13360 18420
rect 12759 18380 13360 18408
rect 12759 18377 12771 18380
rect 12713 18371 12771 18377
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 14274 18368 14280 18420
rect 14332 18368 14338 18420
rect 18874 18408 18880 18420
rect 14476 18380 18880 18408
rect 11440 18340 11468 18368
rect 10336 18312 12020 18340
rect 10336 18281 10364 18312
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18241 9183 18275
rect 9125 18235 9183 18241
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18241 9827 18275
rect 9769 18235 9827 18241
rect 9887 18276 9945 18281
rect 9887 18275 10012 18276
rect 9887 18241 9899 18275
rect 9933 18248 10012 18275
rect 9933 18244 9950 18248
rect 9933 18241 9945 18244
rect 9887 18235 9945 18241
rect 2700 18176 2774 18204
rect 2746 18068 2774 18176
rect 6730 18164 6736 18216
rect 6788 18164 6794 18216
rect 6825 18139 6883 18145
rect 6825 18105 6837 18139
rect 6871 18136 6883 18139
rect 7006 18136 7012 18148
rect 6871 18108 7012 18136
rect 6871 18105 6883 18108
rect 6825 18099 6883 18105
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 9140 18136 9168 18235
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 9692 18204 9720 18235
rect 9364 18176 9720 18204
rect 9784 18204 9812 18235
rect 9784 18176 9904 18204
rect 9364 18164 9370 18176
rect 9876 18148 9904 18176
rect 9766 18136 9772 18148
rect 9140 18108 9772 18136
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 9858 18096 9864 18148
rect 9916 18096 9922 18148
rect 3694 18068 3700 18080
rect 2746 18040 3700 18068
rect 3694 18028 3700 18040
rect 3752 18028 3758 18080
rect 6914 18028 6920 18080
rect 6972 18028 6978 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9582 18068 9588 18080
rect 9447 18040 9588 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 9984 18068 10012 18248
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18241 10379 18275
rect 10321 18235 10379 18241
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 10152 18204 10180 18235
rect 11422 18232 11428 18284
rect 11480 18272 11486 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11480 18244 11897 18272
rect 11480 18232 11486 18244
rect 11885 18241 11897 18244
rect 11931 18241 11943 18275
rect 11992 18272 12020 18312
rect 12066 18300 12072 18352
rect 12124 18340 12130 18352
rect 14292 18340 14320 18368
rect 12124 18312 14320 18340
rect 12124 18300 12130 18312
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 11992 18244 12817 18272
rect 11885 18235 11943 18241
rect 12805 18241 12817 18244
rect 12851 18272 12863 18275
rect 12851 18244 13492 18272
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 13464 18216 13492 18244
rect 13998 18232 14004 18284
rect 14056 18232 14062 18284
rect 14182 18232 14188 18284
rect 14240 18232 14246 18284
rect 14476 18272 14504 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 24394 18408 24400 18420
rect 24228 18380 24400 18408
rect 24228 18349 24256 18380
rect 24394 18368 24400 18380
rect 24452 18368 24458 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 25777 18411 25835 18417
rect 25777 18408 25789 18411
rect 24636 18380 25789 18408
rect 24636 18368 24642 18380
rect 25777 18377 25789 18380
rect 25823 18377 25835 18411
rect 25777 18371 25835 18377
rect 26234 18368 26240 18420
rect 26292 18368 26298 18420
rect 27908 18380 28396 18408
rect 24213 18343 24271 18349
rect 14936 18312 16068 18340
rect 14292 18244 14504 18272
rect 14553 18275 14611 18281
rect 10505 18207 10563 18213
rect 10505 18204 10517 18207
rect 10152 18176 10517 18204
rect 10152 18148 10180 18176
rect 10505 18173 10517 18176
rect 10551 18173 10563 18207
rect 10505 18167 10563 18173
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 11839 18176 11928 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 10134 18096 10140 18148
rect 10192 18096 10198 18148
rect 10594 18096 10600 18148
rect 10652 18136 10658 18148
rect 10781 18139 10839 18145
rect 10781 18136 10793 18139
rect 10652 18108 10793 18136
rect 10652 18096 10658 18108
rect 10781 18105 10793 18108
rect 10827 18105 10839 18139
rect 11517 18139 11575 18145
rect 11517 18136 11529 18139
rect 10781 18099 10839 18105
rect 10888 18108 11529 18136
rect 10888 18068 10916 18108
rect 11517 18105 11529 18108
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 11900 18080 11928 18176
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12676 18176 12909 18204
rect 12676 18164 12682 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 13446 18164 13452 18216
rect 13504 18164 13510 18216
rect 14016 18204 14044 18232
rect 14292 18204 14320 18244
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14016 18176 14320 18204
rect 14458 18164 14464 18216
rect 14516 18164 14522 18216
rect 14568 18204 14596 18235
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 14936 18281 14964 18312
rect 16040 18281 16068 18312
rect 20916 18312 23428 18340
rect 20916 18284 20944 18312
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14884 18244 14933 18272
rect 14884 18232 14890 18244
rect 14921 18241 14933 18244
rect 14967 18241 14979 18275
rect 14921 18235 14979 18241
rect 15197 18275 15255 18281
rect 15197 18241 15209 18275
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18241 15899 18275
rect 15841 18235 15899 18241
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16945 18275 17003 18281
rect 16945 18241 16957 18275
rect 16991 18272 17003 18275
rect 17218 18272 17224 18284
rect 16991 18244 17224 18272
rect 16991 18241 17003 18244
rect 16945 18235 17003 18241
rect 15212 18204 15240 18235
rect 14568 18176 15240 18204
rect 14568 18136 14596 18176
rect 14108 18108 14596 18136
rect 14108 18080 14136 18108
rect 15010 18096 15016 18148
rect 15068 18136 15074 18148
rect 15856 18136 15884 18235
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 19444 18244 19717 18272
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 17586 18204 17592 18216
rect 15988 18176 17592 18204
rect 15988 18164 15994 18176
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 17770 18136 17776 18148
rect 15068 18108 17776 18136
rect 15068 18096 15074 18108
rect 17770 18096 17776 18108
rect 17828 18096 17834 18148
rect 19444 18080 19472 18244
rect 19705 18241 19717 18244
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20530 18272 20536 18284
rect 20027 18244 20536 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20530 18232 20536 18244
rect 20588 18272 20594 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20588 18244 20821 18272
rect 20588 18232 20594 18244
rect 20809 18241 20821 18244
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 20128 18176 20269 18204
rect 20128 18164 20134 18176
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 20824 18204 20852 18235
rect 20898 18232 20904 18284
rect 20956 18232 20962 18284
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 22204 18281 22232 18312
rect 23400 18284 23428 18312
rect 24213 18309 24225 18343
rect 24259 18309 24271 18343
rect 24213 18303 24271 18309
rect 24854 18300 24860 18352
rect 24912 18300 24918 18352
rect 27338 18340 27344 18352
rect 27264 18312 27344 18340
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 21048 18244 21189 18272
rect 21048 18232 21054 18244
rect 21177 18241 21189 18244
rect 21223 18272 21235 18275
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21223 18244 21833 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22465 18275 22523 18281
rect 22235 18244 22269 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 22465 18241 22477 18275
rect 22511 18241 22523 18275
rect 22465 18235 22523 18241
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18272 22891 18275
rect 22922 18272 22928 18284
rect 22879 18244 22928 18272
rect 22879 18241 22891 18244
rect 22833 18235 22891 18241
rect 22480 18204 22508 18235
rect 22922 18232 22928 18244
rect 22980 18232 22986 18284
rect 23014 18232 23020 18284
rect 23072 18232 23078 18284
rect 23382 18232 23388 18284
rect 23440 18232 23446 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 26142 18272 26148 18284
rect 25700 18244 26148 18272
rect 23032 18204 23060 18232
rect 20824 18176 23060 18204
rect 20257 18167 20315 18173
rect 25406 18164 25412 18216
rect 25464 18164 25470 18216
rect 25700 18213 25728 18244
rect 26142 18232 26148 18244
rect 26200 18232 26206 18284
rect 26786 18232 26792 18284
rect 26844 18272 26850 18284
rect 27264 18281 27292 18312
rect 27338 18300 27344 18312
rect 27396 18340 27402 18352
rect 27908 18340 27936 18380
rect 27396 18312 27936 18340
rect 27396 18300 27402 18312
rect 27982 18300 27988 18352
rect 28040 18340 28046 18352
rect 28077 18343 28135 18349
rect 28077 18340 28089 18343
rect 28040 18312 28089 18340
rect 28040 18300 28046 18312
rect 28077 18309 28089 18312
rect 28123 18309 28135 18343
rect 28077 18303 28135 18309
rect 28166 18300 28172 18352
rect 28224 18340 28230 18352
rect 28277 18343 28335 18349
rect 28277 18340 28289 18343
rect 28224 18312 28289 18340
rect 28224 18300 28230 18312
rect 28277 18309 28289 18312
rect 28323 18309 28335 18343
rect 28368 18340 28396 18380
rect 28442 18368 28448 18420
rect 28500 18368 28506 18420
rect 29178 18368 29184 18420
rect 29236 18368 29242 18420
rect 28626 18340 28632 18352
rect 28368 18312 28632 18340
rect 28277 18303 28335 18309
rect 28626 18300 28632 18312
rect 28684 18300 28690 18352
rect 30098 18340 30104 18352
rect 29196 18312 30104 18340
rect 29196 18284 29224 18312
rect 30098 18300 30104 18312
rect 30156 18300 30162 18352
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 26844 18244 26985 18272
rect 26844 18232 26850 18244
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 27249 18275 27307 18281
rect 27249 18241 27261 18275
rect 27295 18241 27307 18275
rect 27249 18235 27307 18241
rect 29178 18232 29184 18284
rect 29236 18232 29242 18284
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18272 29423 18275
rect 30006 18272 30012 18284
rect 29411 18244 30012 18272
rect 29411 18241 29423 18244
rect 29365 18235 29423 18241
rect 30006 18232 30012 18244
rect 30064 18232 30070 18284
rect 25685 18207 25743 18213
rect 25685 18173 25697 18207
rect 25731 18173 25743 18207
rect 26050 18204 26056 18216
rect 25685 18167 25743 18173
rect 25792 18176 26056 18204
rect 25424 18136 25452 18164
rect 25792 18136 25820 18176
rect 26050 18164 26056 18176
rect 26108 18204 26114 18216
rect 26329 18207 26387 18213
rect 26329 18204 26341 18207
rect 26108 18176 26341 18204
rect 26108 18164 26114 18176
rect 26329 18173 26341 18176
rect 26375 18173 26387 18207
rect 26329 18167 26387 18173
rect 25424 18108 25820 18136
rect 27540 18108 28304 18136
rect 27540 18080 27568 18108
rect 9984 18040 10916 18068
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11054 18068 11060 18080
rect 11011 18040 11060 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11882 18028 11888 18080
rect 11940 18028 11946 18080
rect 14090 18028 14096 18080
rect 14148 18028 14154 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16761 18071 16819 18077
rect 16761 18068 16773 18071
rect 16632 18040 16773 18068
rect 16632 18028 16638 18040
rect 16761 18037 16773 18040
rect 16807 18037 16819 18071
rect 16761 18031 16819 18037
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 19242 18068 19248 18080
rect 18012 18040 19248 18068
rect 18012 18028 18018 18040
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19426 18028 19432 18080
rect 19484 18028 19490 18080
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20680 18040 20729 18068
rect 20680 18028 20686 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 22557 18071 22615 18077
rect 22557 18037 22569 18071
rect 22603 18068 22615 18071
rect 23474 18068 23480 18080
rect 22603 18040 23480 18068
rect 22603 18037 22615 18040
rect 22557 18031 22615 18037
rect 23474 18028 23480 18040
rect 23532 18028 23538 18080
rect 27522 18028 27528 18080
rect 27580 18028 27586 18080
rect 27985 18071 28043 18077
rect 27985 18037 27997 18071
rect 28031 18068 28043 18071
rect 28074 18068 28080 18080
rect 28031 18040 28080 18068
rect 28031 18037 28043 18040
rect 27985 18031 28043 18037
rect 28074 18028 28080 18040
rect 28132 18028 28138 18080
rect 28276 18077 28304 18108
rect 28261 18071 28319 18077
rect 28261 18037 28273 18071
rect 28307 18037 28319 18071
rect 28261 18031 28319 18037
rect 1104 17978 30820 18000
rect 1104 17926 4664 17978
rect 4716 17926 4728 17978
rect 4780 17926 4792 17978
rect 4844 17926 4856 17978
rect 4908 17926 4920 17978
rect 4972 17926 12092 17978
rect 12144 17926 12156 17978
rect 12208 17926 12220 17978
rect 12272 17926 12284 17978
rect 12336 17926 12348 17978
rect 12400 17926 19520 17978
rect 19572 17926 19584 17978
rect 19636 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 26948 17978
rect 27000 17926 27012 17978
rect 27064 17926 27076 17978
rect 27128 17926 27140 17978
rect 27192 17926 27204 17978
rect 27256 17926 30820 17978
rect 1104 17904 30820 17926
rect 6365 17867 6423 17873
rect 6365 17833 6377 17867
rect 6411 17864 6423 17867
rect 6454 17864 6460 17876
rect 6411 17836 6460 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6549 17867 6607 17873
rect 6549 17833 6561 17867
rect 6595 17864 6607 17867
rect 6730 17864 6736 17876
rect 6595 17836 6736 17864
rect 6595 17833 6607 17836
rect 6549 17827 6607 17833
rect 5537 17731 5595 17737
rect 5537 17697 5549 17731
rect 5583 17697 5595 17731
rect 5537 17691 5595 17697
rect 3786 17620 3792 17672
rect 3844 17620 3850 17672
rect 5552 17660 5580 17691
rect 5718 17660 5724 17672
rect 5552 17632 5724 17660
rect 5718 17620 5724 17632
rect 5776 17660 5782 17672
rect 6656 17669 6684 17836
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 9858 17864 9864 17876
rect 8352 17836 9864 17864
rect 8352 17824 8358 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 10502 17824 10508 17876
rect 10560 17824 10566 17876
rect 11054 17824 11060 17876
rect 11112 17824 11118 17876
rect 11422 17824 11428 17876
rect 11480 17824 11486 17876
rect 15028 17836 18644 17864
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 7282 17796 7288 17808
rect 6972 17768 7288 17796
rect 6972 17756 6978 17768
rect 7208 17737 7236 17768
rect 7282 17756 7288 17768
rect 7340 17796 7346 17808
rect 11517 17799 11575 17805
rect 11517 17796 11529 17799
rect 7340 17768 11529 17796
rect 7340 17756 7346 17768
rect 11517 17765 11529 17768
rect 11563 17765 11575 17799
rect 11517 17759 11575 17765
rect 12342 17756 12348 17808
rect 12400 17796 12406 17808
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12400 17768 13001 17796
rect 12400 17756 12406 17768
rect 12989 17765 13001 17768
rect 13035 17765 13047 17799
rect 12989 17759 13047 17765
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 7469 17731 7527 17737
rect 7469 17697 7481 17731
rect 7515 17728 7527 17731
rect 8481 17731 8539 17737
rect 7515 17700 8340 17728
rect 7515 17697 7527 17700
rect 7469 17691 7527 17697
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 5776 17632 6101 17660
rect 5776 17620 5782 17632
rect 6089 17629 6101 17632
rect 6135 17660 6147 17663
rect 6641 17663 6699 17669
rect 6135 17632 6500 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 4062 17552 4068 17604
rect 4120 17552 4126 17604
rect 4522 17552 4528 17604
rect 4580 17552 4586 17604
rect 6472 17536 6500 17632
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 6822 17620 6828 17672
rect 6880 17620 6886 17672
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17629 8079 17663
rect 8021 17623 8079 17629
rect 6733 17595 6791 17601
rect 6733 17561 6745 17595
rect 6779 17592 6791 17595
rect 7116 17592 7144 17623
rect 7190 17592 7196 17604
rect 6779 17564 7196 17592
rect 6779 17561 6791 17564
rect 6733 17555 6791 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 6454 17484 6460 17536
rect 6512 17484 6518 17536
rect 7834 17484 7840 17536
rect 7892 17484 7898 17536
rect 8036 17524 8064 17623
rect 8202 17620 8208 17672
rect 8260 17620 8266 17672
rect 8312 17669 8340 17700
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8846 17728 8852 17740
rect 8527 17700 8852 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8846 17688 8852 17700
rect 8904 17728 8910 17740
rect 10042 17728 10048 17740
rect 8904 17700 10048 17728
rect 8904 17688 8910 17700
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 10873 17731 10931 17737
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 10919 17700 11008 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 8312 17663 8381 17669
rect 8312 17632 8335 17663
rect 8323 17629 8335 17632
rect 8369 17629 8381 17663
rect 8323 17623 8381 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 8662 17660 8668 17672
rect 8619 17632 8668 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17660 8815 17663
rect 9306 17660 9312 17672
rect 8803 17632 9312 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 10134 17660 10140 17672
rect 9824 17632 10140 17660
rect 9824 17620 9830 17632
rect 10134 17620 10140 17632
rect 10192 17660 10198 17672
rect 10980 17669 11008 17700
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10192 17632 10425 17660
rect 10192 17620 10198 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11011 17632 11713 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 11793 17663 11851 17669
rect 11793 17629 11805 17663
rect 11839 17660 11851 17663
rect 11839 17632 11928 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 8113 17595 8171 17601
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8478 17592 8484 17604
rect 8159 17564 8484 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8478 17552 8484 17564
rect 8536 17592 8542 17604
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 8536 17564 8953 17592
rect 8536 17552 8542 17564
rect 8941 17561 8953 17564
rect 8987 17561 8999 17595
rect 8941 17555 8999 17561
rect 9125 17595 9183 17601
rect 9125 17561 9137 17595
rect 9171 17561 9183 17595
rect 9125 17555 9183 17561
rect 8573 17527 8631 17533
rect 8573 17524 8585 17527
rect 8036 17496 8585 17524
rect 8573 17493 8585 17496
rect 8619 17493 8631 17527
rect 8573 17487 8631 17493
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 9140 17524 9168 17555
rect 11054 17552 11060 17604
rect 11112 17592 11118 17604
rect 11517 17595 11575 17601
rect 11517 17592 11529 17595
rect 11112 17564 11529 17592
rect 11112 17552 11118 17564
rect 11517 17561 11529 17564
rect 11563 17561 11575 17595
rect 11517 17555 11575 17561
rect 11900 17536 11928 17632
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12124 17632 12817 17660
rect 12124 17620 12130 17632
rect 12805 17629 12817 17632
rect 12851 17660 12863 17663
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 12851 17632 13185 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 13173 17629 13185 17632
rect 13219 17660 13231 17663
rect 14734 17660 14740 17672
rect 13219 17632 14740 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 14734 17620 14740 17632
rect 14792 17660 14798 17672
rect 15028 17660 15056 17836
rect 17954 17756 17960 17808
rect 18012 17756 18018 17808
rect 18616 17796 18644 17836
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19061 17867 19119 17873
rect 19061 17864 19073 17867
rect 19024 17836 19073 17864
rect 19024 17824 19030 17836
rect 19061 17833 19073 17836
rect 19107 17833 19119 17867
rect 19061 17827 19119 17833
rect 19150 17824 19156 17876
rect 19208 17864 19214 17876
rect 19886 17864 19892 17876
rect 19208 17836 19892 17864
rect 19208 17824 19214 17836
rect 19886 17824 19892 17836
rect 19944 17824 19950 17876
rect 20548 17836 22094 17864
rect 20162 17796 20168 17808
rect 18616 17768 20168 17796
rect 20162 17756 20168 17768
rect 20220 17756 20226 17808
rect 15654 17688 15660 17740
rect 15712 17728 15718 17740
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15712 17700 16221 17728
rect 15712 17688 15718 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16209 17691 16267 17697
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 16574 17728 16580 17740
rect 16531 17700 16580 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 16574 17688 16580 17700
rect 16632 17688 16638 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19168 17700 19717 17728
rect 14792 17632 15056 17660
rect 18049 17663 18107 17669
rect 14792 17620 14798 17632
rect 18049 17629 18061 17663
rect 18095 17660 18107 17663
rect 18325 17663 18383 17669
rect 18095 17632 18184 17660
rect 18095 17629 18107 17632
rect 18049 17623 18107 17629
rect 12618 17552 12624 17604
rect 12676 17552 12682 17604
rect 17034 17552 17040 17604
rect 17092 17552 17098 17604
rect 18156 17592 18184 17632
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 19168 17660 19196 17700
rect 19705 17697 19717 17700
rect 19751 17728 19763 17731
rect 20548 17728 20576 17836
rect 22066 17796 22094 17836
rect 24854 17824 24860 17876
rect 24912 17824 24918 17876
rect 27430 17824 27436 17876
rect 27488 17864 27494 17876
rect 27525 17867 27583 17873
rect 27525 17864 27537 17867
rect 27488 17836 27537 17864
rect 27488 17824 27494 17836
rect 27525 17833 27537 17836
rect 27571 17833 27583 17867
rect 27525 17827 27583 17833
rect 27614 17824 27620 17876
rect 27672 17824 27678 17876
rect 28077 17867 28135 17873
rect 28077 17833 28089 17867
rect 28123 17864 28135 17867
rect 28166 17864 28172 17876
rect 28123 17836 28172 17864
rect 28123 17833 28135 17836
rect 28077 17827 28135 17833
rect 28166 17824 28172 17836
rect 28224 17824 28230 17876
rect 28813 17867 28871 17873
rect 28813 17833 28825 17867
rect 28859 17833 28871 17867
rect 28813 17827 28871 17833
rect 27632 17796 27660 17824
rect 28828 17796 28856 17827
rect 29178 17824 29184 17876
rect 29236 17824 29242 17876
rect 29641 17867 29699 17873
rect 29641 17833 29653 17867
rect 29687 17833 29699 17867
rect 29641 17827 29699 17833
rect 22066 17768 27660 17796
rect 28184 17768 28856 17796
rect 19751 17700 20576 17728
rect 22557 17731 22615 17737
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 22557 17697 22569 17731
rect 22603 17728 22615 17731
rect 22922 17728 22928 17740
rect 22603 17700 22928 17728
rect 22603 17697 22615 17700
rect 22557 17691 22615 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23385 17731 23443 17737
rect 23385 17697 23397 17731
rect 23431 17728 23443 17731
rect 25777 17731 25835 17737
rect 25777 17728 25789 17731
rect 23431 17700 25789 17728
rect 23431 17697 23443 17700
rect 23385 17691 23443 17697
rect 25777 17697 25789 17700
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 27338 17688 27344 17740
rect 27396 17688 27402 17740
rect 18371 17632 19196 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 23014 17620 23020 17672
rect 23072 17620 23078 17672
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17660 23351 17663
rect 23339 17632 23428 17660
rect 23339 17629 23351 17632
rect 23293 17623 23351 17629
rect 23400 17604 23428 17632
rect 23566 17620 23572 17672
rect 23624 17620 23630 17672
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 25038 17660 25044 17672
rect 24811 17632 25044 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 25593 17663 25651 17669
rect 25593 17629 25605 17663
rect 25639 17629 25651 17663
rect 25593 17623 25651 17629
rect 27893 17663 27951 17669
rect 27893 17629 27905 17663
rect 27939 17660 27951 17663
rect 27982 17660 27988 17672
rect 27939 17632 27988 17660
rect 27939 17629 27951 17632
rect 27893 17623 27951 17629
rect 19429 17595 19487 17601
rect 18156 17564 19380 17592
rect 19352 17536 19380 17564
rect 19429 17561 19441 17595
rect 19475 17592 19487 17595
rect 19475 17564 19932 17592
rect 19475 17561 19487 17564
rect 19429 17555 19487 17561
rect 19904 17536 19932 17564
rect 23382 17552 23388 17604
rect 23440 17552 23446 17604
rect 25608 17592 25636 17623
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28184 17669 28212 17768
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28721 17663 28779 17669
rect 28721 17629 28733 17663
rect 28767 17629 28779 17663
rect 28828 17660 28856 17768
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 28828 17632 29561 17660
rect 28721 17623 28779 17629
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 27709 17595 27767 17601
rect 25608 17564 26188 17592
rect 26160 17536 26188 17564
rect 27709 17561 27721 17595
rect 27755 17592 27767 17595
rect 28074 17592 28080 17604
rect 27755 17564 28080 17592
rect 27755 17561 27767 17564
rect 27709 17555 27767 17561
rect 28074 17552 28080 17564
rect 28132 17592 28138 17604
rect 28184 17592 28212 17623
rect 28132 17564 28212 17592
rect 28736 17592 28764 17623
rect 29656 17592 29684 17827
rect 30006 17824 30012 17876
rect 30064 17824 30070 17876
rect 28736 17564 29684 17592
rect 28132 17552 28138 17564
rect 8720 17496 9168 17524
rect 8720 17484 8726 17496
rect 11882 17484 11888 17536
rect 11940 17484 11946 17536
rect 19334 17484 19340 17536
rect 19392 17484 19398 17536
rect 19886 17484 19892 17536
rect 19944 17484 19950 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 24026 17524 24032 17536
rect 20220 17496 24032 17524
rect 20220 17484 20226 17496
rect 24026 17484 24032 17496
rect 24084 17484 24090 17536
rect 26142 17484 26148 17536
rect 26200 17524 26206 17536
rect 28736 17524 28764 17564
rect 26200 17496 28764 17524
rect 26200 17484 26206 17496
rect 1104 17434 30820 17456
rect 1104 17382 5324 17434
rect 5376 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 12752 17434
rect 12804 17382 12816 17434
rect 12868 17382 12880 17434
rect 12932 17382 12944 17434
rect 12996 17382 13008 17434
rect 13060 17382 20180 17434
rect 20232 17382 20244 17434
rect 20296 17382 20308 17434
rect 20360 17382 20372 17434
rect 20424 17382 20436 17434
rect 20488 17382 27608 17434
rect 27660 17382 27672 17434
rect 27724 17382 27736 17434
rect 27788 17382 27800 17434
rect 27852 17382 27864 17434
rect 27916 17382 30820 17434
rect 1104 17360 30820 17382
rect 4062 17280 4068 17332
rect 4120 17320 4126 17332
rect 4157 17323 4215 17329
rect 4157 17320 4169 17323
rect 4120 17292 4169 17320
rect 4120 17280 4126 17292
rect 4157 17289 4169 17292
rect 4203 17289 4215 17323
rect 4157 17283 4215 17289
rect 4522 17280 4528 17332
rect 4580 17280 4586 17332
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17289 4767 17323
rect 4709 17283 4767 17289
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 5718 17320 5724 17332
rect 5123 17292 5724 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 4724 17252 4752 17283
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 6822 17280 6828 17332
rect 6880 17280 6886 17332
rect 7834 17280 7840 17332
rect 7892 17280 7898 17332
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 9677 17323 9735 17329
rect 9677 17320 9689 17323
rect 9640 17292 9689 17320
rect 9640 17280 9646 17292
rect 9677 17289 9689 17292
rect 9723 17289 9735 17323
rect 9677 17283 9735 17289
rect 12161 17323 12219 17329
rect 12161 17289 12173 17323
rect 12207 17320 12219 17323
rect 12618 17320 12624 17332
rect 12207 17292 12624 17320
rect 12207 17289 12219 17292
rect 12161 17283 12219 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 14826 17320 14832 17332
rect 13740 17292 14832 17320
rect 4356 17224 4752 17252
rect 5169 17255 5227 17261
rect 4356 17193 4384 17224
rect 5169 17221 5181 17255
rect 5215 17252 5227 17255
rect 7852 17252 7880 17280
rect 13740 17264 13768 17292
rect 14826 17280 14832 17292
rect 14884 17320 14890 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 14884 17292 15577 17320
rect 14884 17280 14890 17292
rect 15565 17289 15577 17292
rect 15611 17320 15623 17323
rect 15611 17292 16804 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 5215 17224 7880 17252
rect 5215 17221 5227 17224
rect 5169 17215 5227 17221
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 7984 17224 12664 17252
rect 7984 17212 7990 17224
rect 12636 17196 12664 17224
rect 13722 17212 13728 17264
rect 13780 17212 13786 17264
rect 14550 17212 14556 17264
rect 14608 17212 14614 17264
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4341 17147 4399 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4479 17156 6316 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4448 17116 4476 17147
rect 6288 17128 6316 17156
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7101 17187 7159 17193
rect 7101 17184 7113 17187
rect 6972 17156 7113 17184
rect 6972 17144 6978 17156
rect 7101 17153 7113 17156
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 9674 17184 9680 17196
rect 9631 17156 9680 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11112 17156 11529 17184
rect 11112 17144 11118 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 12066 17184 12072 17196
rect 11517 17147 11575 17153
rect 11624 17156 12072 17184
rect 4120 17088 4476 17116
rect 4120 17076 4126 17088
rect 5258 17076 5264 17128
rect 5316 17076 5322 17128
rect 6270 17076 6276 17128
rect 6328 17076 6334 17128
rect 7116 17088 7420 17116
rect 4338 17008 4344 17060
rect 4396 17048 4402 17060
rect 7116 17048 7144 17088
rect 4396 17020 7144 17048
rect 7392 17048 7420 17088
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 8168 17088 9781 17116
rect 8168 17076 8174 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 11624 17048 11652 17156
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 7392 17020 11652 17048
rect 11808 17048 11836 17079
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12268 17116 12296 17147
rect 12342 17144 12348 17196
rect 12400 17144 12406 17196
rect 12618 17144 12624 17196
rect 12676 17144 12682 17196
rect 13446 17144 13452 17196
rect 13504 17144 13510 17196
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 15304 17156 15485 17184
rect 12032 17088 12296 17116
rect 12032 17076 12038 17088
rect 13538 17076 13544 17128
rect 13596 17076 13602 17128
rect 13814 17076 13820 17128
rect 13872 17076 13878 17128
rect 15304 17125 15332 17156
rect 15473 17153 15485 17156
rect 15519 17184 15531 17187
rect 15562 17184 15568 17196
rect 15519 17156 15568 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15896 17156 16037 17184
rect 15896 17144 15902 17156
rect 16025 17153 16037 17156
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 16776 17048 16804 17292
rect 16850 17280 16856 17332
rect 16908 17280 16914 17332
rect 17034 17280 17040 17332
rect 17092 17280 17098 17332
rect 17218 17280 17224 17332
rect 17276 17280 17282 17332
rect 17681 17323 17739 17329
rect 17681 17289 17693 17323
rect 17727 17320 17739 17323
rect 17862 17320 17868 17332
rect 17727 17292 17868 17320
rect 17727 17289 17739 17292
rect 17681 17283 17739 17289
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 17954 17280 17960 17332
rect 18012 17280 18018 17332
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 21082 17320 21088 17332
rect 19392 17292 21088 17320
rect 19392 17280 19398 17292
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 24946 17320 24952 17332
rect 23676 17292 24952 17320
rect 16868 17184 16896 17280
rect 17589 17255 17647 17261
rect 17589 17221 17601 17255
rect 17635 17252 17647 17255
rect 17972 17252 18000 17280
rect 17635 17224 18000 17252
rect 17635 17221 17647 17224
rect 17589 17215 17647 17221
rect 19886 17212 19892 17264
rect 19944 17252 19950 17264
rect 20349 17255 20407 17261
rect 20349 17252 20361 17255
rect 19944 17224 20361 17252
rect 19944 17212 19950 17224
rect 20349 17221 20361 17224
rect 20395 17221 20407 17255
rect 20349 17215 20407 17221
rect 23474 17212 23480 17264
rect 23532 17212 23538 17264
rect 23676 17196 23704 17292
rect 24946 17280 24952 17292
rect 25004 17320 25010 17332
rect 25501 17323 25559 17329
rect 25501 17320 25513 17323
rect 25004 17292 25513 17320
rect 25004 17280 25010 17292
rect 25501 17289 25513 17292
rect 25547 17289 25559 17323
rect 25501 17283 25559 17289
rect 26418 17280 26424 17332
rect 26476 17320 26482 17332
rect 27341 17323 27399 17329
rect 27341 17320 27353 17323
rect 26476 17292 27353 17320
rect 26476 17280 26482 17292
rect 27341 17289 27353 17292
rect 27387 17289 27399 17323
rect 27341 17283 27399 17289
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 16868 17156 16957 17184
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 18322 17144 18328 17196
rect 18380 17184 18386 17196
rect 19337 17187 19395 17193
rect 19337 17184 19349 17187
rect 18380 17156 19349 17184
rect 18380 17144 18386 17156
rect 19337 17153 19349 17156
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17184 19579 17187
rect 20070 17184 20076 17196
rect 19567 17156 20076 17184
rect 19567 17153 19579 17156
rect 19521 17147 19579 17153
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20530 17144 20536 17196
rect 20588 17144 20594 17196
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 20898 17184 20904 17196
rect 20855 17156 20904 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 20990 17144 20996 17196
rect 21048 17144 21054 17196
rect 23658 17144 23664 17196
rect 23716 17144 23722 17196
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 25130 17144 25136 17196
rect 25188 17144 25194 17196
rect 27522 17144 27528 17196
rect 27580 17144 27586 17196
rect 27801 17187 27859 17193
rect 27801 17153 27813 17187
rect 27847 17184 27859 17187
rect 28166 17184 28172 17196
rect 27847 17156 28172 17184
rect 27847 17153 27859 17156
rect 27801 17147 27859 17153
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 17865 17119 17923 17125
rect 17865 17085 17877 17119
rect 17911 17116 17923 17119
rect 23109 17119 23167 17125
rect 17911 17088 19932 17116
rect 17911 17085 17923 17088
rect 17865 17079 17923 17085
rect 18322 17048 18328 17060
rect 11808 17020 12434 17048
rect 16776 17020 18328 17048
rect 4396 17008 4402 17020
rect 6454 16940 6460 16992
rect 6512 16940 6518 16992
rect 7282 16940 7288 16992
rect 7340 16940 7346 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7469 16983 7527 16989
rect 7469 16980 7481 16983
rect 7432 16952 7481 16980
rect 7432 16940 7438 16952
rect 7469 16949 7481 16952
rect 7515 16949 7527 16983
rect 7469 16943 7527 16949
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 9088 16952 9229 16980
rect 9088 16940 9094 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 12250 16980 12256 16992
rect 11296 16952 12256 16980
rect 11296 16940 11302 16952
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12406 16980 12434 17020
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 19904 16992 19932 17088
rect 23109 17085 23121 17119
rect 23155 17085 23167 17119
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23109 17079 23167 17085
rect 23768 17088 24041 17116
rect 23124 16992 23152 17079
rect 23198 17008 23204 17060
rect 23256 17048 23262 17060
rect 23768 17048 23796 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17116 27767 17119
rect 28258 17116 28264 17128
rect 27755 17088 28264 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 28258 17076 28264 17088
rect 28316 17076 28322 17128
rect 27798 17048 27804 17060
rect 23256 17020 23796 17048
rect 25056 17020 27804 17048
rect 23256 17008 23262 17020
rect 13262 16980 13268 16992
rect 12406 16952 13268 16980
rect 13262 16940 13268 16952
rect 13320 16940 13326 16992
rect 13998 16940 14004 16992
rect 14056 16980 14062 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 14056 16952 16129 16980
rect 14056 16940 14062 16952
rect 16117 16949 16129 16952
rect 16163 16980 16175 16983
rect 17034 16980 17040 16992
rect 16163 16952 17040 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 23014 16980 23020 16992
rect 19944 16952 23020 16980
rect 19944 16940 19950 16952
rect 23014 16940 23020 16952
rect 23072 16940 23078 16992
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 25056 16980 25084 17020
rect 27798 17008 27804 17020
rect 27856 17008 27862 17060
rect 23164 16952 25084 16980
rect 27709 16983 27767 16989
rect 23164 16940 23170 16952
rect 27709 16949 27721 16983
rect 27755 16980 27767 16983
rect 28074 16980 28080 16992
rect 27755 16952 28080 16980
rect 27755 16949 27767 16952
rect 27709 16943 27767 16949
rect 28074 16940 28080 16952
rect 28132 16940 28138 16992
rect 1104 16890 30820 16912
rect 1104 16838 4664 16890
rect 4716 16838 4728 16890
rect 4780 16838 4792 16890
rect 4844 16838 4856 16890
rect 4908 16838 4920 16890
rect 4972 16838 12092 16890
rect 12144 16838 12156 16890
rect 12208 16838 12220 16890
rect 12272 16838 12284 16890
rect 12336 16838 12348 16890
rect 12400 16838 19520 16890
rect 19572 16838 19584 16890
rect 19636 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 26948 16890
rect 27000 16838 27012 16890
rect 27064 16838 27076 16890
rect 27128 16838 27140 16890
rect 27192 16838 27204 16890
rect 27256 16838 30820 16890
rect 1104 16816 30820 16838
rect 5258 16736 5264 16788
rect 5316 16776 5322 16788
rect 8110 16776 8116 16788
rect 5316 16748 8116 16776
rect 5316 16736 5322 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 9582 16776 9588 16788
rect 8220 16748 9588 16776
rect 5718 16708 5724 16720
rect 4264 16680 5724 16708
rect 4264 16649 4292 16680
rect 5718 16668 5724 16680
rect 5776 16668 5782 16720
rect 5813 16711 5871 16717
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 6178 16708 6184 16720
rect 5859 16680 6184 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 6270 16668 6276 16720
rect 6328 16708 6334 16720
rect 8220 16708 8248 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 10502 16776 10508 16788
rect 9732 16748 10508 16776
rect 9732 16736 9738 16748
rect 10502 16736 10508 16748
rect 10560 16776 10566 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10560 16748 10977 16776
rect 10560 16736 10566 16748
rect 10965 16745 10977 16748
rect 11011 16745 11023 16779
rect 10965 16739 11023 16745
rect 11701 16779 11759 16785
rect 11701 16745 11713 16779
rect 11747 16745 11759 16779
rect 11701 16739 11759 16745
rect 6328 16680 8248 16708
rect 11716 16708 11744 16739
rect 11882 16736 11888 16788
rect 11940 16736 11946 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13872 16748 14105 16776
rect 13872 16736 13878 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14608 16748 14657 16776
rect 14608 16736 14614 16748
rect 14645 16745 14657 16748
rect 14691 16745 14703 16779
rect 14645 16739 14703 16745
rect 15194 16736 15200 16788
rect 15252 16736 15258 16788
rect 15286 16736 15292 16788
rect 15344 16736 15350 16788
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 18874 16776 18880 16788
rect 18472 16748 18880 16776
rect 18472 16736 18478 16748
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19886 16776 19892 16788
rect 19015 16748 19892 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 20530 16736 20536 16788
rect 20588 16776 20594 16788
rect 21082 16776 21088 16788
rect 20588 16748 21088 16776
rect 20588 16736 20594 16748
rect 21082 16736 21088 16748
rect 21140 16776 21146 16788
rect 26786 16776 26792 16788
rect 21140 16748 26792 16776
rect 21140 16736 21146 16748
rect 11790 16708 11796 16720
rect 11716 16680 11796 16708
rect 6328 16668 6334 16680
rect 11790 16668 11796 16680
rect 11848 16708 11854 16720
rect 11848 16680 12112 16708
rect 11848 16668 11854 16680
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16609 4307 16643
rect 4249 16603 4307 16609
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4522 16640 4528 16652
rect 4479 16612 4528 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4522 16600 4528 16612
rect 4580 16640 4586 16652
rect 5258 16640 5264 16652
rect 4580 16612 5264 16640
rect 4580 16600 4586 16612
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 6914 16600 6920 16652
rect 6972 16600 6978 16652
rect 9217 16643 9275 16649
rect 8496 16612 9168 16640
rect 7006 16532 7012 16584
rect 7064 16532 7070 16584
rect 8496 16581 8524 16612
rect 9140 16584 9168 16612
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 9490 16640 9496 16652
rect 9263 16612 9496 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 11146 16640 11152 16652
rect 9640 16612 11152 16640
rect 9640 16600 9646 16612
rect 8481 16575 8539 16581
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8570 16532 8576 16584
rect 8628 16572 8634 16584
rect 8665 16575 8723 16581
rect 8665 16572 8677 16575
rect 8628 16544 8677 16572
rect 8628 16532 8634 16544
rect 8665 16541 8677 16544
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16572 8999 16575
rect 9030 16572 9036 16584
rect 8987 16544 9036 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 9122 16532 9128 16584
rect 9180 16532 9186 16584
rect 11072 16581 11100 16612
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 12084 16649 12112 16680
rect 12069 16643 12127 16649
rect 11440 16612 11928 16640
rect 11440 16581 11468 16612
rect 11057 16575 11115 16581
rect 11057 16541 11069 16575
rect 11103 16541 11115 16575
rect 11057 16535 11115 16541
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 5166 16504 5172 16516
rect 4172 16476 5172 16504
rect 4172 16448 4200 16476
rect 5166 16464 5172 16476
rect 5224 16504 5230 16516
rect 5445 16507 5503 16513
rect 5445 16504 5457 16507
rect 5224 16476 5457 16504
rect 5224 16464 5230 16476
rect 5445 16473 5457 16476
rect 5491 16473 5503 16507
rect 8386 16504 8392 16516
rect 5445 16467 5503 16473
rect 7392 16476 8392 16504
rect 2682 16396 2688 16448
rect 2740 16436 2746 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 2740 16408 3801 16436
rect 2740 16396 2746 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4154 16396 4160 16448
rect 4212 16396 4218 16448
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16436 5963 16439
rect 6546 16436 6552 16448
rect 5951 16408 6552 16436
rect 5951 16405 5963 16408
rect 5905 16399 5963 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 7392 16445 7420 16476
rect 8386 16464 8392 16476
rect 8444 16464 8450 16516
rect 9493 16507 9551 16513
rect 9493 16504 9505 16507
rect 9140 16476 9505 16504
rect 7377 16439 7435 16445
rect 7377 16405 7389 16439
rect 7423 16405 7435 16439
rect 7377 16399 7435 16405
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 9140 16445 9168 16476
rect 9493 16473 9505 16476
rect 9539 16473 9551 16507
rect 11149 16507 11207 16513
rect 11149 16504 11161 16507
rect 10718 16476 11161 16504
rect 9493 16467 9551 16473
rect 11149 16473 11161 16476
rect 11195 16473 11207 16507
rect 11149 16467 11207 16473
rect 11900 16448 11928 16612
rect 12069 16609 12081 16643
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12618 16600 12624 16652
rect 12676 16600 12682 16652
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 15212 16640 15240 16736
rect 17954 16668 17960 16720
rect 18012 16708 18018 16720
rect 18325 16711 18383 16717
rect 18325 16708 18337 16711
rect 18012 16680 18337 16708
rect 18012 16668 18018 16680
rect 18325 16677 18337 16680
rect 18371 16708 18383 16711
rect 19150 16708 19156 16720
rect 18371 16680 19156 16708
rect 18371 16677 18383 16680
rect 18325 16671 18383 16677
rect 19150 16668 19156 16680
rect 19208 16708 19214 16720
rect 20070 16708 20076 16720
rect 19208 16680 20076 16708
rect 19208 16668 19214 16680
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 13320 16612 15240 16640
rect 13320 16600 13326 16612
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 14568 16581 14596 16612
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15620 16612 15669 16640
rect 15620 16600 15626 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 19337 16643 19395 16649
rect 19337 16640 19349 16643
rect 15657 16603 15715 16609
rect 19168 16612 19349 16640
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15838 16572 15844 16584
rect 15519 16544 15844 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 19168 16572 19196 16612
rect 19337 16609 19349 16612
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 19521 16643 19579 16649
rect 19521 16609 19533 16643
rect 19567 16640 19579 16643
rect 19978 16640 19984 16652
rect 19567 16612 19984 16640
rect 19567 16609 19579 16612
rect 19521 16603 19579 16609
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20441 16643 20499 16649
rect 20441 16609 20453 16643
rect 20487 16640 20499 16643
rect 20990 16640 20996 16652
rect 20487 16612 20996 16640
rect 20487 16609 20499 16612
rect 20441 16603 20499 16609
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 21910 16600 21916 16652
rect 21968 16600 21974 16652
rect 22388 16649 22416 16748
rect 26786 16736 26792 16748
rect 26844 16736 26850 16788
rect 27982 16736 27988 16788
rect 28040 16776 28046 16788
rect 28629 16779 28687 16785
rect 28629 16776 28641 16779
rect 28040 16748 28641 16776
rect 28040 16736 28046 16748
rect 28629 16745 28641 16748
rect 28675 16745 28687 16779
rect 28629 16739 28687 16745
rect 23014 16668 23020 16720
rect 23072 16668 23078 16720
rect 23750 16668 23756 16720
rect 23808 16708 23814 16720
rect 23808 16680 24532 16708
rect 23808 16668 23814 16680
rect 22373 16643 22431 16649
rect 22373 16609 22385 16643
rect 22419 16609 22431 16643
rect 23032 16640 23060 16668
rect 24504 16649 24532 16680
rect 24121 16643 24179 16649
rect 24121 16640 24133 16643
rect 23032 16612 24133 16640
rect 22373 16603 22431 16609
rect 24121 16609 24133 16612
rect 24167 16640 24179 16643
rect 24489 16643 24547 16649
rect 24167 16612 24440 16640
rect 24167 16609 24179 16612
rect 24121 16603 24179 16609
rect 18840 16544 19196 16572
rect 19253 16575 19311 16581
rect 18840 16532 18846 16544
rect 19253 16541 19265 16575
rect 19299 16572 19311 16575
rect 22649 16575 22707 16581
rect 19299 16541 19334 16572
rect 19253 16535 19334 16541
rect 22649 16541 22661 16575
rect 22695 16572 22707 16575
rect 23106 16572 23112 16584
rect 22695 16544 23112 16572
rect 22695 16541 22707 16544
rect 22649 16535 22707 16541
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 12253 16507 12311 16513
rect 12253 16504 12265 16507
rect 12032 16476 12265 16504
rect 12032 16464 12038 16476
rect 12253 16473 12265 16476
rect 12299 16473 12311 16507
rect 12253 16467 12311 16473
rect 18138 16464 18144 16516
rect 18196 16464 18202 16516
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 18693 16507 18751 16513
rect 18693 16504 18705 16507
rect 18564 16476 18705 16504
rect 18564 16464 18570 16476
rect 18693 16473 18705 16476
rect 18739 16473 18751 16507
rect 18693 16467 18751 16473
rect 8481 16439 8539 16445
rect 8481 16436 8493 16439
rect 8168 16408 8493 16436
rect 8168 16396 8174 16408
rect 8481 16405 8493 16408
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16405 9183 16439
rect 9125 16399 9183 16405
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 13446 16436 13452 16448
rect 11940 16408 13452 16436
rect 11940 16396 11946 16408
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 18708 16436 18736 16467
rect 18874 16464 18880 16516
rect 18932 16504 18938 16516
rect 19306 16504 19334 16535
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 18932 16476 19840 16504
rect 18932 16464 18938 16476
rect 19705 16439 19763 16445
rect 19705 16436 19717 16439
rect 18708 16408 19717 16436
rect 19705 16405 19717 16408
rect 19751 16405 19763 16439
rect 19812 16436 19840 16476
rect 20622 16464 20628 16516
rect 20680 16464 20686 16516
rect 21082 16464 21088 16516
rect 21140 16504 21146 16516
rect 22002 16504 22008 16516
rect 21140 16476 22008 16504
rect 21140 16464 21146 16476
rect 22002 16464 22008 16476
rect 22060 16464 22066 16516
rect 23676 16504 23704 16532
rect 23845 16507 23903 16513
rect 23845 16504 23857 16507
rect 23676 16476 23857 16504
rect 23845 16473 23857 16476
rect 23891 16473 23903 16507
rect 24412 16504 24440 16612
rect 24489 16609 24501 16643
rect 24535 16609 24547 16643
rect 24489 16603 24547 16609
rect 24765 16643 24823 16649
rect 24765 16609 24777 16643
rect 24811 16640 24823 16643
rect 24854 16640 24860 16652
rect 24811 16612 24860 16640
rect 24811 16609 24823 16612
rect 24765 16603 24823 16609
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 27488 16612 27752 16640
rect 27488 16600 27494 16612
rect 26329 16575 26387 16581
rect 26329 16572 26341 16575
rect 26252 16544 26341 16572
rect 24412 16476 24900 16504
rect 23845 16467 23903 16473
rect 21818 16436 21824 16448
rect 19812 16408 21824 16436
rect 19705 16399 19763 16405
rect 21818 16396 21824 16408
rect 21876 16396 21882 16448
rect 23382 16396 23388 16448
rect 23440 16396 23446 16448
rect 23474 16396 23480 16448
rect 23532 16396 23538 16448
rect 23934 16396 23940 16448
rect 23992 16396 23998 16448
rect 24872 16436 24900 16476
rect 25406 16464 25412 16516
rect 25464 16464 25470 16516
rect 26142 16464 26148 16516
rect 26200 16464 26206 16516
rect 26160 16436 26188 16464
rect 26252 16448 26280 16544
rect 26329 16541 26341 16544
rect 26375 16541 26387 16575
rect 27724 16572 27752 16612
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27724 16544 28181 16572
rect 26329 16535 26387 16541
rect 28169 16541 28181 16544
rect 28215 16572 28227 16575
rect 28215 16544 30420 16572
rect 28215 16541 28227 16544
rect 28169 16535 28227 16541
rect 30392 16516 30420 16544
rect 26510 16464 26516 16516
rect 26568 16464 26574 16516
rect 27522 16464 27528 16516
rect 27580 16464 27586 16516
rect 28258 16464 28264 16516
rect 28316 16464 28322 16516
rect 28445 16507 28503 16513
rect 28445 16473 28457 16507
rect 28491 16473 28503 16507
rect 28445 16467 28503 16473
rect 24872 16408 26188 16436
rect 26234 16396 26240 16448
rect 26292 16396 26298 16448
rect 27540 16436 27568 16464
rect 28460 16436 28488 16467
rect 30374 16464 30380 16516
rect 30432 16464 30438 16516
rect 27540 16408 28488 16436
rect 1104 16346 30820 16368
rect 1104 16294 5324 16346
rect 5376 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 12752 16346
rect 12804 16294 12816 16346
rect 12868 16294 12880 16346
rect 12932 16294 12944 16346
rect 12996 16294 13008 16346
rect 13060 16294 20180 16346
rect 20232 16294 20244 16346
rect 20296 16294 20308 16346
rect 20360 16294 20372 16346
rect 20424 16294 20436 16346
rect 20488 16294 27608 16346
rect 27660 16294 27672 16346
rect 27724 16294 27736 16346
rect 27788 16294 27800 16346
rect 27852 16294 27864 16346
rect 27916 16294 30820 16346
rect 1104 16272 30820 16294
rect 3789 16235 3847 16241
rect 3789 16201 3801 16235
rect 3835 16232 3847 16235
rect 4154 16232 4160 16244
rect 3835 16204 4160 16232
rect 3835 16201 3847 16204
rect 3789 16195 3847 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6914 16232 6920 16244
rect 6227 16204 6920 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 7024 16204 8524 16232
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 7024 16164 7052 16204
rect 4028 16136 7052 16164
rect 4028 16124 4034 16136
rect 8294 16124 8300 16176
rect 8352 16124 8358 16176
rect 8496 16164 8524 16204
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 9398 16232 9404 16244
rect 8720 16204 9404 16232
rect 8720 16192 8726 16204
rect 9398 16192 9404 16204
rect 9456 16232 9462 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 9456 16204 13737 16232
rect 9456 16192 9462 16204
rect 13725 16201 13737 16204
rect 13771 16232 13783 16235
rect 18230 16232 18236 16244
rect 13771 16204 18236 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16201 18475 16235
rect 18417 16195 18475 16201
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 8496 16136 12265 16164
rect 12253 16133 12265 16136
rect 12299 16133 12311 16167
rect 12253 16127 12311 16133
rect 13538 16124 13544 16176
rect 13596 16164 13602 16176
rect 14366 16164 14372 16176
rect 13596 16136 14372 16164
rect 13596 16124 13602 16136
rect 1854 15988 1860 16040
rect 1912 16028 1918 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1912 16000 2053 16028
rect 1912 15988 1918 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2314 15988 2320 16040
rect 2372 15988 2378 16040
rect 3436 16028 3464 16082
rect 3602 16056 3608 16108
rect 3660 16096 3666 16108
rect 4062 16096 4068 16108
rect 3660 16068 4068 16096
rect 3660 16056 3666 16068
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4338 16096 4344 16108
rect 4172 16068 4344 16096
rect 4172 16037 4200 16068
rect 4338 16056 4344 16068
rect 4396 16056 4402 16108
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 5166 16056 5172 16108
rect 5224 16096 5230 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 5224 16068 5457 16096
rect 5224 16056 5230 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5718 16056 5724 16108
rect 5776 16056 5782 16108
rect 5994 16056 6000 16108
rect 6052 16056 6058 16108
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6457 16099 6515 16105
rect 6457 16096 6469 16099
rect 6227 16068 6469 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 6457 16065 6469 16068
rect 6503 16065 6515 16099
rect 6457 16059 6515 16065
rect 3973 16031 4031 16037
rect 3973 16028 3985 16031
rect 3436 16000 3985 16028
rect 3973 15997 3985 16000
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 15997 4215 16031
rect 4157 15991 4215 15997
rect 1670 15852 1676 15904
rect 1728 15892 1734 15904
rect 4172 15892 4200 15991
rect 5736 15960 5764 16056
rect 5905 16031 5963 16037
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6196 16028 6224 16059
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6730 16056 6736 16108
rect 6788 16056 6794 16108
rect 8110 16056 8116 16108
rect 8168 16056 8174 16108
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 5951 16000 6224 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6362 15988 6368 16040
rect 6420 16028 6426 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6420 16000 6653 16028
rect 6420 15988 6426 16000
rect 6641 15997 6653 16000
rect 6687 16028 6699 16031
rect 8220 16028 8248 16059
rect 8386 16056 8392 16108
rect 8444 16105 8450 16108
rect 8444 16099 8473 16105
rect 8461 16065 8473 16099
rect 8444 16059 8473 16065
rect 8444 16056 8450 16059
rect 8570 16056 8576 16108
rect 8628 16096 8634 16108
rect 8846 16096 8852 16108
rect 8628 16068 8852 16096
rect 8628 16056 8634 16068
rect 8846 16056 8852 16068
rect 8904 16056 8910 16108
rect 8938 16056 8944 16108
rect 8996 16056 9002 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11112 16068 11345 16096
rect 11112 16056 11118 16068
rect 11333 16065 11345 16068
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13906 16096 13912 16108
rect 13320 16068 13912 16096
rect 13320 16056 13326 16068
rect 13906 16056 13912 16068
rect 13964 16056 13970 16108
rect 14108 16105 14136 16136
rect 14366 16124 14372 16136
rect 14424 16124 14430 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15594 16136 16037 16164
rect 16025 16133 16037 16136
rect 16071 16133 16083 16167
rect 16025 16127 16083 16133
rect 16850 16124 16856 16176
rect 16908 16124 16914 16176
rect 17034 16124 17040 16176
rect 17092 16124 17098 16176
rect 17589 16167 17647 16173
rect 17589 16133 17601 16167
rect 17635 16164 17647 16167
rect 18138 16164 18144 16176
rect 17635 16136 18144 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 18432 16164 18460 16195
rect 18598 16192 18604 16244
rect 18656 16232 18662 16244
rect 19334 16232 19340 16244
rect 18656 16204 19340 16232
rect 18656 16192 18662 16204
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 23198 16192 23204 16244
rect 23256 16192 23262 16244
rect 24854 16192 24860 16244
rect 24912 16232 24918 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 24912 16204 25053 16232
rect 24912 16192 24918 16204
rect 25041 16201 25053 16204
rect 25087 16201 25099 16235
rect 25041 16195 25099 16201
rect 25130 16192 25136 16244
rect 25188 16192 25194 16244
rect 25406 16192 25412 16244
rect 25464 16192 25470 16244
rect 25593 16235 25651 16241
rect 25593 16201 25605 16235
rect 25639 16201 25651 16235
rect 25593 16195 25651 16201
rect 25700 16204 28212 16232
rect 18690 16164 18696 16176
rect 18432 16136 18696 16164
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 23937 16167 23995 16173
rect 20272 16136 23612 16164
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16868 16096 16896 16124
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16163 16068 16957 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 17052 16096 17080 16124
rect 17681 16099 17739 16105
rect 17681 16096 17693 16099
rect 17052 16068 17693 16096
rect 16945 16059 17003 16065
rect 17681 16065 17693 16068
rect 17727 16065 17739 16099
rect 17681 16059 17739 16065
rect 9398 16028 9404 16040
rect 6687 16000 8064 16028
rect 8220 16000 9404 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 7929 15963 7987 15969
rect 7929 15960 7941 15963
rect 5736 15932 7941 15960
rect 7929 15929 7941 15932
rect 7975 15929 7987 15963
rect 7929 15923 7987 15929
rect 1728 15864 4200 15892
rect 1728 15852 1734 15864
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5179 15895 5237 15901
rect 5179 15892 5191 15895
rect 5040 15864 5191 15892
rect 5040 15852 5046 15864
rect 5179 15861 5191 15864
rect 5225 15892 5237 15895
rect 5721 15895 5779 15901
rect 5721 15892 5733 15895
rect 5225 15864 5733 15892
rect 5225 15861 5237 15864
rect 5179 15855 5237 15861
rect 5721 15861 5733 15864
rect 5767 15892 5779 15895
rect 6178 15892 6184 15904
rect 5767 15864 6184 15892
rect 5767 15861 5779 15864
rect 5721 15855 5779 15861
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 6917 15895 6975 15901
rect 6917 15861 6929 15895
rect 6963 15892 6975 15895
rect 7466 15892 7472 15904
rect 6963 15864 7472 15892
rect 6963 15861 6975 15864
rect 6917 15855 6975 15861
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 8036 15892 8064 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11698 16028 11704 16040
rect 11195 16000 11704 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 13722 16028 13728 16040
rect 13596 16000 13728 16028
rect 13596 15988 13602 16000
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 16028 14427 16031
rect 14826 16028 14832 16040
rect 14415 16000 14832 16028
rect 14415 15997 14427 16000
rect 14369 15991 14427 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15856 15969 15884 16056
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15929 15899 15963
rect 17696 15960 17724 16059
rect 17770 16056 17776 16108
rect 17828 16056 17834 16108
rect 20272 16105 20300 16136
rect 23584 16108 23612 16136
rect 23937 16133 23949 16167
rect 23983 16164 23995 16167
rect 25148 16164 25176 16192
rect 25608 16164 25636 16195
rect 23983 16136 25176 16164
rect 25240 16136 25636 16164
rect 23983 16133 23995 16136
rect 23937 16127 23995 16133
rect 20257 16099 20315 16105
rect 18156 16068 18828 16096
rect 18156 16037 18184 16068
rect 18800 16040 18828 16068
rect 20257 16065 20269 16099
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20588 16068 20637 16096
rect 20588 16056 20594 16068
rect 20625 16065 20637 16068
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 23017 16099 23075 16105
rect 20947 16068 21956 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 18141 16031 18199 16037
rect 18141 15997 18153 16031
rect 18187 15997 18199 16031
rect 18141 15991 18199 15997
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 18598 16028 18604 16040
rect 18380 16000 18604 16028
rect 18380 15988 18386 16000
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 18782 15988 18788 16040
rect 18840 15988 18846 16040
rect 21928 15972 21956 16068
rect 23017 16065 23029 16099
rect 23063 16096 23075 16099
rect 23474 16096 23480 16108
rect 23063 16068 23480 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 23845 16099 23903 16105
rect 23845 16096 23857 16099
rect 23624 16068 23857 16096
rect 23624 16056 23630 16068
rect 23845 16065 23857 16068
rect 23891 16096 23903 16099
rect 25038 16096 25044 16108
rect 23891 16068 25044 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 25038 16056 25044 16068
rect 25096 16056 25102 16108
rect 25240 16105 25268 16136
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25314 16056 25320 16108
rect 25372 16056 25378 16108
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 25700 16028 25728 16204
rect 27430 16124 27436 16176
rect 27488 16124 27494 16176
rect 25961 16099 26019 16105
rect 25961 16065 25973 16099
rect 26007 16096 26019 16099
rect 26234 16096 26240 16108
rect 26007 16068 26240 16096
rect 26007 16065 26019 16068
rect 25961 16059 26019 16065
rect 26234 16056 26240 16068
rect 26292 16096 26298 16108
rect 26694 16096 26700 16108
rect 26292 16068 26700 16096
rect 26292 16056 26298 16068
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 26786 16056 26792 16108
rect 26844 16096 26850 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26844 16068 26985 16096
rect 26844 16056 26850 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27249 16099 27307 16105
rect 27249 16065 27261 16099
rect 27295 16096 27307 16099
rect 27448 16096 27476 16124
rect 27295 16068 27476 16096
rect 27295 16065 27307 16068
rect 27249 16059 27307 16065
rect 27614 16056 27620 16108
rect 27672 16056 27678 16108
rect 27982 16056 27988 16108
rect 28040 16056 28046 16108
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16096 28135 16099
rect 28184 16096 28212 16204
rect 28123 16068 28212 16096
rect 28261 16099 28319 16105
rect 28123 16065 28135 16068
rect 28077 16059 28135 16065
rect 28261 16065 28273 16099
rect 28307 16065 28319 16099
rect 28261 16059 28319 16065
rect 22152 16000 25728 16028
rect 22152 15988 22158 16000
rect 26050 15988 26056 16040
rect 26108 15988 26114 16040
rect 26142 15988 26148 16040
rect 26200 15988 26206 16040
rect 27632 16028 27660 16056
rect 28000 16028 28028 16056
rect 28276 16028 28304 16059
rect 27632 16000 27844 16028
rect 28000 16000 28304 16028
rect 18969 15963 19027 15969
rect 18969 15960 18981 15963
rect 17696 15932 18981 15960
rect 15841 15923 15899 15929
rect 18969 15929 18981 15932
rect 19015 15960 19027 15963
rect 19426 15960 19432 15972
rect 19015 15932 19432 15960
rect 19015 15929 19027 15932
rect 18969 15923 19027 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 21910 15920 21916 15972
rect 21968 15960 21974 15972
rect 21968 15932 26648 15960
rect 21968 15920 21974 15932
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8036 15864 8769 15892
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 8757 15855 8815 15861
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 14182 15892 14188 15904
rect 13136 15864 14188 15892
rect 13136 15852 13142 15864
rect 14182 15852 14188 15864
rect 14240 15892 14246 15904
rect 15654 15892 15660 15904
rect 14240 15864 15660 15892
rect 14240 15852 14246 15864
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 17034 15852 17040 15904
rect 17092 15852 17098 15904
rect 18598 15852 18604 15904
rect 18656 15901 18662 15904
rect 18656 15892 18667 15901
rect 18656 15864 18701 15892
rect 18656 15855 18667 15864
rect 18656 15852 18662 15855
rect 20162 15852 20168 15904
rect 20220 15852 20226 15904
rect 21634 15852 21640 15904
rect 21692 15852 21698 15904
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 26326 15892 26332 15904
rect 23348 15864 26332 15892
rect 23348 15852 23354 15864
rect 26326 15852 26332 15864
rect 26384 15852 26390 15904
rect 26620 15892 26648 15932
rect 27614 15920 27620 15972
rect 27672 15920 27678 15972
rect 27816 15960 27844 16000
rect 27985 15963 28043 15969
rect 27985 15960 27997 15963
rect 27816 15932 27997 15960
rect 27985 15929 27997 15932
rect 28031 15929 28043 15963
rect 27985 15923 28043 15929
rect 27632 15892 27660 15920
rect 26620 15864 27660 15892
rect 28166 15852 28172 15904
rect 28224 15852 28230 15904
rect 1104 15802 30820 15824
rect 1104 15750 4664 15802
rect 4716 15750 4728 15802
rect 4780 15750 4792 15802
rect 4844 15750 4856 15802
rect 4908 15750 4920 15802
rect 4972 15750 12092 15802
rect 12144 15750 12156 15802
rect 12208 15750 12220 15802
rect 12272 15750 12284 15802
rect 12336 15750 12348 15802
rect 12400 15750 19520 15802
rect 19572 15750 19584 15802
rect 19636 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 26948 15802
rect 27000 15750 27012 15802
rect 27064 15750 27076 15802
rect 27128 15750 27140 15802
rect 27192 15750 27204 15802
rect 27256 15750 30820 15802
rect 1104 15728 30820 15750
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2372 15660 2513 15688
rect 2372 15648 2378 15660
rect 2501 15657 2513 15660
rect 2547 15657 2559 15691
rect 2501 15651 2559 15657
rect 5905 15691 5963 15697
rect 5905 15657 5917 15691
rect 5951 15688 5963 15691
rect 5994 15688 6000 15700
rect 5951 15660 6000 15688
rect 5951 15657 5963 15660
rect 5905 15651 5963 15657
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6086 15648 6092 15700
rect 6144 15648 6150 15700
rect 8478 15648 8484 15700
rect 8536 15688 8542 15700
rect 8938 15688 8944 15700
rect 8536 15660 8944 15688
rect 8536 15648 8542 15660
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9398 15648 9404 15700
rect 9456 15648 9462 15700
rect 11238 15688 11244 15700
rect 10336 15660 11244 15688
rect 10336 15620 10364 15660
rect 4356 15592 7052 15620
rect 4356 15564 4384 15592
rect 7024 15564 7052 15592
rect 7208 15592 10364 15620
rect 7208 15564 7236 15592
rect 10888 15564 10916 15660
rect 11238 15648 11244 15660
rect 11296 15648 11302 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12161 15691 12219 15697
rect 12161 15688 12173 15691
rect 12032 15660 12173 15688
rect 12032 15648 12038 15660
rect 12161 15657 12173 15660
rect 12207 15657 12219 15691
rect 12161 15651 12219 15657
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13780 15660 13829 15688
rect 13780 15648 13786 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 14829 15691 14887 15697
rect 13817 15651 13875 15657
rect 14200 15660 14504 15688
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 13648 15620 13676 15648
rect 14200 15620 14228 15660
rect 13412 15592 14228 15620
rect 13412 15580 13418 15592
rect 4338 15512 4344 15564
rect 4396 15512 4402 15564
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 5224 15524 5825 15552
rect 5224 15512 5230 15524
rect 5813 15521 5825 15524
rect 5859 15552 5871 15555
rect 6086 15552 6092 15564
rect 5859 15524 6092 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 6086 15512 6092 15524
rect 6144 15512 6150 15564
rect 6178 15512 6184 15564
rect 6236 15552 6242 15564
rect 6822 15552 6828 15564
rect 6236 15524 6828 15552
rect 6236 15512 6242 15524
rect 2682 15444 2688 15496
rect 2740 15444 2746 15496
rect 6380 15493 6408 15524
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 7006 15512 7012 15564
rect 7064 15512 7070 15564
rect 7190 15512 7196 15564
rect 7248 15512 7254 15564
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 9171 15524 9674 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 6365 15487 6423 15493
rect 6365 15453 6377 15487
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 6546 15444 6552 15496
rect 6604 15444 6610 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9030 15484 9036 15496
rect 8987 15456 9036 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9214 15444 9220 15496
rect 9272 15444 9278 15496
rect 9646 15484 9674 15524
rect 10870 15512 10876 15564
rect 10928 15512 10934 15564
rect 11146 15512 11152 15564
rect 11204 15512 11210 15564
rect 13538 15552 13544 15564
rect 11900 15524 13544 15552
rect 9766 15484 9772 15496
rect 9646 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 9968 15456 10609 15484
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15385 5687 15419
rect 5629 15379 5687 15385
rect 6733 15419 6791 15425
rect 6733 15385 6745 15419
rect 6779 15385 6791 15419
rect 6733 15379 6791 15385
rect 5644 15348 5672 15379
rect 5718 15348 5724 15360
rect 5644 15320 5724 15348
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 6748 15348 6776 15379
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 9232 15416 9260 15444
rect 6880 15388 9260 15416
rect 6880 15376 6886 15388
rect 9968 15360 9996 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15484 11115 15487
rect 11164 15484 11192 15512
rect 11330 15484 11336 15496
rect 11103 15456 11336 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11900 15493 11928 15524
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 14200 15561 14228 15592
rect 13909 15555 13967 15561
rect 13909 15521 13921 15555
rect 13955 15521 13967 15555
rect 13909 15515 13967 15521
rect 14185 15555 14243 15561
rect 14185 15521 14197 15555
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 12437 15487 12495 15493
rect 12437 15453 12449 15487
rect 12483 15453 12495 15487
rect 12437 15447 12495 15453
rect 11517 15419 11575 15425
rect 11517 15385 11529 15419
rect 11563 15416 11575 15419
rect 11606 15416 11612 15428
rect 11563 15388 11612 15416
rect 11563 15385 11575 15388
rect 11517 15379 11575 15385
rect 11606 15376 11612 15388
rect 11664 15376 11670 15428
rect 11808 15416 11836 15447
rect 12452 15416 12480 15447
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13504 15456 13645 15484
rect 13504 15444 13510 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13722 15444 13728 15496
rect 13780 15444 13786 15496
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 13924 15484 13952 15515
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 14476 15552 14504 15660
rect 14829 15657 14841 15691
rect 14875 15688 14887 15691
rect 15010 15688 15016 15700
rect 14875 15660 15016 15688
rect 14875 15657 14887 15660
rect 14829 15651 14887 15657
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 17773 15691 17831 15697
rect 17773 15657 17785 15691
rect 17819 15688 17831 15691
rect 18138 15688 18144 15700
rect 17819 15660 18144 15688
rect 17819 15657 17831 15660
rect 17773 15651 17831 15657
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18874 15688 18880 15700
rect 18472 15660 18880 15688
rect 18472 15648 18478 15660
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 19502 15691 19560 15697
rect 19502 15688 19514 15691
rect 19352 15660 19514 15688
rect 17862 15580 17868 15632
rect 17920 15620 17926 15632
rect 18598 15620 18604 15632
rect 17920 15592 18604 15620
rect 17920 15580 17926 15592
rect 18598 15580 18604 15592
rect 18656 15580 18662 15632
rect 19061 15623 19119 15629
rect 19061 15589 19073 15623
rect 19107 15620 19119 15623
rect 19352 15620 19380 15660
rect 19502 15657 19514 15660
rect 19548 15657 19560 15691
rect 19502 15651 19560 15657
rect 20990 15648 20996 15700
rect 21048 15648 21054 15700
rect 21634 15648 21640 15700
rect 21692 15688 21698 15700
rect 22462 15688 22468 15700
rect 21692 15660 22468 15688
rect 21692 15648 21698 15660
rect 22462 15648 22468 15660
rect 22520 15688 22526 15700
rect 22557 15691 22615 15697
rect 22557 15688 22569 15691
rect 22520 15660 22569 15688
rect 22520 15648 22526 15660
rect 22557 15657 22569 15660
rect 22603 15657 22615 15691
rect 22557 15651 22615 15657
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23290 15688 23296 15700
rect 23063 15660 23296 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 23532 15660 23888 15688
rect 23532 15648 23538 15660
rect 23750 15620 23756 15632
rect 19107 15592 19380 15620
rect 21192 15592 23756 15620
rect 19107 15589 19119 15592
rect 19061 15583 19119 15589
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 14476 15524 15301 15552
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15473 15555 15531 15561
rect 15473 15521 15485 15555
rect 15519 15552 15531 15555
rect 15838 15552 15844 15564
rect 15519 15524 15844 15552
rect 15519 15521 15531 15524
rect 15473 15515 15531 15521
rect 15838 15512 15844 15524
rect 15896 15512 15902 15564
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 16040 15524 19257 15552
rect 13872 15456 13952 15484
rect 14384 15484 14412 15512
rect 16040 15493 16068 15524
rect 19245 15521 19257 15524
rect 19291 15552 19303 15555
rect 19978 15552 19984 15564
rect 19291 15524 19984 15552
rect 19291 15521 19303 15524
rect 19245 15515 19303 15521
rect 19978 15512 19984 15524
rect 20036 15552 20042 15564
rect 21192 15552 21220 15592
rect 23750 15580 23756 15592
rect 23808 15580 23814 15632
rect 23860 15620 23888 15660
rect 23934 15648 23940 15700
rect 23992 15688 23998 15700
rect 24121 15691 24179 15697
rect 24121 15688 24133 15691
rect 23992 15660 24133 15688
rect 23992 15648 23998 15660
rect 24121 15657 24133 15660
rect 24167 15657 24179 15691
rect 25225 15691 25283 15697
rect 25225 15688 25237 15691
rect 24121 15651 24179 15657
rect 24964 15660 25237 15688
rect 24964 15629 24992 15660
rect 25225 15657 25237 15660
rect 25271 15657 25283 15691
rect 25225 15651 25283 15657
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 26329 15691 26387 15697
rect 26329 15688 26341 15691
rect 26108 15660 26341 15688
rect 26108 15648 26114 15660
rect 26329 15657 26341 15660
rect 26375 15657 26387 15691
rect 26329 15651 26387 15657
rect 24949 15623 25007 15629
rect 24949 15620 24961 15623
rect 23860 15592 24961 15620
rect 24949 15589 24961 15592
rect 24995 15589 25007 15623
rect 24949 15583 25007 15589
rect 21634 15552 21640 15564
rect 20036 15524 21220 15552
rect 21560 15524 21640 15552
rect 20036 15512 20042 15524
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 14384 15456 16037 15484
rect 13872 15444 13878 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15484 18567 15487
rect 18690 15484 18696 15496
rect 18555 15456 18696 15484
rect 18555 15453 18567 15456
rect 18509 15447 18567 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 18923 15456 19288 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 14461 15419 14519 15425
rect 14461 15416 14473 15419
rect 11808 15388 12480 15416
rect 6696 15320 6776 15348
rect 6696 15308 6702 15320
rect 9950 15308 9956 15360
rect 10008 15308 10014 15360
rect 11149 15351 11207 15357
rect 11149 15317 11161 15351
rect 11195 15348 11207 15351
rect 11238 15348 11244 15360
rect 11195 15320 11244 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 12452 15348 12480 15388
rect 14292 15388 14473 15416
rect 14090 15348 14096 15360
rect 12452 15320 14096 15348
rect 14090 15308 14096 15320
rect 14148 15348 14154 15360
rect 14292 15348 14320 15388
rect 14461 15385 14473 15388
rect 14507 15385 14519 15419
rect 14461 15379 14519 15385
rect 15856 15388 16068 15416
rect 14148 15320 14320 15348
rect 14369 15351 14427 15357
rect 14148 15308 14154 15320
rect 14369 15317 14381 15351
rect 14415 15348 14427 15351
rect 14642 15348 14648 15360
rect 14415 15320 14648 15348
rect 14415 15317 14427 15320
rect 14369 15311 14427 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 15565 15351 15623 15357
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 15654 15348 15660 15360
rect 15611 15320 15660 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 15654 15308 15660 15320
rect 15712 15348 15718 15360
rect 15856 15348 15884 15388
rect 15712 15320 15884 15348
rect 15712 15308 15718 15320
rect 15930 15308 15936 15360
rect 15988 15308 15994 15360
rect 16040 15348 16068 15388
rect 16298 15376 16304 15428
rect 16356 15376 16362 15428
rect 17034 15376 17040 15428
rect 17092 15376 17098 15428
rect 17972 15348 18000 15444
rect 16040 15320 18000 15348
rect 19260 15348 19288 15456
rect 21358 15444 21364 15496
rect 21416 15444 21422 15496
rect 21560 15493 21588 15524
rect 21634 15512 21640 15524
rect 21692 15512 21698 15564
rect 22741 15555 22799 15561
rect 22741 15552 22753 15555
rect 22480 15524 22753 15552
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 22278 15444 22284 15496
rect 22336 15444 22342 15496
rect 22480 15493 22508 15524
rect 22741 15521 22753 15524
rect 22787 15552 22799 15555
rect 23290 15552 23296 15564
rect 22787 15524 23296 15552
rect 22787 15521 22799 15524
rect 22741 15515 22799 15521
rect 23290 15512 23296 15524
rect 23348 15512 23354 15564
rect 23845 15555 23903 15561
rect 23845 15521 23857 15555
rect 23891 15552 23903 15555
rect 24302 15552 24308 15564
rect 23891 15524 24308 15552
rect 23891 15521 23903 15524
rect 23845 15515 23903 15521
rect 24302 15512 24308 15524
rect 24360 15512 24366 15564
rect 26421 15555 26479 15561
rect 26421 15521 26433 15555
rect 26467 15552 26479 15555
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 26467 15524 27169 15552
rect 26467 15521 26479 15524
rect 26421 15515 26479 15521
rect 27157 15521 27169 15524
rect 27203 15521 27215 15555
rect 28166 15552 28172 15564
rect 27157 15515 27215 15521
rect 27356 15524 28172 15552
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 22830 15444 22836 15496
rect 22888 15444 22894 15496
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 23032 15456 23244 15484
rect 20162 15376 20168 15428
rect 20220 15376 20226 15428
rect 21008 15388 21864 15416
rect 21008 15360 21036 15388
rect 19702 15348 19708 15360
rect 19260 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 20990 15308 20996 15360
rect 21048 15308 21054 15360
rect 21174 15308 21180 15360
rect 21232 15348 21238 15360
rect 21453 15351 21511 15357
rect 21453 15348 21465 15351
rect 21232 15320 21465 15348
rect 21232 15308 21238 15320
rect 21453 15317 21465 15320
rect 21499 15317 21511 15351
rect 21836 15348 21864 15388
rect 21910 15376 21916 15428
rect 21968 15416 21974 15428
rect 22557 15419 22615 15425
rect 22557 15416 22569 15419
rect 21968 15388 22569 15416
rect 21968 15376 21974 15388
rect 22557 15385 22569 15388
rect 22603 15385 22615 15419
rect 23032 15416 23060 15456
rect 22557 15379 22615 15385
rect 22848 15388 23060 15416
rect 23109 15419 23167 15425
rect 22094 15348 22100 15360
rect 21836 15320 22100 15348
rect 21453 15311 21511 15317
rect 22094 15308 22100 15320
rect 22152 15308 22158 15360
rect 22465 15351 22523 15357
rect 22465 15317 22477 15351
rect 22511 15348 22523 15351
rect 22848 15348 22876 15388
rect 23109 15385 23121 15419
rect 23155 15385 23167 15419
rect 23216 15416 23244 15456
rect 23400 15456 23673 15484
rect 23309 15419 23367 15425
rect 23309 15416 23321 15419
rect 23216 15388 23321 15416
rect 23109 15379 23167 15385
rect 23309 15385 23321 15388
rect 23355 15385 23367 15419
rect 23309 15379 23367 15385
rect 22511 15320 22876 15348
rect 23124 15348 23152 15379
rect 23198 15348 23204 15360
rect 23124 15320 23204 15348
rect 22511 15317 22523 15320
rect 22465 15311 22523 15317
rect 23198 15308 23204 15320
rect 23256 15308 23262 15360
rect 23400 15348 23428 15456
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15484 23811 15487
rect 23799 15456 23888 15484
rect 23799 15453 23811 15456
rect 23753 15447 23811 15453
rect 23860 15428 23888 15456
rect 23934 15444 23940 15496
rect 23992 15444 23998 15496
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24946 15484 24952 15496
rect 24627 15456 24952 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24946 15444 24952 15456
rect 25004 15484 25010 15496
rect 25133 15487 25191 15493
rect 25133 15484 25145 15487
rect 25004 15456 25145 15484
rect 25004 15444 25010 15456
rect 25133 15453 25145 15456
rect 25179 15453 25191 15487
rect 25133 15447 25191 15453
rect 25958 15444 25964 15496
rect 26016 15484 26022 15496
rect 26145 15487 26203 15493
rect 26145 15484 26157 15487
rect 26016 15456 26157 15484
rect 26016 15444 26022 15456
rect 26145 15453 26157 15456
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 26234 15444 26240 15496
rect 26292 15444 26298 15496
rect 26326 15444 26332 15496
rect 26384 15444 26390 15496
rect 27356 15493 27384 15524
rect 28166 15512 28172 15524
rect 28224 15512 28230 15564
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 27522 15444 27528 15496
rect 27580 15444 27586 15496
rect 27617 15487 27675 15493
rect 27617 15453 27629 15487
rect 27663 15484 27675 15487
rect 28258 15484 28264 15496
rect 27663 15456 28264 15484
rect 27663 15453 27675 15456
rect 27617 15447 27675 15453
rect 23842 15376 23848 15428
rect 23900 15376 23906 15428
rect 26344 15416 26372 15444
rect 27632 15416 27660 15447
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 26344 15388 27660 15416
rect 23477 15351 23535 15357
rect 23477 15348 23489 15351
rect 23400 15320 23489 15348
rect 23477 15317 23489 15320
rect 23523 15317 23535 15351
rect 23477 15311 23535 15317
rect 25038 15308 25044 15360
rect 25096 15308 25102 15360
rect 25590 15308 25596 15360
rect 25648 15308 25654 15360
rect 1104 15258 30820 15280
rect 1104 15206 5324 15258
rect 5376 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 12752 15258
rect 12804 15206 12816 15258
rect 12868 15206 12880 15258
rect 12932 15206 12944 15258
rect 12996 15206 13008 15258
rect 13060 15206 20180 15258
rect 20232 15206 20244 15258
rect 20296 15206 20308 15258
rect 20360 15206 20372 15258
rect 20424 15206 20436 15258
rect 20488 15206 27608 15258
rect 27660 15206 27672 15258
rect 27724 15206 27736 15258
rect 27788 15206 27800 15258
rect 27852 15206 27864 15258
rect 27916 15206 30820 15258
rect 1104 15184 30820 15206
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 6730 15144 6736 15156
rect 6043 15116 6736 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 6932 15116 8432 15144
rect 3605 15079 3663 15085
rect 3605 15045 3617 15079
rect 3651 15045 3663 15079
rect 6546 15076 6552 15088
rect 3605 15039 3663 15045
rect 5920 15048 6552 15076
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 3620 15008 3648 15039
rect 5920 15017 5948 15048
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 5905 15011 5963 15017
rect 3620 14980 5856 15008
rect 3786 14900 3792 14952
rect 3844 14940 3850 14952
rect 4522 14940 4528 14952
rect 3844 14912 4528 14940
rect 3844 14900 3850 14912
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 5828 14940 5856 14980
rect 5905 14977 5917 15011
rect 5951 14977 5963 15011
rect 5905 14971 5963 14977
rect 6730 14940 6736 14952
rect 5828 14912 6736 14940
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 6932 14872 6960 15116
rect 7006 15036 7012 15088
rect 7064 15036 7070 15088
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 8202 15076 8208 15088
rect 7156 15048 8208 15076
rect 7156 15036 7162 15048
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 8404 15076 8432 15116
rect 8478 15104 8484 15156
rect 8536 15104 8542 15156
rect 10226 15144 10232 15156
rect 9416 15116 10232 15144
rect 9416 15076 9444 15116
rect 10226 15104 10232 15116
rect 10284 15144 10290 15156
rect 11054 15144 11060 15156
rect 10284 15116 11060 15144
rect 10284 15104 10290 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 13814 15144 13820 15156
rect 11992 15116 13820 15144
rect 9674 15076 9680 15088
rect 8404 15048 9444 15076
rect 9508 15048 9680 15076
rect 7024 15008 7052 15036
rect 9508 15017 9536 15048
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 11992 15085 12020 15116
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14921 15147 14979 15153
rect 14921 15113 14933 15147
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16298 15144 16304 15156
rect 16071 15116 16304 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15045 12035 15079
rect 11977 15039 12035 15045
rect 12066 15036 12072 15088
rect 12124 15036 12130 15088
rect 12207 15079 12265 15085
rect 12207 15045 12219 15079
rect 12253 15076 12265 15079
rect 13630 15076 13636 15088
rect 12253 15048 13636 15076
rect 12253 15045 12265 15048
rect 12207 15039 12265 15045
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 14936 15076 14964 15107
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 18046 15144 18052 15156
rect 18003 15116 18052 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 18414 15144 18420 15156
rect 18248 15116 18420 15144
rect 18248 15085 18276 15116
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 19702 15104 19708 15156
rect 19760 15104 19766 15156
rect 20073 15147 20131 15153
rect 20073 15113 20085 15147
rect 20119 15144 20131 15147
rect 20990 15144 20996 15156
rect 20119 15116 20996 15144
rect 20119 15113 20131 15116
rect 20073 15107 20131 15113
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21140 15116 21312 15144
rect 21140 15104 21146 15116
rect 17681 15079 17739 15085
rect 14936 15048 16068 15076
rect 7745 15011 7803 15017
rect 7745 15008 7757 15011
rect 7024 14980 7757 15008
rect 7745 14977 7757 14980
rect 7791 14977 7803 15011
rect 7745 14971 7803 14977
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11204 14980 11713 15008
rect 11204 14968 11210 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 11992 14980 13308 15008
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7469 14943 7527 14949
rect 7469 14940 7481 14943
rect 7248 14912 7481 14940
rect 7248 14900 7254 14912
rect 7469 14909 7481 14912
rect 7515 14909 7527 14943
rect 7469 14903 7527 14909
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9766 14940 9772 14952
rect 9723 14912 9772 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 9950 14900 9956 14952
rect 10008 14900 10014 14952
rect 10870 14900 10876 14952
rect 10928 14940 10934 14952
rect 11992 14940 12020 14980
rect 10928 14912 12020 14940
rect 12345 14943 12403 14949
rect 10928 14900 10934 14912
rect 12345 14909 12357 14943
rect 12391 14940 12403 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12391 14912 12449 14940
rect 12391 14909 12403 14912
rect 12345 14903 12403 14909
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 9968 14872 9996 14900
rect 3896 14844 6960 14872
rect 9692 14844 9996 14872
rect 3896 14816 3924 14844
rect 2958 14764 2964 14816
rect 3016 14804 3022 14816
rect 3145 14807 3203 14813
rect 3145 14804 3157 14807
rect 3016 14776 3157 14804
rect 3016 14764 3022 14776
rect 3145 14773 3157 14776
rect 3191 14773 3203 14807
rect 3145 14767 3203 14773
rect 3878 14764 3884 14816
rect 3936 14764 3942 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 9692 14804 9720 14844
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 11974 14872 11980 14884
rect 11848 14844 11980 14872
rect 11848 14832 11854 14844
rect 11974 14832 11980 14844
rect 12032 14872 12038 14884
rect 13004 14872 13032 14903
rect 12032 14844 13032 14872
rect 13280 14872 13308 14980
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14093 15011 14151 15017
rect 14093 15008 14105 15011
rect 14056 14980 14105 15008
rect 14056 14968 14062 14980
rect 14093 14977 14105 14980
rect 14139 15008 14151 15011
rect 14139 14980 14688 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 13354 14900 13360 14952
rect 13412 14900 13418 14952
rect 13446 14900 13452 14952
rect 13504 14900 13510 14952
rect 14660 14940 14688 14980
rect 14734 14968 14740 15020
rect 14792 14968 14798 15020
rect 15120 15017 15148 15048
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15841 15011 15899 15017
rect 15841 14977 15853 15011
rect 15887 15008 15899 15011
rect 15930 15008 15936 15020
rect 15887 14980 15936 15008
rect 15887 14977 15899 14980
rect 15841 14971 15899 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 16040 15008 16068 15048
rect 17681 15045 17693 15079
rect 17727 15076 17739 15079
rect 18233 15079 18291 15085
rect 18233 15076 18245 15079
rect 17727 15048 18245 15076
rect 17727 15045 17739 15048
rect 17681 15039 17739 15045
rect 18233 15045 18245 15048
rect 18279 15045 18291 15079
rect 18233 15039 18291 15045
rect 18340 15048 19288 15076
rect 18340 15008 18368 15048
rect 19260 15020 19288 15048
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 21284 15085 21312 15116
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 22646 15144 22652 15156
rect 21876 15116 22652 15144
rect 21876 15104 21882 15116
rect 22646 15104 22652 15116
rect 22704 15104 22710 15156
rect 25590 15104 25596 15156
rect 25648 15144 25654 15156
rect 25685 15147 25743 15153
rect 25685 15144 25697 15147
rect 25648 15116 25697 15144
rect 25648 15104 25654 15116
rect 25685 15113 25697 15116
rect 25731 15144 25743 15147
rect 25731 15116 26188 15144
rect 25731 15113 25743 15116
rect 25685 15107 25743 15113
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 19392 15048 19441 15076
rect 19392 15036 19398 15048
rect 19429 15045 19441 15048
rect 19475 15045 19487 15079
rect 19429 15039 19487 15045
rect 21269 15079 21327 15085
rect 21269 15045 21281 15079
rect 21315 15045 21327 15079
rect 21269 15039 21327 15045
rect 21407 15079 21465 15085
rect 21407 15045 21419 15079
rect 21453 15076 21465 15079
rect 21453 15048 22416 15076
rect 21453 15045 21465 15048
rect 21407 15039 21465 15045
rect 16040 14980 18368 15008
rect 18782 14968 18788 15020
rect 18840 14968 18846 15020
rect 19242 14968 19248 15020
rect 19300 14968 19306 15020
rect 20165 15011 20223 15017
rect 20165 14977 20177 15011
rect 20211 15008 20223 15011
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20211 14980 20913 15008
rect 20211 14977 20223 14980
rect 20165 14971 20223 14977
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21545 15011 21603 15017
rect 21223 14980 21312 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 18506 14940 18512 14952
rect 13832 14912 14596 14940
rect 14660 14912 18512 14940
rect 13832 14872 13860 14912
rect 13280 14844 13860 14872
rect 13909 14875 13967 14881
rect 12032 14832 12038 14844
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 14274 14872 14280 14884
rect 13955 14844 14280 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 14568 14872 14596 14912
rect 18506 14900 18512 14912
rect 18564 14940 18570 14952
rect 20257 14943 20315 14949
rect 20257 14940 20269 14943
rect 18564 14912 20269 14940
rect 18564 14900 18570 14912
rect 20257 14909 20269 14912
rect 20303 14940 20315 14943
rect 20806 14940 20812 14952
rect 20303 14912 20812 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 14568 14844 18981 14872
rect 18969 14841 18981 14844
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 4120 14776 9720 14804
rect 4120 14764 4126 14776
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 13814 14804 13820 14816
rect 13688 14776 13820 14804
rect 13688 14764 13694 14776
rect 13814 14764 13820 14776
rect 13872 14804 13878 14816
rect 14185 14807 14243 14813
rect 14185 14804 14197 14807
rect 13872 14776 14197 14804
rect 13872 14764 13878 14776
rect 14185 14773 14197 14776
rect 14231 14773 14243 14807
rect 14185 14767 14243 14773
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15378 14804 15384 14816
rect 15335 14776 15384 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15378 14764 15384 14776
rect 15436 14804 15442 14816
rect 15654 14804 15660 14816
rect 15436 14776 15660 14804
rect 15436 14764 15442 14776
rect 15654 14764 15660 14776
rect 15712 14804 15718 14816
rect 17218 14804 17224 14816
rect 15712 14776 17224 14804
rect 15712 14764 15718 14776
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 18509 14807 18567 14813
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 18690 14804 18696 14816
rect 18555 14776 18696 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 18984 14804 19012 14835
rect 19058 14832 19064 14884
rect 19116 14872 19122 14884
rect 19245 14875 19303 14881
rect 19245 14872 19257 14875
rect 19116 14844 19257 14872
rect 19116 14832 19122 14844
rect 19245 14841 19257 14844
rect 19291 14841 19303 14875
rect 21100 14872 21128 14971
rect 21174 14872 21180 14884
rect 21100 14844 21180 14872
rect 19245 14835 19303 14841
rect 21174 14832 21180 14844
rect 21232 14832 21238 14884
rect 21082 14804 21088 14816
rect 18984 14776 21088 14804
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 21284 14804 21312 14980
rect 21545 14977 21557 15011
rect 21591 15008 21603 15011
rect 21726 15008 21732 15020
rect 21591 14980 21732 15008
rect 21591 14977 21603 14980
rect 21545 14971 21603 14977
rect 21726 14968 21732 14980
rect 21784 14968 21790 15020
rect 21821 15011 21879 15017
rect 21821 14977 21833 15011
rect 21867 15008 21879 15011
rect 21910 15008 21916 15020
rect 21867 14980 21916 15008
rect 21867 14977 21879 14980
rect 21821 14971 21879 14977
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22281 15011 22339 15017
rect 22060 14980 22103 15008
rect 22060 14968 22066 14980
rect 22281 14977 22293 15011
rect 22327 14977 22339 15011
rect 22388 15008 22416 15048
rect 22462 15036 22468 15088
rect 22520 15036 22526 15088
rect 26160 15020 26188 15116
rect 26234 15104 26240 15156
rect 26292 15144 26298 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 26292 15116 26525 15144
rect 26292 15104 26298 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 26513 15107 26571 15113
rect 23750 15008 23756 15020
rect 22388 14980 23756 15008
rect 22281 14971 22339 14977
rect 21358 14900 21364 14952
rect 21416 14900 21422 14952
rect 21376 14872 21404 14900
rect 22189 14875 22247 14881
rect 22189 14872 22201 14875
rect 21376 14844 22201 14872
rect 22189 14841 22201 14844
rect 22235 14872 22247 14875
rect 22296 14872 22324 14971
rect 23750 14968 23756 14980
rect 23808 14968 23814 15020
rect 24302 14968 24308 15020
rect 24360 15008 24366 15020
rect 25593 15011 25651 15017
rect 25593 15008 25605 15011
rect 24360 14980 25605 15008
rect 24360 14968 24366 14980
rect 25593 14977 25605 14980
rect 25639 14977 25651 15011
rect 25593 14971 25651 14977
rect 22235 14844 22324 14872
rect 22235 14841 22247 14844
rect 22189 14835 22247 14841
rect 22278 14804 22284 14816
rect 21284 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14804 22342 14816
rect 22649 14807 22707 14813
rect 22649 14804 22661 14807
rect 22336 14776 22661 14804
rect 22336 14764 22342 14776
rect 22649 14773 22661 14776
rect 22695 14773 22707 14807
rect 25608 14804 25636 14971
rect 25866 14968 25872 15020
rect 25924 15008 25930 15020
rect 25924 14980 26004 15008
rect 25924 14968 25930 14980
rect 25976 14940 26004 14980
rect 26050 14968 26056 15020
rect 26108 14968 26114 15020
rect 26142 14968 26148 15020
rect 26200 14968 26206 15020
rect 26694 14968 26700 15020
rect 26752 15008 26758 15020
rect 27249 15011 27307 15017
rect 27249 15008 27261 15011
rect 26752 14980 27261 15008
rect 26752 14968 26758 14980
rect 27249 14977 27261 14980
rect 27295 15008 27307 15011
rect 27801 15011 27859 15017
rect 27801 15008 27813 15011
rect 27295 14980 27813 15008
rect 27295 14977 27307 14980
rect 27249 14971 27307 14977
rect 27801 14977 27813 14980
rect 27847 14977 27859 15011
rect 27801 14971 27859 14977
rect 26237 14943 26295 14949
rect 26237 14940 26249 14943
rect 25976 14912 26249 14940
rect 26237 14909 26249 14912
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14909 26387 14943
rect 26329 14903 26387 14909
rect 25869 14875 25927 14881
rect 25869 14841 25881 14875
rect 25915 14872 25927 14875
rect 25958 14872 25964 14884
rect 25915 14844 25964 14872
rect 25915 14841 25927 14844
rect 25869 14835 25927 14841
rect 25958 14832 25964 14844
rect 26016 14832 26022 14884
rect 26344 14804 26372 14903
rect 27522 14900 27528 14952
rect 27580 14940 27586 14952
rect 27580 14912 27660 14940
rect 27580 14900 27586 14912
rect 27632 14881 27660 14912
rect 27617 14875 27675 14881
rect 27617 14841 27629 14875
rect 27663 14872 27675 14875
rect 27663 14844 27936 14872
rect 27663 14841 27675 14844
rect 27617 14835 27675 14841
rect 25608 14776 26372 14804
rect 22649 14767 22707 14773
rect 27706 14764 27712 14816
rect 27764 14764 27770 14816
rect 27908 14813 27936 14844
rect 27893 14807 27951 14813
rect 27893 14773 27905 14807
rect 27939 14773 27951 14807
rect 27893 14767 27951 14773
rect 28258 14764 28264 14816
rect 28316 14764 28322 14816
rect 1104 14714 30820 14736
rect 1104 14662 4664 14714
rect 4716 14662 4728 14714
rect 4780 14662 4792 14714
rect 4844 14662 4856 14714
rect 4908 14662 4920 14714
rect 4972 14662 12092 14714
rect 12144 14662 12156 14714
rect 12208 14662 12220 14714
rect 12272 14662 12284 14714
rect 12336 14662 12348 14714
rect 12400 14662 19520 14714
rect 19572 14662 19584 14714
rect 19636 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 26948 14714
rect 27000 14662 27012 14714
rect 27064 14662 27076 14714
rect 27128 14662 27140 14714
rect 27192 14662 27204 14714
rect 27256 14662 30820 14714
rect 1104 14640 30820 14662
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 3605 14603 3663 14609
rect 3605 14600 3617 14603
rect 3568 14572 3617 14600
rect 3568 14560 3574 14572
rect 3605 14569 3617 14572
rect 3651 14569 3663 14603
rect 3605 14563 3663 14569
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 5718 14600 5724 14612
rect 4571 14572 5724 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6638 14560 6644 14612
rect 6696 14560 6702 14612
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 9674 14600 9680 14612
rect 6880 14572 9680 14600
rect 6880 14560 6886 14572
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 9766 14560 9772 14612
rect 9824 14560 9830 14612
rect 10768 14603 10826 14609
rect 10768 14569 10780 14603
rect 10814 14600 10826 14603
rect 11146 14600 11152 14612
rect 10814 14572 11152 14600
rect 10814 14569 10826 14572
rect 10768 14563 10826 14569
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 11940 14572 13001 14600
rect 11940 14560 11946 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 12989 14563 13047 14569
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14569 13415 14603
rect 16942 14600 16948 14612
rect 13357 14563 13415 14569
rect 16684 14572 16948 14600
rect 4982 14532 4988 14544
rect 4540 14504 4988 14532
rect 4540 14464 4568 14504
rect 4982 14492 4988 14504
rect 5040 14532 5046 14544
rect 6840 14532 6868 14560
rect 5040 14504 6868 14532
rect 6932 14504 10012 14532
rect 5040 14492 5046 14504
rect 6932 14464 6960 14504
rect 4448 14436 4568 14464
rect 4816 14436 6960 14464
rect 1854 14356 1860 14408
rect 1912 14356 1918 14408
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 4028 14368 4077 14396
rect 4028 14356 4034 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4338 14356 4344 14408
rect 4396 14396 4402 14408
rect 4448 14405 4476 14436
rect 4816 14405 4844 14436
rect 6288 14405 6316 14436
rect 7374 14424 7380 14476
rect 7432 14424 7438 14476
rect 7576 14436 9904 14464
rect 4433 14399 4491 14405
rect 4433 14396 4445 14399
rect 4396 14368 4445 14396
rect 4396 14356 4402 14368
rect 4433 14365 4445 14368
rect 4479 14365 4491 14399
rect 4433 14359 4491 14365
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14365 4859 14399
rect 4801 14359 4859 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5997 14399 6055 14405
rect 5997 14396 6009 14399
rect 5123 14368 6009 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5997 14365 6009 14368
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 6549 14399 6607 14405
rect 6549 14365 6561 14399
rect 6595 14396 6607 14399
rect 6822 14396 6828 14408
rect 6595 14368 6828 14396
rect 6595 14365 6607 14368
rect 6549 14359 6607 14365
rect 2130 14288 2136 14340
rect 2188 14288 2194 14340
rect 3142 14288 3148 14340
rect 3200 14288 3206 14340
rect 4522 14328 4528 14340
rect 4080 14300 4528 14328
rect 4080 14272 4108 14300
rect 4522 14288 4528 14300
rect 4580 14328 4586 14340
rect 4816 14328 4844 14359
rect 4580 14300 4844 14328
rect 4580 14288 4586 14300
rect 1670 14220 1676 14272
rect 1728 14260 1734 14272
rect 3878 14260 3884 14272
rect 1728 14232 3884 14260
rect 1728 14220 1734 14232
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4062 14220 4068 14272
rect 4120 14220 4126 14272
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 5092 14260 5120 14359
rect 6012 14328 6040 14359
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 6917 14399 6975 14405
rect 6917 14365 6929 14399
rect 6963 14396 6975 14399
rect 7098 14396 7104 14408
rect 6963 14368 7104 14396
rect 6963 14365 6975 14368
rect 6917 14359 6975 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7466 14356 7472 14408
rect 7524 14356 7530 14408
rect 7576 14328 7604 14436
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 8036 14368 8309 14396
rect 8036 14340 8064 14368
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 6012 14300 7604 14328
rect 7742 14288 7748 14340
rect 7800 14288 7806 14340
rect 8018 14288 8024 14340
rect 8076 14288 8082 14340
rect 8110 14288 8116 14340
rect 8168 14288 8174 14340
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 9324 14328 9352 14359
rect 9674 14356 9680 14408
rect 9732 14356 9738 14408
rect 9876 14328 9904 14436
rect 9984 14408 10012 14504
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13372 14532 13400 14563
rect 16684 14532 16712 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 20530 14600 20536 14612
rect 17276 14572 20536 14600
rect 17276 14560 17282 14572
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 21416 14572 21465 14600
rect 21416 14560 21422 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 22925 14603 22983 14609
rect 22925 14600 22937 14603
rect 21453 14563 21511 14569
rect 21560 14572 22416 14600
rect 11848 14504 16712 14532
rect 11848 14492 11854 14504
rect 11514 14464 11520 14476
rect 10336 14436 11520 14464
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10336 14405 10364 14436
rect 11514 14424 11520 14436
rect 11572 14464 11578 14476
rect 11572 14436 12020 14464
rect 11572 14424 11578 14436
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14365 10379 14399
rect 10321 14359 10379 14365
rect 10336 14328 10364 14359
rect 10502 14356 10508 14408
rect 10560 14356 10566 14408
rect 11992 14396 12020 14436
rect 12066 14424 12072 14476
rect 12124 14464 12130 14476
rect 17236 14473 17264 14560
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 21560 14532 21588 14572
rect 21821 14535 21879 14541
rect 21821 14532 21833 14535
rect 18840 14504 21588 14532
rect 21652 14504 21833 14532
rect 18840 14492 18846 14504
rect 12253 14467 12311 14473
rect 12253 14464 12265 14467
rect 12124 14436 12265 14464
rect 12124 14424 12130 14436
rect 12253 14433 12265 14436
rect 12299 14464 12311 14467
rect 17221 14467 17279 14473
rect 12299 14436 13492 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12529 14399 12587 14405
rect 12529 14396 12541 14399
rect 11992 14368 12541 14396
rect 12529 14365 12541 14368
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14396 12863 14399
rect 13170 14396 13176 14408
rect 12851 14368 13176 14396
rect 12851 14365 12863 14368
rect 12805 14359 12863 14365
rect 13170 14356 13176 14368
rect 13228 14356 13234 14408
rect 13464 14405 13492 14436
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 17221 14427 17279 14433
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14433 17463 14467
rect 17405 14427 17463 14433
rect 17972 14436 19196 14464
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13596 14368 13737 14396
rect 13596 14356 13602 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 14182 14356 14188 14408
rect 14240 14356 14246 14408
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16114 14396 16120 14408
rect 16071 14368 16120 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16868 14368 16957 14396
rect 8260 14300 9674 14328
rect 9876 14300 10364 14328
rect 8260 14288 8266 14300
rect 4212 14232 5120 14260
rect 4212 14220 4218 14232
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7926 14260 7932 14272
rect 6788 14232 7932 14260
rect 6788 14220 6794 14232
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 9646 14260 9674 14300
rect 11238 14288 11244 14340
rect 11296 14288 11302 14340
rect 14369 14331 14427 14337
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 16574 14328 16580 14340
rect 14415 14300 16580 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 16574 14288 16580 14300
rect 16632 14288 16638 14340
rect 16868 14272 16896 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 17420 14396 17448 14427
rect 17770 14396 17776 14408
rect 17420 14368 17776 14396
rect 16945 14359 17003 14365
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 17862 14356 17868 14408
rect 17920 14396 17926 14408
rect 17972 14405 18000 14436
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 17920 14368 17969 14396
rect 17920 14356 17926 14368
rect 17957 14365 17969 14368
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14365 18199 14399
rect 18141 14359 18199 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 18463 14368 18828 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 17678 14288 17684 14340
rect 17736 14288 17742 14340
rect 18156 14272 18184 14359
rect 18800 14337 18828 14368
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 19061 14399 19119 14405
rect 19061 14396 19073 14399
rect 19024 14368 19073 14396
rect 19024 14356 19030 14368
rect 19061 14365 19073 14368
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19168 14340 19196 14436
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19300 14436 19993 14464
rect 19300 14424 19306 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19576 14368 19717 14396
rect 19576 14356 19582 14368
rect 19705 14365 19717 14368
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14396 19855 14399
rect 20070 14396 20076 14408
rect 19843 14368 20076 14396
rect 19843 14365 19855 14368
rect 19797 14359 19855 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 18785 14331 18843 14337
rect 18785 14297 18797 14331
rect 18831 14328 18843 14331
rect 18874 14328 18880 14340
rect 18831 14300 18880 14328
rect 18831 14297 18843 14300
rect 18785 14291 18843 14297
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 21284 14337 21312 14504
rect 21652 14396 21680 14504
rect 21821 14501 21833 14504
rect 21867 14501 21879 14535
rect 21821 14495 21879 14501
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22152 14436 22293 14464
rect 22152 14424 22158 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22388 14464 22416 14572
rect 22572 14572 22937 14600
rect 22462 14492 22468 14544
rect 22520 14532 22526 14544
rect 22572 14541 22600 14572
rect 22925 14569 22937 14572
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 23106 14560 23112 14612
rect 23164 14560 23170 14612
rect 23658 14560 23664 14612
rect 23716 14560 23722 14612
rect 23934 14560 23940 14612
rect 23992 14560 23998 14612
rect 24302 14560 24308 14612
rect 24360 14600 24366 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 24360 14572 24409 14600
rect 24360 14560 24366 14572
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 24946 14600 24952 14612
rect 24397 14563 24455 14569
rect 24504 14572 24952 14600
rect 22557 14535 22615 14541
rect 22557 14532 22569 14535
rect 22520 14504 22569 14532
rect 22520 14492 22526 14504
rect 22557 14501 22569 14504
rect 22603 14501 22615 14535
rect 23124 14532 23152 14560
rect 22557 14495 22615 14501
rect 22664 14504 23152 14532
rect 23477 14535 23535 14541
rect 22664 14464 22692 14504
rect 23477 14501 23489 14535
rect 23523 14532 23535 14535
rect 23952 14532 23980 14560
rect 23523 14504 23980 14532
rect 23523 14501 23535 14504
rect 23477 14495 23535 14501
rect 24504 14464 24532 14572
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 25038 14560 25044 14612
rect 25096 14600 25102 14612
rect 26053 14603 26111 14609
rect 26053 14600 26065 14603
rect 25096 14572 26065 14600
rect 25096 14560 25102 14572
rect 22388 14436 22692 14464
rect 23952 14436 24532 14464
rect 22281 14427 22339 14433
rect 21500 14371 21680 14396
rect 21499 14368 21680 14371
rect 21729 14399 21787 14405
rect 21499 14365 21557 14368
rect 19429 14331 19487 14337
rect 19429 14328 19441 14331
rect 19208 14300 19441 14328
rect 19208 14288 19214 14300
rect 19429 14297 19441 14300
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 21269 14331 21327 14337
rect 21269 14297 21281 14331
rect 21315 14297 21327 14331
rect 21499 14331 21511 14365
rect 21545 14331 21557 14365
rect 21729 14365 21741 14399
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21499 14325 21557 14331
rect 21744 14328 21772 14359
rect 21910 14356 21916 14408
rect 21968 14356 21974 14408
rect 22296 14396 22324 14427
rect 23952 14405 23980 14436
rect 25148 14415 25176 14572
rect 26053 14569 26065 14572
rect 26099 14569 26111 14603
rect 26053 14563 26111 14569
rect 27433 14603 27491 14609
rect 27433 14569 27445 14603
rect 27479 14569 27491 14603
rect 27433 14563 27491 14569
rect 25777 14535 25835 14541
rect 25777 14501 25789 14535
rect 25823 14501 25835 14535
rect 25777 14495 25835 14501
rect 25792 14464 25820 14495
rect 25866 14492 25872 14544
rect 25924 14532 25930 14544
rect 27448 14532 27476 14563
rect 27706 14560 27712 14612
rect 27764 14560 27770 14612
rect 28258 14560 28264 14612
rect 28316 14560 28322 14612
rect 25924 14504 27476 14532
rect 25924 14492 25930 14504
rect 27157 14467 27215 14473
rect 27157 14464 27169 14467
rect 25792 14436 27169 14464
rect 27157 14433 27169 14436
rect 27203 14433 27215 14467
rect 27157 14427 27215 14433
rect 27249 14467 27307 14473
rect 27249 14433 27261 14467
rect 27295 14464 27307 14467
rect 27724 14464 27752 14560
rect 27295 14436 27752 14464
rect 27295 14433 27307 14436
rect 27249 14427 27307 14433
rect 25133 14409 25191 14415
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22296 14368 22845 14396
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 23937 14399 23995 14405
rect 23937 14365 23949 14399
rect 23983 14365 23995 14399
rect 23937 14359 23995 14365
rect 24026 14356 24032 14408
rect 24084 14396 24090 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24084 14368 24593 14396
rect 24084 14356 24090 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24762 14356 24768 14408
rect 24820 14356 24826 14408
rect 24922 14399 24980 14405
rect 24922 14365 24934 14399
rect 24968 14396 24980 14399
rect 24968 14365 24992 14396
rect 24922 14359 24992 14365
rect 22002 14328 22008 14340
rect 21744 14300 22008 14328
rect 21269 14291 21327 14297
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 22278 14288 22284 14340
rect 22336 14328 22342 14340
rect 23842 14328 23848 14340
rect 22336 14300 23848 14328
rect 22336 14288 22342 14300
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 24673 14331 24731 14337
rect 24673 14297 24685 14331
rect 24719 14328 24731 14331
rect 24719 14300 24900 14328
rect 24719 14297 24731 14300
rect 24673 14291 24731 14297
rect 24872 14272 24900 14300
rect 24964 14272 24992 14359
rect 25038 14356 25044 14408
rect 25096 14356 25102 14408
rect 25133 14375 25145 14409
rect 25179 14375 25191 14409
rect 25133 14369 25191 14375
rect 25222 14356 25228 14408
rect 25280 14356 25286 14408
rect 25314 14356 25320 14408
rect 25372 14396 25378 14408
rect 25372 14368 25452 14396
rect 25372 14356 25378 14368
rect 25424 14337 25452 14368
rect 25590 14356 25596 14408
rect 25648 14356 25654 14408
rect 26142 14356 26148 14408
rect 26200 14396 26206 14408
rect 26329 14399 26387 14405
rect 26329 14396 26341 14399
rect 26200 14368 26341 14396
rect 26200 14356 26206 14368
rect 26329 14365 26341 14368
rect 26375 14396 26387 14399
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26375 14368 26985 14396
rect 26375 14365 26387 14368
rect 26329 14359 26387 14365
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 27065 14399 27123 14405
rect 27065 14365 27077 14399
rect 27111 14396 27123 14399
rect 27893 14399 27951 14405
rect 27893 14396 27905 14399
rect 27111 14368 27905 14396
rect 27111 14365 27123 14368
rect 27065 14359 27123 14365
rect 27893 14365 27905 14368
rect 27939 14396 27951 14399
rect 28276 14396 28304 14560
rect 27939 14368 28304 14396
rect 27939 14365 27951 14368
rect 27893 14359 27951 14365
rect 25409 14331 25467 14337
rect 25409 14297 25421 14331
rect 25455 14297 25467 14331
rect 25409 14291 25467 14297
rect 25498 14288 25504 14340
rect 25556 14288 25562 14340
rect 13262 14260 13268 14272
rect 9646 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14260 13326 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13320 14232 13645 14260
rect 13320 14220 13326 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14642 14220 14648 14272
rect 14700 14260 14706 14272
rect 16206 14260 16212 14272
rect 14700 14232 16212 14260
rect 14700 14220 14706 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16850 14220 16856 14272
rect 16908 14220 16914 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 19242 14260 19248 14272
rect 18196 14232 19248 14260
rect 18196 14220 18202 14232
rect 19242 14220 19248 14232
rect 19300 14220 19306 14272
rect 21637 14263 21695 14269
rect 21637 14229 21649 14263
rect 21683 14260 21695 14263
rect 22186 14260 22192 14272
rect 21683 14232 22192 14260
rect 21683 14229 21695 14232
rect 21637 14223 21695 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22738 14220 22744 14272
rect 22796 14220 22802 14272
rect 23198 14220 23204 14272
rect 23256 14260 23262 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 23256 14232 23305 14260
rect 23256 14220 23262 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 25869 14263 25927 14269
rect 25869 14260 25881 14263
rect 25004 14232 25881 14260
rect 25004 14220 25010 14232
rect 25869 14229 25881 14232
rect 25915 14260 25927 14263
rect 26142 14260 26148 14272
rect 25915 14232 26148 14260
rect 25915 14229 25927 14232
rect 25869 14223 25927 14229
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26326 14220 26332 14272
rect 26384 14260 26390 14272
rect 26789 14263 26847 14269
rect 26789 14260 26801 14263
rect 26384 14232 26801 14260
rect 26384 14220 26390 14232
rect 26789 14229 26801 14232
rect 26835 14229 26847 14263
rect 26789 14223 26847 14229
rect 1104 14170 30820 14192
rect 1104 14118 5324 14170
rect 5376 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 12752 14170
rect 12804 14118 12816 14170
rect 12868 14118 12880 14170
rect 12932 14118 12944 14170
rect 12996 14118 13008 14170
rect 13060 14118 20180 14170
rect 20232 14118 20244 14170
rect 20296 14118 20308 14170
rect 20360 14118 20372 14170
rect 20424 14118 20436 14170
rect 20488 14118 27608 14170
rect 27660 14118 27672 14170
rect 27724 14118 27736 14170
rect 27788 14118 27800 14170
rect 27852 14118 27864 14170
rect 27916 14118 30820 14170
rect 1104 14096 30820 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 2409 14059 2467 14065
rect 2409 14056 2421 14059
rect 2188 14028 2421 14056
rect 2188 14016 2194 14028
rect 2409 14025 2421 14028
rect 2455 14025 2467 14059
rect 2958 14056 2964 14068
rect 2409 14019 2467 14025
rect 2746 14028 2964 14056
rect 934 13880 940 13932
rect 992 13920 998 13932
rect 1397 13923 1455 13929
rect 1397 13920 1409 13923
rect 992 13892 1409 13920
rect 992 13880 998 13892
rect 1397 13889 1409 13892
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 1670 13880 1676 13932
rect 1728 13880 1734 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2746 13920 2774 14028
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 3053 14059 3111 14065
rect 3053 14025 3065 14059
rect 3099 14056 3111 14059
rect 3142 14056 3148 14068
rect 3099 14028 3148 14056
rect 3099 14025 3111 14028
rect 3053 14019 3111 14025
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3510 14016 3516 14068
rect 3568 14016 3574 14068
rect 4338 14056 4344 14068
rect 3804 14028 4344 14056
rect 2639 13892 2774 13920
rect 3145 13923 3203 13929
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3191 13892 3464 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3252 13716 3280 13815
rect 3436 13784 3464 13892
rect 3528 13852 3556 14016
rect 3804 13929 3832 14028
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 7745 14059 7803 14065
rect 7340 14028 7604 14056
rect 7340 14016 7346 14028
rect 3896 13960 6592 13988
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3896 13852 3924 13960
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13920 4031 13923
rect 4062 13920 4068 13932
rect 4019 13892 4068 13920
rect 4019 13889 4031 13892
rect 3973 13883 4031 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4356 13929 4384 13960
rect 6564 13932 6592 13960
rect 7466 13948 7472 14000
rect 7524 13948 7530 14000
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 3528 13824 3924 13852
rect 4525 13855 4583 13861
rect 4525 13836 4537 13855
rect 4448 13821 4537 13836
rect 4571 13821 4583 13855
rect 4448 13815 4583 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 4448 13808 4568 13815
rect 3602 13784 3608 13796
rect 3436 13756 3608 13784
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 3697 13787 3755 13793
rect 3697 13753 3709 13787
rect 3743 13784 3755 13787
rect 4448 13784 4476 13808
rect 4816 13784 4844 13815
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 7484 13852 7512 13948
rect 7576 13929 7604 14028
rect 7745 14025 7757 14059
rect 7791 14056 7803 14059
rect 8110 14056 8116 14068
rect 7791 14028 8116 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 7852 13929 7880 14028
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 8297 14059 8355 14065
rect 8297 14025 8309 14059
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8312 13988 8340 14019
rect 8478 14016 8484 14068
rect 8536 14016 8542 14068
rect 9122 14016 9128 14068
rect 9180 14016 9186 14068
rect 9398 14016 9404 14068
rect 9456 14016 9462 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 11057 14059 11115 14065
rect 9732 14028 11008 14056
rect 9732 14016 9738 14028
rect 7984 13960 8340 13988
rect 7984 13948 7990 13960
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13889 7619 13923
rect 7561 13883 7619 13889
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 7760 13852 7788 13883
rect 8018 13880 8024 13932
rect 8076 13880 8082 13932
rect 8496 13929 8524 14016
rect 9140 13988 9168 14016
rect 8772 13960 9168 13988
rect 9217 13991 9275 13997
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 7484 13824 7788 13852
rect 7926 13812 7932 13864
rect 7984 13812 7990 13864
rect 5534 13784 5540 13796
rect 3743 13756 4476 13784
rect 4724 13756 5540 13784
rect 3743 13753 3755 13756
rect 3697 13747 3755 13753
rect 3970 13716 3976 13728
rect 3252 13688 3976 13716
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 4724 13716 4752 13756
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 6917 13787 6975 13793
rect 6917 13753 6929 13787
rect 6963 13784 6975 13787
rect 8036 13784 8064 13880
rect 8110 13812 8116 13864
rect 8168 13852 8174 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 8168 13824 8585 13852
rect 8168 13812 8174 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 8662 13812 8668 13864
rect 8720 13812 8726 13864
rect 8772 13861 8800 13960
rect 9217 13957 9229 13991
rect 9263 13988 9275 13991
rect 9553 13991 9611 13997
rect 9553 13988 9565 13991
rect 9263 13960 9565 13988
rect 9263 13957 9275 13960
rect 9217 13951 9275 13957
rect 9553 13957 9565 13960
rect 9599 13957 9611 13991
rect 9553 13951 9611 13957
rect 9769 13991 9827 13997
rect 9769 13957 9781 13991
rect 9815 13988 9827 13991
rect 10134 13988 10140 14000
rect 9815 13960 10140 13988
rect 9815 13957 9827 13960
rect 9769 13951 9827 13957
rect 10134 13948 10140 13960
rect 10192 13988 10198 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10192 13960 10793 13988
rect 10192 13948 10198 13960
rect 10781 13957 10793 13960
rect 10827 13988 10839 13991
rect 10870 13988 10876 14000
rect 10827 13960 10876 13988
rect 10827 13957 10839 13960
rect 10781 13951 10839 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 10980 13988 11008 14028
rect 11057 14025 11069 14059
rect 11103 14056 11115 14059
rect 11146 14056 11152 14068
rect 11103 14028 11152 14056
rect 11103 14025 11115 14028
rect 11057 14019 11115 14025
rect 11146 14016 11152 14028
rect 11204 14056 11210 14068
rect 11790 14056 11796 14068
rect 11204 14028 11796 14056
rect 11204 14016 11210 14028
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 14550 14056 14556 14068
rect 14016 14028 14556 14056
rect 11606 13988 11612 14000
rect 10980 13960 11612 13988
rect 11606 13948 11612 13960
rect 11664 13948 11670 14000
rect 11698 13948 11704 14000
rect 11756 13988 11762 14000
rect 13173 13991 13231 13997
rect 13173 13988 13185 13991
rect 11756 13960 13185 13988
rect 11756 13948 11762 13960
rect 13173 13957 13185 13960
rect 13219 13957 13231 13991
rect 13173 13951 13231 13957
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9309 13923 9367 13929
rect 9171 13892 9260 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9232 13864 9260 13892
rect 9309 13889 9321 13923
rect 9355 13920 9367 13923
rect 9355 13892 9628 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 9600 13864 9628 13892
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9732 13892 9873 13920
rect 9732 13880 9738 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 13078 13920 13084 13932
rect 12299 13892 13084 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 9214 13812 9220 13864
rect 9272 13812 9278 13864
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 10060 13852 10088 13883
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 13906 13920 13912 13932
rect 13495 13892 13912 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14016 13929 14044 14028
rect 14550 14016 14556 14028
rect 14608 14056 14614 14068
rect 17678 14056 17684 14068
rect 14608 14028 16712 14056
rect 14608 14016 14614 14028
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16114 13920 16120 13932
rect 15427 13892 16120 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16684 13929 16712 14028
rect 16868 14028 17684 14056
rect 16868 13997 16896 14028
rect 17678 14016 17684 14028
rect 17736 14016 17742 14068
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 19058 14056 19064 14068
rect 17828 14028 19064 14056
rect 17828 14016 17834 14028
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13957 16911 13991
rect 16853 13951 16911 13957
rect 18616 13929 18644 14028
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 22738 14016 22744 14068
rect 22796 14016 22802 14068
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14056 23259 14059
rect 23658 14056 23664 14068
rect 23247 14028 23664 14056
rect 23247 14025 23259 14028
rect 23201 14019 23259 14025
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25498 14056 25504 14068
rect 24912 14028 25504 14056
rect 24912 14016 24918 14028
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 21450 13988 21456 14000
rect 18892 13960 19564 13988
rect 18892 13932 18920 13960
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18874 13880 18880 13932
rect 18932 13880 18938 13932
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19242 13880 19248 13932
rect 19300 13880 19306 13932
rect 19536 13929 19564 13960
rect 19812 13960 21456 13988
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 19812 13929 19840 13960
rect 21450 13948 21456 13960
rect 21508 13948 21514 14000
rect 22756 13988 22784 14016
rect 24673 13991 24731 13997
rect 24673 13988 24685 13991
rect 22756 13960 24685 13988
rect 23297 13957 23355 13960
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19668 13892 19809 13920
rect 19668 13880 19674 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20990 13920 20996 13932
rect 20119 13892 20996 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21082 13880 21088 13932
rect 21140 13920 21146 13932
rect 22094 13920 22100 13932
rect 21140 13892 22100 13920
rect 21140 13880 21146 13892
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13889 23075 13923
rect 23198 13920 23204 13932
rect 23017 13883 23075 13889
rect 23124 13892 23204 13920
rect 9640 13824 10088 13852
rect 9640 13812 9646 13824
rect 11974 13812 11980 13864
rect 12032 13812 12038 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 13596 13824 14044 13852
rect 13596 13812 13602 13824
rect 6963 13756 8064 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 9950 13744 9956 13796
rect 10008 13784 10014 13796
rect 11992 13784 12020 13812
rect 10008 13756 12020 13784
rect 10008 13744 10014 13756
rect 4120 13688 4752 13716
rect 4120 13676 4126 13688
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 9548 13688 9597 13716
rect 9548 13676 9554 13688
rect 9585 13685 9597 13688
rect 9631 13716 9643 13719
rect 10229 13719 10287 13725
rect 10229 13716 10241 13719
rect 9631 13688 10241 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 10229 13685 10241 13688
rect 10275 13685 10287 13719
rect 14016 13716 14044 13824
rect 14090 13812 14096 13864
rect 14148 13852 14154 13864
rect 14642 13852 14648 13864
rect 14148 13824 14648 13852
rect 14148 13812 14154 13824
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15654 13812 15660 13864
rect 15712 13812 15718 13864
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 16908 13824 17141 13852
rect 16908 13812 16914 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 19426 13812 19432 13864
rect 19484 13812 19490 13864
rect 14369 13787 14427 13793
rect 14369 13753 14381 13787
rect 14415 13784 14427 13787
rect 20809 13787 20867 13793
rect 14415 13756 15148 13784
rect 14415 13753 14427 13756
rect 14369 13747 14427 13753
rect 14645 13719 14703 13725
rect 14645 13716 14657 13719
rect 14016 13688 14657 13716
rect 10229 13679 10287 13685
rect 14645 13685 14657 13688
rect 14691 13685 14703 13719
rect 15120 13716 15148 13756
rect 20809 13753 20821 13787
rect 20855 13784 20867 13787
rect 22002 13784 22008 13796
rect 20855 13756 22008 13784
rect 20855 13753 20867 13756
rect 20809 13747 20867 13753
rect 22002 13744 22008 13756
rect 22060 13784 22066 13796
rect 22830 13784 22836 13796
rect 22060 13756 22836 13784
rect 22060 13744 22066 13756
rect 22830 13744 22836 13756
rect 22888 13744 22894 13796
rect 15286 13716 15292 13728
rect 15120 13688 15292 13716
rect 14645 13679 14703 13685
rect 15286 13676 15292 13688
rect 15344 13676 15350 13728
rect 22738 13676 22744 13728
rect 22796 13716 22802 13728
rect 22940 13716 22968 13883
rect 23032 13784 23060 13883
rect 23124 13861 23152 13892
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23297 13923 23309 13957
rect 23343 13923 23355 13957
rect 24673 13957 24685 13960
rect 24719 13988 24731 13991
rect 25038 13988 25044 14000
rect 24719 13960 25044 13988
rect 24719 13957 24731 13960
rect 24673 13951 24731 13957
rect 25038 13948 25044 13960
rect 25096 13948 25102 14000
rect 23297 13917 23355 13923
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24762 13920 24768 13932
rect 23532 13892 24768 13920
rect 23532 13880 23538 13892
rect 24762 13880 24768 13892
rect 24820 13920 24826 13932
rect 25314 13920 25320 13932
rect 24820 13892 25320 13920
rect 24820 13880 24826 13892
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23842 13784 23848 13796
rect 23032 13756 23848 13784
rect 23842 13744 23848 13756
rect 23900 13744 23906 13796
rect 24026 13744 24032 13796
rect 24084 13744 24090 13796
rect 24964 13793 24992 13892
rect 25314 13880 25320 13892
rect 25372 13880 25378 13932
rect 25884 13920 25912 14016
rect 26145 13923 26203 13929
rect 26145 13920 26157 13923
rect 25884 13892 26157 13920
rect 26145 13889 26157 13892
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 26234 13812 26240 13864
rect 26292 13812 26298 13864
rect 24949 13787 25007 13793
rect 24949 13753 24961 13787
rect 24995 13753 25007 13787
rect 24949 13747 25007 13753
rect 24044 13716 24072 13744
rect 22796 13688 24072 13716
rect 22796 13676 22802 13688
rect 25130 13676 25136 13728
rect 25188 13676 25194 13728
rect 26142 13676 26148 13728
rect 26200 13676 26206 13728
rect 26510 13676 26516 13728
rect 26568 13676 26574 13728
rect 1104 13626 30820 13648
rect 1104 13574 4664 13626
rect 4716 13574 4728 13626
rect 4780 13574 4792 13626
rect 4844 13574 4856 13626
rect 4908 13574 4920 13626
rect 4972 13574 12092 13626
rect 12144 13574 12156 13626
rect 12208 13574 12220 13626
rect 12272 13574 12284 13626
rect 12336 13574 12348 13626
rect 12400 13574 19520 13626
rect 19572 13574 19584 13626
rect 19636 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 26948 13626
rect 27000 13574 27012 13626
rect 27064 13574 27076 13626
rect 27128 13574 27140 13626
rect 27192 13574 27204 13626
rect 27256 13574 30820 13626
rect 1104 13552 30820 13574
rect 6638 13512 6644 13524
rect 4632 13484 6644 13512
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 4632 13317 4660 13484
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8846 13512 8852 13524
rect 8352 13484 8852 13512
rect 8352 13472 8358 13484
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 10229 13515 10287 13521
rect 10229 13512 10241 13515
rect 8904 13484 10241 13512
rect 8904 13472 8910 13484
rect 10229 13481 10241 13484
rect 10275 13481 10287 13515
rect 10229 13475 10287 13481
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 16632 13484 17693 13512
rect 16632 13472 16638 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 17681 13475 17739 13481
rect 23474 13472 23480 13524
rect 23532 13472 23538 13524
rect 23750 13472 23756 13524
rect 23808 13512 23814 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 23808 13484 24593 13512
rect 23808 13472 23814 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 26234 13512 26240 13524
rect 25547 13484 26240 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 26789 13515 26847 13521
rect 26789 13481 26801 13515
rect 26835 13512 26847 13515
rect 28350 13512 28356 13524
rect 26835 13484 28356 13512
rect 26835 13481 26847 13484
rect 26789 13475 26847 13481
rect 28350 13472 28356 13484
rect 28408 13472 28414 13524
rect 6656 13444 6684 13472
rect 9398 13444 9404 13456
rect 6656 13416 9404 13444
rect 9398 13404 9404 13416
rect 9456 13444 9462 13456
rect 9582 13444 9588 13456
rect 9456 13416 9588 13444
rect 9456 13404 9462 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 19426 13404 19432 13456
rect 19484 13404 19490 13456
rect 22112 13416 24992 13444
rect 7190 13376 7196 13388
rect 5736 13348 7196 13376
rect 5736 13320 5764 13348
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 10873 13379 10931 13385
rect 10873 13345 10885 13379
rect 10919 13376 10931 13379
rect 11882 13376 11888 13388
rect 10919 13348 11888 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12897 13379 12955 13385
rect 12897 13345 12909 13379
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4304 13280 4629 13308
rect 4304 13268 4310 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5534 13308 5540 13320
rect 5491 13280 5540 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 5534 13268 5540 13280
rect 5592 13268 5598 13320
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 6546 13268 6552 13320
rect 6604 13268 6610 13320
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 7852 13240 7880 13271
rect 8018 13268 8024 13320
rect 8076 13268 8082 13320
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10594 13308 10600 13320
rect 10284 13280 10600 13308
rect 10284 13268 10290 13280
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13277 11207 13311
rect 12912 13308 12940 13339
rect 13630 13336 13636 13388
rect 13688 13336 13694 13388
rect 15194 13336 15200 13388
rect 15252 13336 15258 13388
rect 16206 13336 16212 13388
rect 16264 13376 16270 13388
rect 17405 13379 17463 13385
rect 16264 13348 16896 13376
rect 16264 13336 16270 13348
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12912 13280 13369 13308
rect 11149 13271 11207 13277
rect 13357 13277 13369 13280
rect 13403 13308 13415 13311
rect 14550 13308 14556 13320
rect 13403 13280 14556 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 11164 13240 11192 13271
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15286 13308 15292 13320
rect 15151 13280 15292 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16666 13308 16672 13320
rect 15396 13280 16672 13308
rect 7024 13212 8708 13240
rect 11164 13212 11284 13240
rect 7024 13181 7052 13212
rect 8680 13184 8708 13212
rect 11256 13184 11284 13212
rect 11422 13200 11428 13252
rect 11480 13200 11486 13252
rect 12158 13200 12164 13252
rect 12216 13200 12222 13252
rect 13449 13243 13507 13249
rect 13449 13209 13461 13243
rect 13495 13240 13507 13243
rect 15396 13240 15424 13280
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 16868 13317 16896 13348
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 17770 13376 17776 13388
rect 17451 13348 17776 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 18506 13376 18512 13388
rect 18156 13348 18512 13376
rect 18156 13320 18184 13348
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 19444 13376 19472 13404
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 19444 13348 19533 13376
rect 19521 13345 19533 13348
rect 19567 13345 19579 13379
rect 19521 13339 19579 13345
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 21082 13376 21088 13388
rect 20864 13348 21088 13376
rect 20864 13336 20870 13348
rect 21082 13336 21088 13348
rect 21140 13376 21146 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21140 13348 21833 13376
rect 21140 13336 21146 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 17034 13268 17040 13320
rect 17092 13268 17098 13320
rect 17862 13268 17868 13320
rect 17920 13268 17926 13320
rect 18138 13268 18144 13320
rect 18196 13268 18202 13320
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13308 18475 13311
rect 18874 13308 18880 13320
rect 18463 13280 18880 13308
rect 18463 13277 18475 13280
rect 18417 13271 18475 13277
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13277 19395 13311
rect 19337 13271 19395 13277
rect 16942 13240 16948 13252
rect 13495 13212 15424 13240
rect 15488 13212 16948 13240
rect 13495 13209 13507 13212
rect 13449 13203 13507 13209
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13141 7067 13175
rect 7009 13135 7067 13141
rect 7834 13132 7840 13184
rect 7892 13132 7898 13184
rect 8662 13132 8668 13184
rect 8720 13132 8726 13184
rect 11238 13132 11244 13184
rect 11296 13132 11302 13184
rect 12989 13175 13047 13181
rect 12989 13141 13001 13175
rect 13035 13172 13047 13175
rect 13078 13172 13084 13184
rect 13035 13144 13084 13172
rect 13035 13141 13047 13144
rect 12989 13135 13047 13141
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 15488 13181 15516 13212
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 17880 13240 17908 13268
rect 18322 13240 18328 13252
rect 17880 13212 18328 13240
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 19352 13240 19380 13271
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21177 13311 21235 13317
rect 21177 13308 21189 13311
rect 21048 13280 21189 13308
rect 21048 13268 21054 13280
rect 21177 13277 21189 13280
rect 21223 13308 21235 13311
rect 22112 13308 22140 13416
rect 22186 13336 22192 13388
rect 22244 13336 22250 13388
rect 22278 13336 22284 13388
rect 22336 13336 22342 13388
rect 22373 13379 22431 13385
rect 22373 13345 22385 13379
rect 22419 13376 22431 13379
rect 22738 13376 22744 13388
rect 22419 13348 22744 13376
rect 22419 13345 22431 13348
rect 22373 13339 22431 13345
rect 22738 13336 22744 13348
rect 22796 13336 22802 13388
rect 22830 13336 22836 13388
rect 22888 13376 22894 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22888 13348 23029 13376
rect 22888 13336 22894 13348
rect 23017 13345 23029 13348
rect 23063 13376 23075 13379
rect 23474 13376 23480 13388
rect 23063 13348 23480 13376
rect 23063 13345 23075 13348
rect 23017 13339 23075 13345
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 23842 13336 23848 13388
rect 23900 13376 23906 13388
rect 24762 13376 24768 13388
rect 23900 13348 24768 13376
rect 23900 13336 23906 13348
rect 21223 13280 22140 13308
rect 21223 13277 21235 13280
rect 21177 13271 21235 13277
rect 22462 13268 22468 13320
rect 22520 13268 22526 13320
rect 22925 13311 22983 13317
rect 22925 13277 22937 13311
rect 22971 13308 22983 13311
rect 23385 13311 23443 13317
rect 23385 13308 23397 13311
rect 22971 13280 23397 13308
rect 22971 13277 22983 13280
rect 22925 13271 22983 13277
rect 23385 13277 23397 13280
rect 23431 13277 23443 13311
rect 23385 13271 23443 13277
rect 21358 13240 21364 13252
rect 19352 13212 21364 13240
rect 21358 13200 21364 13212
rect 21416 13240 21422 13252
rect 21637 13243 21695 13249
rect 21637 13240 21649 13243
rect 21416 13212 21649 13240
rect 21416 13200 21422 13212
rect 21637 13209 21649 13212
rect 21683 13240 21695 13243
rect 22940 13240 22968 13271
rect 24026 13268 24032 13320
rect 24084 13268 24090 13320
rect 24228 13317 24256 13348
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 24964 13376 24992 13416
rect 26510 13404 26516 13456
rect 26568 13404 26574 13456
rect 27338 13376 27344 13388
rect 24964 13348 27344 13376
rect 24857 13339 24915 13345
rect 24213 13311 24271 13317
rect 24213 13277 24225 13311
rect 24259 13277 24271 13311
rect 24213 13271 24271 13277
rect 21683 13212 22968 13240
rect 24121 13243 24179 13249
rect 21683 13209 21695 13212
rect 21637 13203 21695 13209
rect 24121 13209 24133 13243
rect 24167 13240 24179 13243
rect 24872 13240 24900 13339
rect 27338 13336 27344 13348
rect 27396 13336 27402 13388
rect 24949 13311 25007 13317
rect 24949 13277 24961 13311
rect 24995 13308 25007 13311
rect 25130 13308 25136 13320
rect 24995 13280 25136 13308
rect 24995 13277 25007 13280
rect 24949 13271 25007 13277
rect 25130 13268 25136 13280
rect 25188 13308 25194 13320
rect 25409 13311 25467 13317
rect 25409 13308 25421 13311
rect 25188 13280 25421 13308
rect 25188 13268 25194 13280
rect 25409 13277 25421 13280
rect 25455 13277 25467 13311
rect 25409 13271 25467 13277
rect 25593 13311 25651 13317
rect 25593 13277 25605 13311
rect 25639 13277 25651 13311
rect 25593 13271 25651 13277
rect 24167 13212 24900 13240
rect 24167 13209 24179 13212
rect 24121 13203 24179 13209
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13141 15531 13175
rect 15473 13135 15531 13141
rect 16850 13132 16856 13184
rect 16908 13132 16914 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 21269 13175 21327 13181
rect 21269 13172 21281 13175
rect 20680 13144 21281 13172
rect 20680 13132 20686 13144
rect 21269 13141 21281 13144
rect 21315 13141 21327 13175
rect 21269 13135 21327 13141
rect 21729 13175 21787 13181
rect 21729 13141 21741 13175
rect 21775 13172 21787 13175
rect 22649 13175 22707 13181
rect 22649 13172 22661 13175
rect 21775 13144 22661 13172
rect 21775 13141 21787 13144
rect 21729 13135 21787 13141
rect 22649 13141 22661 13144
rect 22695 13141 22707 13175
rect 22649 13135 22707 13141
rect 23293 13175 23351 13181
rect 23293 13141 23305 13175
rect 23339 13172 23351 13175
rect 24670 13172 24676 13184
rect 23339 13144 24676 13172
rect 23339 13141 23351 13144
rect 23293 13135 23351 13141
rect 24670 13132 24676 13144
rect 24728 13172 24734 13184
rect 25498 13172 25504 13184
rect 24728 13144 25504 13172
rect 24728 13132 24734 13144
rect 25498 13132 25504 13144
rect 25556 13172 25562 13184
rect 25608 13172 25636 13271
rect 26326 13268 26332 13320
rect 26384 13268 26390 13320
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 26605 13311 26663 13317
rect 26605 13277 26617 13311
rect 26651 13277 26663 13311
rect 26605 13271 26663 13277
rect 26142 13200 26148 13252
rect 26200 13240 26206 13252
rect 26620 13240 26648 13271
rect 26200 13212 26648 13240
rect 26200 13200 26206 13212
rect 25556 13144 25636 13172
rect 25556 13132 25562 13144
rect 1104 13082 30820 13104
rect 1104 13030 5324 13082
rect 5376 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 12752 13082
rect 12804 13030 12816 13082
rect 12868 13030 12880 13082
rect 12932 13030 12944 13082
rect 12996 13030 13008 13082
rect 13060 13030 20180 13082
rect 20232 13030 20244 13082
rect 20296 13030 20308 13082
rect 20360 13030 20372 13082
rect 20424 13030 20436 13082
rect 20488 13030 27608 13082
rect 27660 13030 27672 13082
rect 27724 13030 27736 13082
rect 27788 13030 27800 13082
rect 27852 13030 27864 13082
rect 27916 13030 30820 13082
rect 1104 13008 30820 13030
rect 7098 12928 7104 12980
rect 7156 12928 7162 12980
rect 8754 12968 8760 12980
rect 8404 12940 8760 12968
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 5721 12903 5779 12909
rect 4028 12872 5396 12900
rect 4028 12860 4034 12872
rect 2774 12792 2780 12844
rect 2832 12792 2838 12844
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4212 12804 4353 12832
rect 4212 12792 4218 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 4617 12835 4675 12841
rect 4617 12832 4629 12835
rect 4580 12804 4629 12832
rect 4580 12792 4586 12804
rect 4617 12801 4629 12804
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5368 12841 5396 12872
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 6454 12900 6460 12912
rect 5767 12872 6460 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 7116 12832 7144 12928
rect 8404 12909 8432 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9766 12968 9772 12980
rect 8956 12940 9772 12968
rect 8389 12903 8447 12909
rect 8389 12869 8401 12903
rect 8435 12869 8447 12903
rect 8389 12863 8447 12869
rect 8846 12860 8852 12912
rect 8904 12860 8910 12912
rect 8956 12909 8984 12940
rect 9766 12928 9772 12940
rect 9824 12968 9830 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9824 12940 9873 12968
rect 9824 12928 9830 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 11330 12968 11336 12980
rect 9861 12931 9919 12937
rect 11072 12940 11336 12968
rect 8941 12903 8999 12909
rect 8941 12869 8953 12903
rect 8987 12869 8999 12903
rect 8941 12863 8999 12869
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 11072 12909 11100 12940
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 11480 12940 11621 12968
rect 11480 12928 11486 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 13078 12968 13084 12980
rect 11609 12931 11667 12937
rect 11808 12940 13084 12968
rect 10229 12903 10287 12909
rect 10229 12900 10241 12903
rect 9640 12872 10241 12900
rect 9640 12860 9646 12872
rect 10229 12869 10241 12872
rect 10275 12869 10287 12903
rect 10229 12863 10287 12869
rect 11057 12903 11115 12909
rect 11057 12869 11069 12903
rect 11103 12869 11115 12903
rect 11057 12863 11115 12869
rect 5399 12804 7144 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8711 12835 8769 12841
rect 8711 12832 8723 12835
rect 8352 12804 8723 12832
rect 8352 12792 8358 12804
rect 8711 12801 8723 12804
rect 8757 12801 8769 12835
rect 8711 12795 8769 12801
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9306 12832 9312 12844
rect 9079 12804 9312 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 9456 12804 9505 12832
rect 9456 12792 9462 12804
rect 9493 12801 9505 12804
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9674 12792 9680 12844
rect 9732 12832 9738 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9732 12804 9781 12832
rect 9732 12792 9738 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10042 12792 10048 12844
rect 10100 12792 10106 12844
rect 10594 12792 10600 12844
rect 10652 12832 10658 12844
rect 11808 12841 11836 12940
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 13906 12968 13912 12980
rect 13863 12940 13912 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 13906 12928 13912 12940
rect 13964 12968 13970 12980
rect 13964 12940 15424 12968
rect 13964 12928 13970 12940
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 11940 12872 12112 12900
rect 11940 12860 11946 12872
rect 12084 12841 12112 12872
rect 12158 12860 12164 12912
rect 12216 12860 12222 12912
rect 14550 12900 14556 12912
rect 14292 12872 14556 12900
rect 14292 12841 14320 12872
rect 14550 12860 14556 12872
rect 14608 12860 14614 12912
rect 11333 12835 11391 12841
rect 11333 12832 11345 12835
rect 10652 12804 11345 12832
rect 10652 12792 10658 12804
rect 11333 12801 11345 12804
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11793 12835 11851 12841
rect 11793 12801 11805 12835
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 15396 12841 15424 12940
rect 16666 12928 16672 12980
rect 16724 12928 16730 12980
rect 16850 12928 16856 12980
rect 16908 12928 16914 12980
rect 16942 12928 16948 12980
rect 17000 12928 17006 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17678 12968 17684 12980
rect 17092 12940 17684 12968
rect 17092 12928 17098 12940
rect 17678 12928 17684 12940
rect 17736 12968 17742 12980
rect 17736 12940 17816 12968
rect 17736 12928 17742 12940
rect 16868 12841 16896 12928
rect 16960 12900 16988 12928
rect 17788 12909 17816 12940
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 20036 12940 20085 12968
rect 20036 12928 20042 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 22278 12928 22284 12980
rect 22336 12928 22342 12980
rect 22462 12928 22468 12980
rect 22520 12968 22526 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 22520 12940 25053 12968
rect 22520 12928 22526 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 25590 12928 25596 12980
rect 25648 12928 25654 12980
rect 26418 12928 26424 12980
rect 26476 12928 26482 12980
rect 17155 12903 17213 12909
rect 17155 12900 17167 12903
rect 16960 12872 17167 12900
rect 17155 12869 17167 12872
rect 17201 12869 17213 12903
rect 17773 12903 17831 12909
rect 17155 12863 17213 12869
rect 17420 12872 17724 12900
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 1854 12724 1860 12776
rect 1912 12724 1918 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 2746 12736 6653 12764
rect 1872 12696 1900 12724
rect 2746 12696 2774 12736
rect 6641 12733 6653 12736
rect 6687 12764 6699 12767
rect 7006 12764 7012 12776
rect 6687 12736 7012 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8938 12764 8944 12776
rect 8628 12736 8944 12764
rect 8628 12724 8634 12736
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9582 12724 9588 12776
rect 9640 12724 9646 12776
rect 10502 12764 10508 12776
rect 9692 12736 10508 12764
rect 1872 12668 2774 12696
rect 6086 12656 6092 12708
rect 6144 12656 6150 12708
rect 7024 12696 7052 12724
rect 9692 12696 9720 12736
rect 10502 12724 10508 12736
rect 10560 12764 10566 12776
rect 15013 12767 15071 12773
rect 10560 12736 11284 12764
rect 10560 12724 10566 12736
rect 11256 12708 11284 12736
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15105 12767 15163 12773
rect 15105 12764 15117 12767
rect 15059 12736 15117 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 15105 12733 15117 12736
rect 15151 12733 15163 12767
rect 15105 12727 15163 12733
rect 7024 12668 9720 12696
rect 11238 12656 11244 12708
rect 11296 12656 11302 12708
rect 14829 12699 14887 12705
rect 14829 12696 14841 12699
rect 14108 12668 14841 12696
rect 14108 12640 14136 12668
rect 14829 12665 14841 12668
rect 14875 12665 14887 12699
rect 16960 12696 16988 12795
rect 17052 12764 17080 12795
rect 17126 12764 17132 12776
rect 17052 12736 17132 12764
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 17276 12736 17325 12764
rect 17276 12724 17282 12736
rect 17313 12733 17325 12736
rect 17359 12764 17371 12767
rect 17420 12764 17448 12872
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17696 12832 17724 12872
rect 17773 12869 17785 12903
rect 17819 12869 17831 12903
rect 17773 12863 17831 12869
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 18601 12903 18659 12909
rect 18601 12900 18613 12903
rect 18288 12872 18613 12900
rect 18288 12860 18294 12872
rect 18601 12869 18613 12872
rect 18647 12869 18659 12903
rect 20530 12900 20536 12912
rect 18601 12863 18659 12869
rect 19306 12872 20536 12900
rect 18690 12832 18696 12844
rect 17696 12804 18696 12832
rect 17589 12795 17647 12801
rect 17359 12736 17448 12764
rect 17359 12733 17371 12736
rect 17313 12727 17371 12733
rect 17402 12696 17408 12708
rect 16960 12668 17408 12696
rect 14829 12659 14887 12665
rect 17402 12656 17408 12668
rect 17460 12656 17466 12708
rect 2590 12588 2596 12640
rect 2648 12588 2654 12640
rect 5074 12588 5080 12640
rect 5132 12588 5138 12640
rect 6181 12631 6239 12637
rect 6181 12597 6193 12631
rect 6227 12628 6239 12631
rect 7466 12628 7472 12640
rect 6227 12600 7472 12628
rect 6227 12597 6239 12600
rect 6181 12591 6239 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9309 12631 9367 12637
rect 9309 12597 9321 12631
rect 9355 12628 9367 12631
rect 9398 12628 9404 12640
rect 9355 12600 9404 12628
rect 9355 12597 9367 12600
rect 9309 12591 9367 12597
rect 9398 12588 9404 12600
rect 9456 12588 9462 12640
rect 9766 12588 9772 12640
rect 9824 12588 9830 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 11974 12628 11980 12640
rect 11664 12600 11980 12628
rect 11664 12588 11670 12600
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 14090 12588 14096 12640
rect 14148 12588 14154 12640
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 16206 12588 16212 12640
rect 16264 12628 16270 12640
rect 17604 12628 17632 12795
rect 18690 12792 18696 12804
rect 18748 12832 18754 12844
rect 19306 12832 19334 12872
rect 20530 12860 20536 12872
rect 20588 12900 20594 12912
rect 22296 12900 22324 12928
rect 25958 12900 25964 12912
rect 20588 12872 22324 12900
rect 25424 12872 25820 12900
rect 20588 12860 20594 12872
rect 18748 12804 19334 12832
rect 21637 12835 21695 12841
rect 18748 12792 18754 12804
rect 21637 12801 21649 12835
rect 21683 12801 21695 12835
rect 21637 12795 21695 12801
rect 21652 12764 21680 12795
rect 23198 12792 23204 12844
rect 23256 12792 23262 12844
rect 23477 12835 23535 12841
rect 23477 12801 23489 12835
rect 23523 12832 23535 12835
rect 23566 12832 23572 12844
rect 23523 12804 23572 12832
rect 23523 12801 23535 12804
rect 23477 12795 23535 12801
rect 23014 12764 23020 12776
rect 21652 12736 23020 12764
rect 23014 12724 23020 12736
rect 23072 12764 23078 12776
rect 23492 12764 23520 12795
rect 23566 12792 23572 12804
rect 23624 12792 23630 12844
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 24305 12835 24363 12841
rect 24305 12832 24317 12835
rect 24084 12804 24317 12832
rect 24084 12792 24090 12804
rect 24305 12801 24317 12804
rect 24351 12801 24363 12835
rect 24305 12795 24363 12801
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24489 12835 24547 12841
rect 24489 12832 24501 12835
rect 24443 12804 24501 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24489 12801 24501 12804
rect 24535 12801 24547 12835
rect 24489 12795 24547 12801
rect 24670 12792 24676 12844
rect 24728 12792 24734 12844
rect 25424 12841 25452 12872
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 24903 12804 25421 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25498 12792 25504 12844
rect 25556 12792 25562 12844
rect 25685 12835 25743 12841
rect 25685 12801 25697 12835
rect 25731 12801 25743 12835
rect 25685 12795 25743 12801
rect 23072 12736 23520 12764
rect 23072 12724 23078 12736
rect 16264 12600 17632 12628
rect 16264 12588 16270 12600
rect 21542 12588 21548 12640
rect 21600 12588 21606 12640
rect 24688 12628 24716 12792
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12764 25007 12767
rect 25130 12764 25136 12776
rect 24995 12736 25136 12764
rect 24995 12733 25007 12736
rect 24949 12727 25007 12733
rect 25130 12724 25136 12736
rect 25188 12764 25194 12776
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 25188 12736 25329 12764
rect 25188 12724 25194 12736
rect 25317 12733 25329 12736
rect 25363 12764 25375 12767
rect 25700 12764 25728 12795
rect 25363 12736 25728 12764
rect 25792 12764 25820 12872
rect 25884 12872 25964 12900
rect 25884 12841 25912 12872
rect 25958 12860 25964 12872
rect 26016 12900 26022 12912
rect 26436 12900 26464 12928
rect 26016 12872 26464 12900
rect 26016 12860 26022 12872
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12832 26111 12835
rect 26142 12832 26148 12844
rect 26099 12804 26148 12832
rect 26099 12801 26111 12804
rect 26053 12795 26111 12801
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 25961 12767 26019 12773
rect 25961 12764 25973 12767
rect 25792 12736 25973 12764
rect 25363 12733 25375 12736
rect 25317 12727 25375 12733
rect 25961 12733 25973 12736
rect 26007 12733 26019 12767
rect 25961 12727 26019 12733
rect 25225 12631 25283 12637
rect 25225 12628 25237 12631
rect 24688 12600 25237 12628
rect 25225 12597 25237 12600
rect 25271 12597 25283 12631
rect 25225 12591 25283 12597
rect 1104 12538 30820 12560
rect 1104 12486 4664 12538
rect 4716 12486 4728 12538
rect 4780 12486 4792 12538
rect 4844 12486 4856 12538
rect 4908 12486 4920 12538
rect 4972 12486 12092 12538
rect 12144 12486 12156 12538
rect 12208 12486 12220 12538
rect 12272 12486 12284 12538
rect 12336 12486 12348 12538
rect 12400 12486 19520 12538
rect 19572 12486 19584 12538
rect 19636 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 26948 12538
rect 27000 12486 27012 12538
rect 27064 12486 27076 12538
rect 27128 12486 27140 12538
rect 27192 12486 27204 12538
rect 27256 12486 30820 12538
rect 1104 12464 30820 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 2832 12396 3801 12424
rect 2832 12384 2838 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 6748 12396 8064 12424
rect 3988 12328 5212 12356
rect 3988 12300 4016 12328
rect 5184 12300 5212 12328
rect 1854 12248 1860 12300
rect 1912 12248 1918 12300
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2590 12288 2596 12300
rect 2179 12260 2596 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 3970 12248 3976 12300
rect 4028 12248 4034 12300
rect 4338 12248 4344 12300
rect 4396 12248 4402 12300
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 5074 12288 5080 12300
rect 4939 12260 5080 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5166 12248 5172 12300
rect 5224 12248 5230 12300
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3786 12180 3792 12232
rect 3844 12220 3850 12232
rect 4356 12220 4384 12248
rect 3844 12192 4384 12220
rect 4709 12223 4767 12229
rect 3844 12180 3850 12192
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3620 12124 4169 12152
rect 3620 12093 3648 12124
rect 4157 12121 4169 12124
rect 4203 12152 4215 12155
rect 4724 12152 4752 12183
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 6472 12152 6500 12180
rect 4203 12124 6500 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 3605 12087 3663 12093
rect 3605 12053 3617 12087
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 6748 12084 6776 12396
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 8036 12356 8064 12396
rect 8294 12384 8300 12436
rect 8352 12384 8358 12436
rect 9214 12424 9220 12436
rect 8404 12396 9220 12424
rect 8404 12356 8432 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 9364 12396 9413 12424
rect 9364 12384 9370 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9674 12424 9680 12436
rect 9401 12387 9459 12393
rect 9646 12384 9680 12424
rect 9732 12424 9738 12436
rect 10042 12424 10048 12436
rect 9732 12396 10048 12424
rect 9732 12384 9738 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 14182 12424 14188 12436
rect 13464 12396 14188 12424
rect 7524 12328 7972 12356
rect 8036 12328 8432 12356
rect 7524 12316 7530 12328
rect 7484 12229 7512 12316
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 7944 12288 7972 12328
rect 8478 12297 8484 12300
rect 8461 12291 8484 12297
rect 7944 12260 8064 12288
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12189 7527 12223
rect 7469 12183 7527 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 8036 12220 8064 12260
rect 8461 12257 8473 12291
rect 8461 12251 8484 12257
rect 8478 12248 8484 12251
rect 8536 12248 8542 12300
rect 9646 12288 9674 12384
rect 9324 12260 9674 12288
rect 8379 12223 8437 12229
rect 8379 12220 8391 12223
rect 8036 12192 8391 12220
rect 7929 12183 7987 12189
rect 8379 12189 8391 12192
rect 8425 12189 8437 12223
rect 8379 12183 8437 12189
rect 4295 12056 6776 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7024 12084 7052 12183
rect 7285 12155 7343 12161
rect 7285 12121 7297 12155
rect 7331 12152 7343 12155
rect 7650 12152 7656 12164
rect 7331 12124 7656 12152
rect 7331 12121 7343 12124
rect 7285 12115 7343 12121
rect 7650 12112 7656 12124
rect 7708 12152 7714 12164
rect 7944 12152 7972 12183
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9324 12229 9352 12260
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 9582 12180 9588 12232
rect 9640 12180 9646 12232
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 13464 12229 13492 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 21358 12384 21364 12436
rect 21416 12384 21422 12436
rect 13817 12359 13875 12365
rect 13817 12325 13829 12359
rect 13863 12325 13875 12359
rect 18049 12359 18107 12365
rect 18049 12356 18061 12359
rect 13817 12319 13875 12325
rect 17144 12328 18061 12356
rect 13538 12248 13544 12300
rect 13596 12248 13602 12300
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 7708 12124 7972 12152
rect 13556 12152 13584 12248
rect 13832 12220 13860 12319
rect 17144 12300 17172 12328
rect 18049 12325 18061 12328
rect 18095 12325 18107 12359
rect 18049 12319 18107 12325
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15562 12288 15568 12300
rect 14967 12260 15568 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 19334 12248 19340 12300
rect 19392 12288 19398 12300
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19392 12260 19625 12288
rect 19392 12248 19398 12260
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 19978 12288 19984 12300
rect 19659 12260 19984 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 13832 12192 14841 12220
rect 14829 12189 14841 12192
rect 14875 12220 14887 12223
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 14875 12192 15301 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 16206 12180 16212 12232
rect 16264 12220 16270 12232
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 16264 12192 16865 12220
rect 16264 12180 16270 12192
rect 16853 12189 16865 12192
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17083 12192 17325 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17052 12152 17080 12183
rect 17494 12180 17500 12232
rect 17552 12180 17558 12232
rect 18785 12223 18843 12229
rect 18785 12220 18797 12223
rect 18708 12192 18797 12220
rect 13556 12124 17080 12152
rect 17221 12155 17279 12161
rect 7708 12112 7714 12124
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 17267 12124 17816 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 17788 12096 17816 12124
rect 18708 12096 18736 12192
rect 18785 12189 18797 12192
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 19061 12223 19119 12229
rect 19061 12189 19073 12223
rect 19107 12220 19119 12223
rect 19242 12220 19248 12232
rect 19107 12192 19248 12220
rect 19107 12189 19119 12192
rect 19061 12183 19119 12189
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 21542 12220 21548 12232
rect 21022 12192 21548 12220
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21726 12180 21732 12232
rect 21784 12180 21790 12232
rect 23014 12180 23020 12232
rect 23072 12180 23078 12232
rect 19889 12155 19947 12161
rect 19889 12121 19901 12155
rect 19935 12152 19947 12155
rect 19978 12152 19984 12164
rect 19935 12124 19984 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 6972 12056 8585 12084
rect 6972 12044 6978 12056
rect 8573 12053 8585 12056
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 9674 12044 9680 12096
rect 9732 12044 9738 12096
rect 15194 12044 15200 12096
rect 15252 12044 15258 12096
rect 15378 12044 15384 12096
rect 15436 12044 15442 12096
rect 17310 12044 17316 12096
rect 17368 12044 17374 12096
rect 17770 12044 17776 12096
rect 17828 12044 17834 12096
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 21910 12044 21916 12096
rect 21968 12044 21974 12096
rect 23014 12044 23020 12096
rect 23072 12084 23078 12096
rect 23109 12087 23167 12093
rect 23109 12084 23121 12087
rect 23072 12056 23121 12084
rect 23072 12044 23078 12056
rect 23109 12053 23121 12056
rect 23155 12053 23167 12087
rect 23109 12047 23167 12053
rect 1104 11994 30820 12016
rect 1104 11942 5324 11994
rect 5376 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 12752 11994
rect 12804 11942 12816 11994
rect 12868 11942 12880 11994
rect 12932 11942 12944 11994
rect 12996 11942 13008 11994
rect 13060 11942 20180 11994
rect 20232 11942 20244 11994
rect 20296 11942 20308 11994
rect 20360 11942 20372 11994
rect 20424 11942 20436 11994
rect 20488 11942 27608 11994
rect 27660 11942 27672 11994
rect 27724 11942 27736 11994
rect 27788 11942 27800 11994
rect 27852 11942 27864 11994
rect 27916 11942 30820 11994
rect 1104 11920 30820 11942
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 3602 11840 3608 11892
rect 3660 11840 3666 11892
rect 5166 11840 5172 11892
rect 5224 11840 5230 11892
rect 6454 11840 6460 11892
rect 6512 11840 6518 11892
rect 6914 11840 6920 11892
rect 6972 11840 6978 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9969 11883 10027 11889
rect 9969 11880 9981 11883
rect 9732 11852 9981 11880
rect 9732 11840 9738 11852
rect 9969 11849 9981 11852
rect 10015 11849 10027 11883
rect 9969 11843 10027 11849
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 10836 11852 15148 11880
rect 10836 11840 10842 11852
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3620 11744 3648 11840
rect 3384 11716 3648 11744
rect 5184 11744 5212 11840
rect 6472 11753 6500 11840
rect 9769 11815 9827 11821
rect 9769 11781 9781 11815
rect 9815 11812 9827 11815
rect 10134 11812 10140 11824
rect 9815 11784 10140 11812
rect 9815 11781 9827 11784
rect 9769 11775 9827 11781
rect 10134 11772 10140 11784
rect 10192 11772 10198 11824
rect 12434 11772 12440 11824
rect 12492 11772 12498 11824
rect 14182 11812 14188 11824
rect 13832 11784 14188 11812
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5184 11716 5457 11744
rect 3384 11704 3390 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 11146 11704 11152 11756
rect 11204 11704 11210 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11296 11716 11529 11744
rect 11296 11704 11302 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 13446 11744 13452 11756
rect 11517 11707 11575 11713
rect 13280 11716 13452 11744
rect 5166 11636 5172 11688
rect 5224 11636 5230 11688
rect 13280 11685 13308 11716
rect 13446 11704 13452 11716
rect 13504 11744 13510 11756
rect 13832 11753 13860 11784
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13504 11716 13829 11744
rect 13504 11704 13510 11716
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 15120 11744 15148 11852
rect 15194 11840 15200 11892
rect 15252 11840 15258 11892
rect 17405 11883 17463 11889
rect 17405 11849 17417 11883
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 15212 11812 15240 11840
rect 16807 11815 16865 11821
rect 16807 11812 16819 11815
rect 15212 11784 16819 11812
rect 16807 11781 16819 11784
rect 16853 11781 16865 11815
rect 16807 11775 16865 11781
rect 16942 11772 16948 11824
rect 17000 11772 17006 11824
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17420 11812 17448 11843
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 20036 11852 20085 11880
rect 20036 11840 20042 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11880 21695 11883
rect 21726 11880 21732 11892
rect 21683 11852 21732 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 21968 11852 22324 11880
rect 21968 11840 21974 11852
rect 22296 11821 22324 11852
rect 22281 11815 22339 11821
rect 17083 11784 19840 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15120 11716 16681 11744
rect 13817 11707 13875 11713
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17310 11744 17316 11756
rect 17175 11716 17316 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11348 11648 11805 11676
rect 6178 11568 6184 11620
rect 6236 11608 6242 11620
rect 10042 11608 10048 11620
rect 6236 11580 10048 11608
rect 6236 11568 6242 11580
rect 6748 11549 6776 11580
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 11348 11617 11376 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11645 13323 11679
rect 16684 11676 16712 11707
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 17402 11704 17408 11756
rect 17460 11744 17466 11756
rect 17589 11747 17647 11753
rect 17589 11744 17601 11747
rect 17460 11716 17601 11744
rect 17460 11704 17466 11716
rect 17589 11713 17601 11716
rect 17635 11744 17647 11747
rect 17678 11744 17684 11756
rect 17635 11716 17684 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11713 17831 11747
rect 17773 11707 17831 11713
rect 17218 11676 17224 11688
rect 16684 11648 17224 11676
rect 13265 11639 13323 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 11333 11611 11391 11617
rect 11333 11577 11345 11611
rect 11379 11577 11391 11611
rect 11333 11571 11391 11577
rect 17788 11552 17816 11707
rect 18141 11679 18199 11685
rect 18141 11645 18153 11679
rect 18187 11676 18199 11679
rect 18325 11679 18383 11685
rect 18187 11648 18276 11676
rect 18187 11645 18199 11648
rect 18141 11639 18199 11645
rect 18248 11552 18276 11648
rect 18325 11645 18337 11679
rect 18371 11645 18383 11679
rect 18325 11639 18383 11645
rect 18340 11552 18368 11639
rect 18690 11636 18696 11688
rect 18748 11636 18754 11688
rect 19812 11676 19840 11784
rect 20088 11784 22048 11812
rect 20088 11756 20116 11784
rect 20070 11704 20076 11756
rect 20128 11704 20134 11756
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20622 11744 20628 11756
rect 20303 11716 20628 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 22020 11753 22048 11784
rect 22281 11781 22293 11815
rect 22327 11781 22339 11815
rect 22281 11775 22339 11781
rect 23014 11772 23020 11824
rect 23072 11772 23078 11824
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11713 21327 11747
rect 21269 11707 21327 11713
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 20990 11676 20996 11688
rect 19812 11648 20996 11676
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21082 11636 21088 11688
rect 21140 11636 21146 11688
rect 21174 11636 21180 11688
rect 21232 11636 21238 11688
rect 21284 11676 21312 11707
rect 23934 11704 23940 11756
rect 23992 11744 23998 11756
rect 24213 11747 24271 11753
rect 24213 11744 24225 11747
rect 23992 11716 24225 11744
rect 23992 11704 23998 11716
rect 24213 11713 24225 11716
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 23753 11679 23811 11685
rect 23753 11676 23765 11679
rect 21284 11648 23765 11676
rect 6733 11543 6791 11549
rect 6733 11509 6745 11543
rect 6779 11540 6791 11543
rect 6779 11512 6813 11540
rect 6779 11509 6791 11512
rect 6733 11503 6791 11509
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 9674 11540 9680 11552
rect 9456 11512 9680 11540
rect 9456 11500 9462 11512
rect 9674 11500 9680 11512
rect 9732 11540 9738 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9732 11512 9965 11540
rect 9732 11500 9738 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10134 11500 10140 11552
rect 10192 11500 10198 11552
rect 13354 11500 13360 11552
rect 13412 11500 13418 11552
rect 13538 11500 13544 11552
rect 13596 11500 13602 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 17313 11543 17371 11549
rect 17313 11540 17325 11543
rect 14976 11512 17325 11540
rect 14976 11500 14982 11512
rect 17313 11509 17325 11512
rect 17359 11509 17371 11543
rect 17313 11503 17371 11509
rect 17770 11500 17776 11552
rect 17828 11500 17834 11552
rect 18230 11500 18236 11552
rect 18288 11500 18294 11552
rect 18322 11500 18328 11552
rect 18380 11500 18386 11552
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 19426 11540 19432 11552
rect 18472 11512 19432 11540
rect 18472 11500 18478 11512
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 21284 11540 21312 11648
rect 23753 11645 23765 11648
rect 23799 11676 23811 11679
rect 23842 11676 23848 11688
rect 23799 11648 23848 11676
rect 23799 11645 23811 11648
rect 23753 11639 23811 11645
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 20036 11512 21312 11540
rect 20036 11500 20042 11512
rect 24302 11500 24308 11552
rect 24360 11500 24366 11552
rect 1104 11450 30820 11472
rect 1104 11398 4664 11450
rect 4716 11398 4728 11450
rect 4780 11398 4792 11450
rect 4844 11398 4856 11450
rect 4908 11398 4920 11450
rect 4972 11398 12092 11450
rect 12144 11398 12156 11450
rect 12208 11398 12220 11450
rect 12272 11398 12284 11450
rect 12336 11398 12348 11450
rect 12400 11398 19520 11450
rect 19572 11398 19584 11450
rect 19636 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 26948 11450
rect 27000 11398 27012 11450
rect 27064 11398 27076 11450
rect 27128 11398 27140 11450
rect 27192 11398 27204 11450
rect 27256 11398 30820 11450
rect 1104 11376 30820 11398
rect 1854 11296 1860 11348
rect 1912 11296 1918 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 9582 11336 9588 11348
rect 6880 11308 9588 11336
rect 6880 11296 6886 11308
rect 9582 11296 9588 11308
rect 9640 11296 9646 11348
rect 10134 11296 10140 11348
rect 10192 11296 10198 11348
rect 11146 11296 11152 11348
rect 11204 11296 11210 11348
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12434 11336 12440 11348
rect 12023 11308 12440 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 14918 11336 14924 11348
rect 12728 11308 14924 11336
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 1872 11200 1900 11296
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11268 7159 11271
rect 9122 11268 9128 11280
rect 7147 11240 9128 11268
rect 7147 11237 7159 11240
rect 7101 11231 7159 11237
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 1811 11172 1900 11200
rect 3513 11203 3571 11209
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 3559 11172 4200 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 2038 11024 2044 11076
rect 2096 11024 2102 11076
rect 4172 11073 4200 11172
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 4632 11172 8800 11200
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4632 11132 4660 11172
rect 4295 11104 4660 11132
rect 4709 11135 4767 11141
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4724 11064 4752 11095
rect 4203 11036 4844 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 4816 10996 4844 11036
rect 4890 11024 4896 11076
rect 4948 11024 4954 11076
rect 5000 11036 5580 11064
rect 5000 10996 5028 11036
rect 4816 10968 5028 10996
rect 5552 10996 5580 11036
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 5776 11036 6561 11064
rect 5776 11024 5782 11036
rect 6549 11033 6561 11036
rect 6595 11033 6607 11067
rect 6549 11027 6607 11033
rect 6656 11008 6684 11095
rect 7374 11092 7380 11144
rect 7432 11092 7438 11144
rect 7650 11092 7656 11144
rect 7708 11092 7714 11144
rect 8294 11092 8300 11144
rect 8352 11092 8358 11144
rect 8386 11092 8392 11144
rect 8444 11092 8450 11144
rect 8665 11067 8723 11073
rect 8665 11033 8677 11067
rect 8711 11033 8723 11067
rect 8772 11064 8800 11172
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10042 11132 10048 11144
rect 9999 11104 10048 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10152 11132 10180 11296
rect 10321 11271 10379 11277
rect 10321 11237 10333 11271
rect 10367 11237 10379 11271
rect 11164 11268 11192 11296
rect 12161 11271 12219 11277
rect 12161 11268 12173 11271
rect 11164 11240 12173 11268
rect 10321 11231 10379 11237
rect 12161 11237 12173 11240
rect 12207 11237 12219 11271
rect 12728 11268 12756 11308
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 15528 11308 15761 11336
rect 15528 11296 15534 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 19337 11339 19395 11345
rect 19337 11336 19349 11339
rect 17000 11308 19349 11336
rect 17000 11296 17006 11308
rect 19337 11305 19349 11308
rect 19383 11305 19395 11339
rect 21082 11336 21088 11348
rect 19337 11299 19395 11305
rect 19628 11308 21088 11336
rect 12161 11231 12219 11237
rect 12636 11240 12756 11268
rect 10336 11200 10364 11231
rect 12636 11209 12664 11240
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 13596 11240 13645 11268
rect 13596 11228 13602 11240
rect 13633 11237 13645 11240
rect 13679 11237 13691 11271
rect 13633 11231 13691 11237
rect 15838 11228 15844 11280
rect 15896 11228 15902 11280
rect 17144 11240 19564 11268
rect 12621 11203 12679 11209
rect 10336 11172 10916 11200
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10152 11104 10609 11132
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 10888 11141 10916 11172
rect 12621 11169 12633 11203
rect 12667 11169 12679 11203
rect 12621 11163 12679 11169
rect 12805 11203 12863 11209
rect 12805 11169 12817 11203
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 13446 11200 13452 11212
rect 13403 11172 13452 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11101 10931 11135
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 10873 11095 10931 11101
rect 11808 11104 11897 11132
rect 11808 11076 11836 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 12820 11132 12848 11163
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 15010 11160 15016 11212
rect 15068 11160 15074 11212
rect 13630 11132 13636 11144
rect 12820 11104 13636 11132
rect 11885 11095 11943 11101
rect 13630 11092 13636 11104
rect 13688 11132 13694 11144
rect 15028 11132 15056 11160
rect 13688 11104 15056 11132
rect 15565 11135 15623 11141
rect 13688 11092 13694 11104
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15856 11132 15884 11228
rect 17144 11144 17172 11240
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 19337 11203 19395 11209
rect 19337 11200 19349 11203
rect 17828 11172 19349 11200
rect 17828 11160 17834 11172
rect 19337 11169 19349 11172
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 17126 11132 17132 11144
rect 15856 11104 17132 11132
rect 15565 11095 15623 11101
rect 10413 11067 10471 11073
rect 10413 11064 10425 11067
rect 8772 11036 10425 11064
rect 8665 11027 8723 11033
rect 10413 11033 10425 11036
rect 10459 11033 10471 11067
rect 10413 11027 10471 11033
rect 6638 10996 6644 11008
rect 5552 10968 6644 10996
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 8680 10996 8708 11027
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 12529 11067 12587 11073
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 13446 11064 13452 11076
rect 12575 11036 13452 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 13446 11024 13452 11036
rect 13504 11024 13510 11076
rect 15580 11008 15608 11095
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18874 11092 18880 11144
rect 18932 11092 18938 11144
rect 19536 11141 19564 11240
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 16209 11067 16267 11073
rect 16209 11033 16221 11067
rect 16255 11064 16267 11067
rect 16482 11064 16488 11076
rect 16255 11036 16488 11064
rect 16255 11033 16267 11036
rect 16209 11027 16267 11033
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 16942 11024 16948 11076
rect 17000 11024 17006 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 17402 11064 17408 11076
rect 17359 11036 17408 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 17402 11024 17408 11036
rect 17460 11024 17466 11076
rect 18141 11067 18199 11073
rect 18141 11033 18153 11067
rect 18187 11064 18199 11067
rect 18322 11064 18328 11076
rect 18187 11036 18328 11064
rect 18187 11033 18199 11036
rect 18141 11027 18199 11033
rect 18322 11024 18328 11036
rect 18380 11024 18386 11076
rect 18892 11064 18920 11092
rect 19260 11064 19288 11095
rect 19628 11064 19656 11308
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21232 11308 22017 11336
rect 21232 11296 21238 11308
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 25038 11336 25044 11348
rect 24360 11308 25044 11336
rect 24360 11296 24366 11308
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 25130 11296 25136 11348
rect 25188 11296 25194 11348
rect 25317 11339 25375 11345
rect 25317 11305 25329 11339
rect 25363 11305 25375 11339
rect 25317 11299 25375 11305
rect 19705 11271 19763 11277
rect 19705 11237 19717 11271
rect 19751 11268 19763 11271
rect 21818 11268 21824 11280
rect 19751 11240 21824 11268
rect 19751 11237 19763 11240
rect 19705 11231 19763 11237
rect 21818 11228 21824 11240
rect 21876 11268 21882 11280
rect 23934 11268 23940 11280
rect 21876 11240 22324 11268
rect 21876 11228 21882 11240
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22296 11141 22324 11240
rect 23768 11240 23940 11268
rect 23768 11209 23796 11240
rect 23934 11228 23940 11240
rect 23992 11228 23998 11280
rect 25332 11268 25360 11299
rect 24044 11240 25360 11268
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11169 23811 11203
rect 23753 11163 23811 11169
rect 22281 11135 22339 11141
rect 22281 11101 22293 11135
rect 22327 11101 22339 11135
rect 22281 11095 22339 11101
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 22646 11092 22652 11144
rect 22704 11132 22710 11144
rect 23474 11132 23480 11144
rect 22704 11104 23480 11132
rect 22704 11092 22710 11104
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 24044 11132 24072 11240
rect 24854 11200 24860 11212
rect 24780 11172 24860 11200
rect 23952 11104 24072 11132
rect 18892 11036 19104 11064
rect 19260 11036 19656 11064
rect 8628 10968 8708 10996
rect 8628 10956 8634 10968
rect 13814 10956 13820 11008
rect 13872 10956 13878 11008
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 15105 10999 15163 11005
rect 15105 10996 15117 10999
rect 14884 10968 15117 10996
rect 14884 10956 14890 10968
rect 15105 10965 15117 10968
rect 15151 10965 15163 10999
rect 15105 10959 15163 10965
rect 15562 10956 15568 11008
rect 15620 10956 15626 11008
rect 19076 10996 19104 11036
rect 19886 11024 19892 11076
rect 19944 11064 19950 11076
rect 20165 11067 20223 11073
rect 20165 11064 20177 11067
rect 19944 11036 20177 11064
rect 19944 11024 19950 11036
rect 20165 11033 20177 11036
rect 20211 11033 20223 11067
rect 20165 11027 20223 11033
rect 21818 11024 21824 11076
rect 21876 11024 21882 11076
rect 22511 11067 22569 11073
rect 22511 11033 22523 11067
rect 22557 11064 22569 11067
rect 23952 11064 23980 11104
rect 24486 11092 24492 11144
rect 24544 11092 24550 11144
rect 24670 11141 24676 11144
rect 24637 11135 24676 11141
rect 24637 11101 24649 11135
rect 24637 11095 24676 11101
rect 24670 11092 24676 11095
rect 24728 11092 24734 11144
rect 24780 11141 24808 11172
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 25038 11160 25044 11212
rect 25096 11160 25102 11212
rect 25498 11160 25504 11212
rect 25556 11160 25562 11212
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 24954 11135 25012 11141
rect 24954 11101 24966 11135
rect 25000 11132 25012 11135
rect 25056 11132 25084 11160
rect 25000 11104 25084 11132
rect 25593 11135 25651 11141
rect 25000 11101 25012 11104
rect 24954 11095 25012 11101
rect 25593 11101 25605 11135
rect 25639 11101 25651 11135
rect 25593 11095 25651 11101
rect 24857 11067 24915 11073
rect 24857 11064 24869 11067
rect 22557 11036 23980 11064
rect 24044 11036 24869 11064
rect 22557 11033 22569 11036
rect 22511 11027 22569 11033
rect 20070 10996 20076 11008
rect 19076 10968 20076 10996
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 20622 10956 20628 11008
rect 20680 10996 20686 11008
rect 23198 10996 23204 11008
rect 20680 10968 23204 10996
rect 20680 10956 20686 10968
rect 23198 10956 23204 10968
rect 23256 10956 23262 11008
rect 23842 10956 23848 11008
rect 23900 10996 23906 11008
rect 24044 10996 24072 11036
rect 24857 11033 24869 11036
rect 24903 11033 24915 11067
rect 24857 11027 24915 11033
rect 23900 10968 24072 10996
rect 24213 10999 24271 11005
rect 23900 10956 23906 10968
rect 24213 10965 24225 10999
rect 24259 10996 24271 10999
rect 25406 10996 25412 11008
rect 24259 10968 25412 10996
rect 24259 10965 24271 10968
rect 24213 10959 24271 10965
rect 25406 10956 25412 10968
rect 25464 10996 25470 11008
rect 25608 10996 25636 11095
rect 25464 10968 25636 10996
rect 25464 10956 25470 10968
rect 1104 10906 30820 10928
rect 1104 10854 5324 10906
rect 5376 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 12752 10906
rect 12804 10854 12816 10906
rect 12868 10854 12880 10906
rect 12932 10854 12944 10906
rect 12996 10854 13008 10906
rect 13060 10854 20180 10906
rect 20232 10854 20244 10906
rect 20296 10854 20308 10906
rect 20360 10854 20372 10906
rect 20424 10854 20436 10906
rect 20488 10854 27608 10906
rect 27660 10854 27672 10906
rect 27724 10854 27736 10906
rect 27788 10854 27800 10906
rect 27852 10854 27864 10906
rect 27916 10854 30820 10906
rect 1104 10832 30820 10854
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2096 10764 2697 10792
rect 2096 10752 2102 10764
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3200 10764 3249 10792
rect 3200 10752 3206 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 3237 10755 3295 10761
rect 3786 10752 3792 10804
rect 3844 10752 3850 10804
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4028 10764 5304 10792
rect 4028 10752 4034 10764
rect 3804 10724 3832 10752
rect 2884 10696 3832 10724
rect 2884 10665 2912 10696
rect 4890 10684 4896 10736
rect 4948 10684 4954 10736
rect 5276 10724 5304 10764
rect 7374 10752 7380 10804
rect 7432 10752 7438 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7708 10764 7757 10792
rect 7708 10752 7714 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 8021 10795 8079 10801
rect 8021 10761 8033 10795
rect 8067 10792 8079 10795
rect 8386 10792 8392 10804
rect 8067 10764 8392 10792
rect 8067 10761 8079 10764
rect 8021 10755 8079 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 13354 10752 13360 10804
rect 13412 10752 13418 10804
rect 15102 10792 15108 10804
rect 14200 10764 15108 10792
rect 5718 10724 5724 10736
rect 5276 10696 5724 10724
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 3326 10616 3332 10668
rect 3384 10616 3390 10668
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 4172 10520 4200 10616
rect 4448 10588 4476 10619
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4580 10628 4721 10656
rect 4580 10616 4586 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 4816 10588 4844 10616
rect 4908 10597 4936 10684
rect 5460 10665 5488 10696
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 4448 10560 4844 10588
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 5000 10520 5028 10619
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6822 10616 6828 10668
rect 6880 10616 6886 10668
rect 7392 10656 7420 10752
rect 8665 10727 8723 10733
rect 8665 10724 8677 10727
rect 8312 10696 8677 10724
rect 8312 10668 8340 10696
rect 8665 10693 8677 10696
rect 8711 10693 8723 10727
rect 9214 10724 9220 10736
rect 8665 10687 8723 10693
rect 8772 10696 9220 10724
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7392 10628 7665 10656
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 7975 10628 8217 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 5166 10548 5172 10600
rect 5224 10548 5230 10600
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 6840 10588 6868 10616
rect 6779 10560 6868 10588
rect 7469 10591 7527 10597
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 7469 10557 7481 10591
rect 7515 10557 7527 10591
rect 8220 10588 8248 10619
rect 8294 10616 8300 10668
rect 8352 10616 8358 10668
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10656 8631 10659
rect 8772 10656 8800 10696
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 10152 10696 10333 10724
rect 8619 10628 8800 10656
rect 8619 10625 8631 10628
rect 8573 10619 8631 10625
rect 8404 10588 8432 10616
rect 8220 10560 8432 10588
rect 8496 10588 8524 10619
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 10152 10665 10180 10696
rect 10321 10693 10333 10696
rect 10367 10693 10379 10727
rect 10321 10687 10379 10693
rect 9493 10659 9551 10665
rect 9493 10625 9505 10659
rect 9539 10656 9551 10659
rect 9585 10659 9643 10665
rect 9585 10656 9597 10659
rect 9539 10628 9597 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 9585 10625 9597 10628
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 8496 10560 8984 10588
rect 7469 10551 7527 10557
rect 5074 10520 5080 10532
rect 4172 10492 5080 10520
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 6181 10523 6239 10529
rect 6181 10489 6193 10523
rect 6227 10520 6239 10523
rect 6748 10520 6776 10551
rect 6227 10492 6776 10520
rect 7484 10520 7512 10551
rect 8956 10520 8984 10560
rect 9030 10548 9036 10600
rect 9088 10548 9094 10600
rect 9140 10588 9168 10616
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9140 10560 9873 10588
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10244 10588 10272 10619
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12805 10659 12863 10665
rect 12805 10656 12817 10659
rect 12676 10628 12817 10656
rect 12676 10616 12682 10628
rect 12805 10625 12817 10628
rect 12851 10625 12863 10659
rect 13372 10656 13400 10752
rect 13633 10727 13691 10733
rect 13633 10693 13645 10727
rect 13679 10724 13691 10727
rect 14093 10727 14151 10733
rect 14093 10724 14105 10727
rect 13679 10696 14105 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 14093 10693 14105 10696
rect 14139 10693 14151 10727
rect 14093 10687 14151 10693
rect 13449 10659 13507 10665
rect 13449 10656 13461 10659
rect 13372 10628 13461 10656
rect 12805 10619 12863 10625
rect 13449 10625 13461 10628
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13872 10628 13921 10656
rect 13872 10616 13878 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 10100 10560 10272 10588
rect 10100 10548 10106 10560
rect 9677 10523 9735 10529
rect 9677 10520 9689 10523
rect 7484 10492 8524 10520
rect 8956 10492 9689 10520
rect 6227 10489 6239 10492
rect 6181 10483 6239 10489
rect 7926 10412 7932 10464
rect 7984 10412 7990 10464
rect 8496 10452 8524 10492
rect 9677 10489 9689 10492
rect 9723 10489 9735 10523
rect 10244 10520 10272 10560
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 14200 10588 14228 10764
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15286 10752 15292 10804
rect 15344 10752 15350 10804
rect 15378 10752 15384 10804
rect 15436 10752 15442 10804
rect 17126 10752 17132 10804
rect 17184 10752 17190 10804
rect 18506 10752 18512 10804
rect 18564 10792 18570 10804
rect 19978 10792 19984 10804
rect 18564 10764 19984 10792
rect 18564 10752 18570 10764
rect 15396 10724 15424 10752
rect 14660 10696 15424 10724
rect 17144 10724 17172 10752
rect 17144 10696 17724 10724
rect 14660 10665 14688 10696
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14369 10659 14427 10665
rect 14369 10625 14381 10659
rect 14415 10625 14427 10659
rect 14369 10619 14427 10625
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 14553 10619 14611 10625
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 15470 10656 15476 10668
rect 14875 10628 15476 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 12943 10560 14228 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 9677 10483 9735 10489
rect 9876 10492 10272 10520
rect 13817 10523 13875 10529
rect 8846 10452 8852 10464
rect 8496 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10452 8910 10464
rect 9876 10452 9904 10492
rect 13817 10489 13829 10523
rect 13863 10520 13875 10523
rect 13906 10520 13912 10532
rect 13863 10492 13912 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 8904 10424 9904 10452
rect 8904 10412 8910 10424
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 13170 10412 13176 10464
rect 13228 10412 13234 10464
rect 14292 10452 14320 10619
rect 14384 10520 14412 10619
rect 14568 10588 14596 10619
rect 14844 10588 14872 10619
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 14568 10560 14872 10588
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 14936 10520 14964 10548
rect 14384 10492 14964 10520
rect 15028 10520 15056 10551
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 16316 10588 16344 10619
rect 16942 10616 16948 10668
rect 17000 10616 17006 10668
rect 17310 10616 17316 10668
rect 17368 10616 17374 10668
rect 17696 10665 17724 10696
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17865 10659 17923 10665
rect 17865 10625 17877 10659
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 16482 10588 16488 10600
rect 16316 10560 16488 10588
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 16960 10588 16988 10616
rect 17880 10588 17908 10619
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18012 10628 19073 10656
rect 18012 10616 18018 10628
rect 19061 10625 19073 10628
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19426 10616 19432 10668
rect 19484 10616 19490 10668
rect 19536 10656 19564 10764
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 21361 10795 21419 10801
rect 21361 10761 21373 10795
rect 21407 10792 21419 10795
rect 21407 10764 22094 10792
rect 21407 10761 21419 10764
rect 21361 10755 21419 10761
rect 19886 10684 19892 10736
rect 19944 10684 19950 10736
rect 21818 10684 21824 10736
rect 21876 10684 21882 10736
rect 22066 10724 22094 10764
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22244 10764 22385 10792
rect 22244 10752 22250 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23934 10752 23940 10804
rect 23992 10752 23998 10804
rect 24486 10752 24492 10804
rect 24544 10792 24550 10804
rect 24581 10795 24639 10801
rect 24581 10792 24593 10795
rect 24544 10764 24593 10792
rect 24544 10752 24550 10764
rect 24581 10761 24593 10764
rect 24627 10761 24639 10795
rect 24581 10755 24639 10761
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25225 10795 25283 10801
rect 25225 10792 25237 10795
rect 24912 10764 25237 10792
rect 24912 10752 24918 10764
rect 25225 10761 25237 10764
rect 25271 10761 25283 10795
rect 25225 10755 25283 10761
rect 25406 10752 25412 10804
rect 25464 10752 25470 10804
rect 22281 10727 22339 10733
rect 22066 10696 22140 10724
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19536 10628 19717 10656
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 19904 10597 19932 10684
rect 20070 10616 20076 10668
rect 20128 10616 20134 10668
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10656 20683 10659
rect 21836 10656 21864 10684
rect 20671 10628 21864 10656
rect 20671 10625 20683 10628
rect 20625 10619 20683 10625
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 22112 10656 22140 10696
rect 22281 10693 22293 10727
rect 22327 10724 22339 10727
rect 23952 10724 23980 10752
rect 22327 10696 23980 10724
rect 22327 10693 22339 10696
rect 22281 10687 22339 10693
rect 22388 10665 22416 10696
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22112 10628 22385 10656
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10656 22891 10659
rect 23014 10656 23020 10668
rect 22879 10628 23020 10656
rect 22879 10625 22891 10628
rect 22833 10619 22891 10625
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24121 10659 24179 10665
rect 24121 10656 24133 10659
rect 23900 10628 24133 10656
rect 23900 10616 23906 10628
rect 24121 10625 24133 10628
rect 24167 10625 24179 10659
rect 24121 10619 24179 10625
rect 24213 10659 24271 10665
rect 24213 10625 24225 10659
rect 24259 10656 24271 10659
rect 24302 10656 24308 10668
rect 24259 10628 24308 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10656 24455 10659
rect 24578 10656 24584 10668
rect 24443 10628 24584 10656
rect 24443 10625 24455 10628
rect 24397 10619 24455 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 25424 10665 25452 10752
rect 25409 10659 25467 10665
rect 25409 10625 25421 10659
rect 25455 10625 25467 10659
rect 25409 10619 25467 10625
rect 16960 10560 17908 10588
rect 19889 10591 19947 10597
rect 19889 10557 19901 10591
rect 19935 10557 19947 10591
rect 19889 10551 19947 10557
rect 20349 10591 20407 10597
rect 20349 10557 20361 10591
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 15562 10520 15568 10532
rect 15028 10492 15568 10520
rect 15028 10452 15056 10492
rect 15562 10480 15568 10492
rect 15620 10520 15626 10532
rect 15841 10523 15899 10529
rect 15841 10520 15853 10523
rect 15620 10492 15853 10520
rect 15620 10480 15626 10492
rect 15841 10489 15853 10492
rect 15887 10489 15899 10523
rect 15841 10483 15899 10489
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 17184 10492 17785 10520
rect 17184 10480 17190 10492
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 19242 10480 19248 10532
rect 19300 10520 19306 10532
rect 20364 10520 20392 10551
rect 21082 10548 21088 10600
rect 21140 10548 21146 10600
rect 22738 10597 22744 10600
rect 22189 10591 22247 10597
rect 22189 10557 22201 10591
rect 22235 10588 22247 10591
rect 22695 10591 22744 10597
rect 22695 10588 22707 10591
rect 22235 10560 22707 10588
rect 22235 10557 22247 10560
rect 22189 10551 22247 10557
rect 22695 10557 22707 10560
rect 22741 10557 22744 10591
rect 22695 10551 22744 10557
rect 22738 10548 22744 10551
rect 22796 10548 22802 10600
rect 25314 10548 25320 10600
rect 25372 10588 25378 10600
rect 25593 10591 25651 10597
rect 25593 10588 25605 10591
rect 25372 10560 25605 10588
rect 25372 10548 25378 10560
rect 25593 10557 25605 10560
rect 25639 10557 25651 10591
rect 25593 10551 25651 10557
rect 19300 10492 20392 10520
rect 19300 10480 19306 10492
rect 19904 10464 19932 10492
rect 14292 10424 15056 10452
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 15988 10424 16037 10452
rect 15988 10412 15994 10424
rect 16025 10421 16037 10424
rect 16071 10421 16083 10455
rect 16025 10415 16083 10421
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 19886 10412 19892 10464
rect 19944 10412 19950 10464
rect 21100 10452 21128 10548
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 21100 10424 21833 10452
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 22278 10412 22284 10464
rect 22336 10412 22342 10464
rect 22554 10412 22560 10464
rect 22612 10412 22618 10464
rect 1104 10362 30820 10384
rect 1104 10310 4664 10362
rect 4716 10310 4728 10362
rect 4780 10310 4792 10362
rect 4844 10310 4856 10362
rect 4908 10310 4920 10362
rect 4972 10310 12092 10362
rect 12144 10310 12156 10362
rect 12208 10310 12220 10362
rect 12272 10310 12284 10362
rect 12336 10310 12348 10362
rect 12400 10310 19520 10362
rect 19572 10310 19584 10362
rect 19636 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 26948 10362
rect 27000 10310 27012 10362
rect 27064 10310 27076 10362
rect 27128 10310 27140 10362
rect 27192 10310 27204 10362
rect 27256 10310 30820 10362
rect 1104 10288 30820 10310
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 9858 10248 9864 10260
rect 7984 10220 9864 10248
rect 7984 10208 7990 10220
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 13170 10208 13176 10260
rect 13228 10208 13234 10260
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 9968 10112 9996 10208
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 8956 10084 9352 10112
rect 9968 10084 10149 10112
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 6270 10044 6276 10056
rect 5224 10016 6276 10044
rect 5224 10004 5230 10016
rect 6270 10004 6276 10016
rect 6328 10044 6334 10056
rect 8956 10053 8984 10084
rect 9324 10056 9352 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 13188 10112 13216 10208
rect 10137 10075 10195 10081
rect 12544 10084 13216 10112
rect 13464 10180 13492 10211
rect 13538 10208 13544 10260
rect 13596 10248 13602 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 13596 10220 13645 10248
rect 13596 10208 13602 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14323 10220 14657 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 15378 10248 15384 10260
rect 14645 10211 14703 10217
rect 14752 10220 15384 10248
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 13464 10152 14473 10180
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6328 10016 6469 10044
rect 6328 10004 6334 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9214 10044 9220 10056
rect 9171 10016 9220 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 6748 9920 6776 10007
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9306 10004 9312 10056
rect 9364 10004 9370 10056
rect 12544 10053 12572 10084
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13078 10044 13084 10056
rect 12851 10016 13084 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 9030 9936 9036 9988
rect 9088 9976 9094 9988
rect 10244 9976 10272 10007
rect 9088 9948 10272 9976
rect 9088 9936 9094 9948
rect 6730 9868 6736 9920
rect 6788 9868 6794 9920
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9908 7527 9911
rect 8570 9908 8576 9920
rect 7515 9880 8576 9908
rect 7515 9877 7527 9880
rect 7469 9871 7527 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 10594 9868 10600 9920
rect 10652 9868 10658 9920
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12636 9908 12664 10007
rect 12728 9976 12756 10007
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13173 10047 13231 10053
rect 13173 10013 13185 10047
rect 13219 10044 13231 10047
rect 13354 10044 13360 10056
rect 13219 10016 13360 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13464 9976 13492 10152
rect 14461 10149 14473 10152
rect 14507 10149 14519 10183
rect 14461 10143 14519 10149
rect 14752 10121 14780 10220
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17310 10248 17316 10260
rect 17267 10220 17316 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17420 10220 22232 10248
rect 17420 10180 17448 10220
rect 15856 10152 17448 10180
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 15059 10084 15485 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 15473 10081 15485 10084
rect 15519 10081 15531 10115
rect 15473 10075 15531 10081
rect 14182 10004 14188 10056
rect 14240 10004 14246 10056
rect 14826 10004 14832 10056
rect 14884 10004 14890 10056
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 15565 10047 15623 10053
rect 15565 10013 15577 10047
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 12728 9948 13492 9976
rect 14844 9976 14872 10004
rect 15580 9976 15608 10007
rect 14844 9948 15608 9976
rect 12584 9880 12664 9908
rect 12989 9911 13047 9917
rect 12584 9868 12590 9880
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 15856 9908 15884 10152
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 16850 10112 16856 10124
rect 16715 10084 16856 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17310 10072 17316 10124
rect 17368 10112 17374 10124
rect 19334 10112 19340 10124
rect 17368 10084 19340 10112
rect 17368 10072 17374 10084
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19444 10112 19472 10220
rect 20806 10180 20812 10192
rect 19720 10152 20812 10180
rect 19613 10115 19671 10121
rect 19613 10112 19625 10115
rect 19444 10084 19625 10112
rect 19613 10081 19625 10084
rect 19659 10081 19671 10115
rect 19613 10075 19671 10081
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 19518 10044 19524 10056
rect 19475 10016 19524 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 19518 10004 19524 10016
rect 19576 10004 19582 10056
rect 19720 10053 19748 10152
rect 20806 10140 20812 10152
rect 20864 10140 20870 10192
rect 20898 10140 20904 10192
rect 20956 10180 20962 10192
rect 20956 10152 22140 10180
rect 20956 10140 20962 10152
rect 20165 10115 20223 10121
rect 20165 10081 20177 10115
rect 20211 10112 20223 10115
rect 20530 10112 20536 10124
rect 20211 10084 20536 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 21453 10115 21511 10121
rect 21453 10112 21465 10115
rect 20732 10084 21465 10112
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 20441 10047 20499 10053
rect 20441 10044 20453 10047
rect 19705 10007 19763 10013
rect 19812 10016 20453 10044
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16540 9948 16896 9976
rect 16540 9936 16546 9948
rect 13035 9880 15884 9908
rect 15933 9911 15991 9917
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 15933 9877 15945 9911
rect 15979 9908 15991 9911
rect 16574 9908 16580 9920
rect 15979 9880 16580 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 16758 9868 16764 9920
rect 16816 9868 16822 9920
rect 16868 9917 16896 9948
rect 17494 9936 17500 9988
rect 17552 9976 17558 9988
rect 17589 9979 17647 9985
rect 17589 9976 17601 9979
rect 17552 9948 17601 9976
rect 17552 9936 17558 9948
rect 17589 9945 17601 9948
rect 17635 9945 17647 9979
rect 19337 9979 19395 9985
rect 19337 9976 19349 9979
rect 18814 9948 19349 9976
rect 17589 9939 17647 9945
rect 19337 9945 19349 9948
rect 19383 9945 19395 9979
rect 19812 9976 19840 10016
rect 20441 10013 20453 10016
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 20624 10047 20682 10053
rect 20624 10013 20636 10047
rect 20670 10046 20682 10047
rect 20732 10046 20760 10084
rect 21453 10081 21465 10084
rect 21499 10081 21511 10115
rect 22002 10112 22008 10124
rect 21453 10075 21511 10081
rect 21560 10084 22008 10112
rect 20670 10018 20760 10046
rect 20670 10013 20682 10018
rect 20624 10007 20682 10013
rect 21174 10004 21180 10056
rect 21232 10044 21238 10056
rect 21560 10053 21588 10084
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 21269 10047 21327 10053
rect 21269 10044 21281 10047
rect 21232 10016 21281 10044
rect 21232 10004 21238 10016
rect 21269 10013 21281 10016
rect 21315 10044 21327 10047
rect 21361 10047 21419 10053
rect 21361 10044 21373 10047
rect 21315 10016 21373 10044
rect 21315 10013 21327 10016
rect 21269 10007 21327 10013
rect 21361 10013 21373 10016
rect 21407 10013 21419 10047
rect 21361 10007 21419 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10013 21603 10047
rect 22112 10044 22140 10152
rect 22204 10112 22232 10220
rect 22278 10208 22284 10260
rect 22336 10248 22342 10260
rect 23014 10248 23020 10260
rect 22336 10220 23020 10248
rect 22336 10208 22342 10220
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 24949 10251 25007 10257
rect 24949 10217 24961 10251
rect 24995 10248 25007 10251
rect 25498 10248 25504 10260
rect 24995 10220 25504 10248
rect 24995 10217 25007 10220
rect 24949 10211 25007 10217
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 25958 10208 25964 10260
rect 26016 10208 26022 10260
rect 24762 10140 24768 10192
rect 24820 10140 24826 10192
rect 25774 10112 25780 10124
rect 22204 10084 25780 10112
rect 25774 10072 25780 10084
rect 25832 10072 25838 10124
rect 22370 10044 22376 10056
rect 22112 10016 22376 10044
rect 21545 10007 21603 10013
rect 20303 9979 20361 9985
rect 20303 9976 20315 9979
rect 19337 9939 19395 9945
rect 19444 9948 19840 9976
rect 20088 9948 20315 9976
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 18230 9908 18236 9920
rect 16899 9880 18236 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 18230 9868 18236 9880
rect 18288 9908 18294 9920
rect 19061 9911 19119 9917
rect 19061 9908 19073 9911
rect 18288 9880 19073 9908
rect 18288 9868 18294 9880
rect 19061 9877 19073 9880
rect 19107 9877 19119 9911
rect 19061 9871 19119 9877
rect 19150 9868 19156 9920
rect 19208 9908 19214 9920
rect 19444 9908 19472 9948
rect 20088 9917 20116 9948
rect 20303 9945 20315 9948
rect 20349 9945 20361 9979
rect 20303 9939 20361 9945
rect 20533 9979 20591 9985
rect 20533 9945 20545 9979
rect 20579 9976 20591 9979
rect 20898 9976 20904 9988
rect 20579 9948 20904 9976
rect 20579 9945 20591 9948
rect 20533 9939 20591 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21085 9979 21143 9985
rect 21085 9945 21097 9979
rect 21131 9945 21143 9979
rect 21085 9939 21143 9945
rect 19208 9880 19472 9908
rect 20073 9911 20131 9917
rect 19208 9868 19214 9880
rect 20073 9877 20085 9911
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 20622 9868 20628 9920
rect 20680 9908 20686 9920
rect 20809 9911 20867 9917
rect 20809 9908 20821 9911
rect 20680 9880 20821 9908
rect 20680 9868 20686 9880
rect 20809 9877 20821 9880
rect 20855 9877 20867 9911
rect 21100 9908 21128 9939
rect 21560 9908 21588 10007
rect 22370 10004 22376 10016
rect 22428 10044 22434 10056
rect 22554 10044 22560 10056
rect 22428 10016 22560 10044
rect 22428 10004 22434 10016
rect 22554 10004 22560 10016
rect 22612 10004 22618 10056
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10044 22799 10047
rect 22787 10016 23060 10044
rect 22787 10013 22799 10016
rect 22741 10007 22799 10013
rect 23032 9920 23060 10016
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 24912 10016 25697 10044
rect 24912 10004 24918 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 25961 10047 26019 10053
rect 25961 10013 25973 10047
rect 26007 10013 26019 10047
rect 25961 10007 26019 10013
rect 24489 9979 24547 9985
rect 24489 9945 24501 9979
rect 24535 9976 24547 9979
rect 24578 9976 24584 9988
rect 24535 9948 24584 9976
rect 24535 9945 24547 9948
rect 24489 9939 24547 9945
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 25406 9936 25412 9988
rect 25464 9976 25470 9988
rect 25869 9979 25927 9985
rect 25869 9976 25881 9979
rect 25464 9948 25881 9976
rect 25464 9936 25470 9948
rect 25869 9945 25881 9948
rect 25915 9945 25927 9979
rect 25869 9939 25927 9945
rect 25976 9920 26004 10007
rect 21100 9880 21588 9908
rect 20809 9871 20867 9877
rect 22646 9868 22652 9920
rect 22704 9868 22710 9920
rect 23014 9868 23020 9920
rect 23072 9868 23078 9920
rect 25958 9868 25964 9920
rect 26016 9868 26022 9920
rect 1104 9818 30820 9840
rect 1104 9766 5324 9818
rect 5376 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 12752 9818
rect 12804 9766 12816 9818
rect 12868 9766 12880 9818
rect 12932 9766 12944 9818
rect 12996 9766 13008 9818
rect 13060 9766 20180 9818
rect 20232 9766 20244 9818
rect 20296 9766 20308 9818
rect 20360 9766 20372 9818
rect 20424 9766 20436 9818
rect 20488 9766 27608 9818
rect 27660 9766 27672 9818
rect 27724 9766 27736 9818
rect 27788 9766 27800 9818
rect 27852 9766 27864 9818
rect 27916 9766 30820 9818
rect 1104 9744 30820 9766
rect 8757 9707 8815 9713
rect 5828 9676 6684 9704
rect 3602 9596 3608 9648
rect 3660 9596 3666 9648
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 5828 9636 5856 9676
rect 4120 9608 5856 9636
rect 5905 9639 5963 9645
rect 4120 9596 4126 9608
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 5951 9608 6561 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 6656 9636 6684 9676
rect 8757 9673 8769 9707
rect 8803 9704 8815 9707
rect 9306 9704 9312 9716
rect 8803 9676 9312 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 12618 9664 12624 9716
rect 12676 9664 12682 9716
rect 13262 9704 13268 9716
rect 12728 9676 13268 9704
rect 6730 9636 6736 9648
rect 6656 9608 6736 9636
rect 6549 9599 6607 9605
rect 6730 9596 6736 9608
rect 6788 9636 6794 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 6788 9608 8217 9636
rect 6788 9596 6794 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 12342 9636 12348 9648
rect 8205 9599 8263 9605
rect 10796 9608 12348 9636
rect 10796 9580 10824 9608
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4080 9540 4537 9568
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 2332 9364 2360 9463
rect 2590 9460 2596 9512
rect 2648 9460 2654 9512
rect 4080 9509 4108 9540
rect 4525 9537 4537 9540
rect 4571 9568 4583 9571
rect 4571 9540 5120 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 5092 9500 5120 9540
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 5408 9540 5457 9568
rect 5408 9528 5414 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5592 9540 5641 9568
rect 5592 9528 5598 9540
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5736 9540 6408 9568
rect 5736 9500 5764 9540
rect 5092 9472 5764 9500
rect 4801 9463 4859 9469
rect 3326 9364 3332 9376
rect 2332 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4154 9324 4160 9376
rect 4212 9324 4218 9376
rect 4632 9364 4660 9463
rect 4816 9432 4844 9463
rect 6178 9460 6184 9512
rect 6236 9460 6242 9512
rect 6380 9509 6408 9540
rect 8570 9528 8576 9580
rect 8628 9568 8634 9580
rect 9306 9568 9312 9580
rect 8628 9540 9312 9568
rect 8628 9528 8634 9540
rect 9306 9528 9312 9540
rect 9364 9568 9370 9580
rect 9674 9577 9680 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9364 9540 9505 9568
rect 9364 9528 9370 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9670 9568 9680 9577
rect 9635 9540 9680 9568
rect 9493 9531 9551 9537
rect 9670 9531 9680 9540
rect 9674 9528 9680 9531
rect 9732 9528 9738 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11514 9528 11520 9580
rect 11572 9528 11578 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12492 9540 12541 9568
rect 12492 9528 12498 9540
rect 12529 9537 12541 9540
rect 12575 9568 12587 9571
rect 12728 9568 12756 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 16945 9707 17003 9713
rect 16945 9704 16957 9707
rect 16816 9676 16957 9704
rect 16816 9664 16822 9676
rect 16945 9673 16957 9676
rect 16991 9673 17003 9707
rect 19150 9704 19156 9716
rect 16945 9667 17003 9673
rect 17880 9676 19156 9704
rect 12820 9608 14228 9636
rect 12820 9577 12848 9608
rect 14200 9580 14228 9608
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17431 9639 17489 9645
rect 17431 9636 17443 9639
rect 16632 9608 17443 9636
rect 16632 9596 16638 9608
rect 17431 9605 17443 9608
rect 17477 9605 17489 9639
rect 17431 9599 17489 9605
rect 12575 9540 12756 9568
rect 12805 9571 12863 9577
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12805 9537 12817 9571
rect 12851 9537 12863 9571
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12805 9531 12863 9537
rect 13004 9540 13185 9568
rect 6365 9503 6423 9509
rect 6365 9469 6377 9503
rect 6411 9500 6423 9503
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 6411 9472 8309 9500
rect 6411 9469 6423 9472
rect 6365 9463 6423 9469
rect 8297 9469 8309 9472
rect 8343 9500 8355 9503
rect 8849 9503 8907 9509
rect 8343 9472 8708 9500
rect 8343 9469 8355 9472
rect 8297 9463 8355 9469
rect 5166 9432 5172 9444
rect 4816 9404 5172 9432
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 8570 9392 8576 9444
rect 8628 9392 8634 9444
rect 8680 9432 8708 9472
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 9214 9500 9220 9512
rect 8895 9472 9220 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9631 9472 9965 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 9953 9469 9965 9472
rect 9999 9469 10011 9503
rect 9953 9463 10011 9469
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 10689 9503 10747 9509
rect 10689 9500 10701 9503
rect 10275 9472 10701 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 10689 9469 10701 9472
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 8941 9435 8999 9441
rect 8941 9432 8953 9435
rect 8680 9404 8953 9432
rect 8941 9401 8953 9404
rect 8987 9401 8999 9435
rect 8941 9395 8999 9401
rect 9490 9392 9496 9444
rect 9548 9432 9554 9444
rect 10060 9432 10088 9463
rect 9548 9404 10088 9432
rect 10152 9432 10180 9463
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 11256 9432 11284 9460
rect 10152 9404 11284 9432
rect 12253 9435 12311 9441
rect 9548 9392 9554 9404
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12710 9432 12716 9444
rect 12299 9404 12716 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 4632 9336 9781 9364
rect 9769 9333 9781 9336
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 13004 9373 13032 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13354 9528 13360 9580
rect 13412 9528 13418 9580
rect 14182 9528 14188 9580
rect 14240 9528 14246 9580
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 15838 9568 15844 9580
rect 15068 9540 15844 9568
rect 15068 9528 15074 9540
rect 15838 9528 15844 9540
rect 15896 9568 15902 9580
rect 16850 9568 16856 9580
rect 15896 9540 16856 9568
rect 15896 9528 15902 9540
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17126 9528 17132 9580
rect 17184 9528 17190 9580
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9537 17279 9571
rect 17221 9531 17279 9537
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9500 13139 9503
rect 13372 9500 13400 9528
rect 13127 9472 13400 9500
rect 13127 9469 13139 9472
rect 13081 9463 13139 9469
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16942 9500 16948 9512
rect 16080 9472 16948 9500
rect 16080 9460 16086 9472
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17236 9500 17264 9531
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 17880 9568 17908 9676
rect 19150 9664 19156 9676
rect 19208 9704 19214 9716
rect 22554 9704 22560 9716
rect 19208 9676 22560 9704
rect 19208 9664 19214 9676
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 22646 9664 22652 9716
rect 22704 9664 22710 9716
rect 22465 9639 22523 9645
rect 22465 9605 22477 9639
rect 22511 9636 22523 9639
rect 22572 9636 22600 9664
rect 22511 9608 22600 9636
rect 22511 9605 22523 9608
rect 22465 9599 22523 9605
rect 17368 9540 17908 9568
rect 17368 9528 17374 9540
rect 18138 9528 18144 9580
rect 18196 9528 18202 9580
rect 22664 9577 22692 9664
rect 22830 9596 22836 9648
rect 22888 9596 22894 9648
rect 23474 9596 23480 9648
rect 23532 9636 23538 9648
rect 23845 9639 23903 9645
rect 23845 9636 23857 9639
rect 23532 9608 23857 9636
rect 23532 9596 23538 9608
rect 23845 9605 23857 9608
rect 23891 9605 23903 9639
rect 23845 9599 23903 9605
rect 23937 9639 23995 9645
rect 23937 9605 23949 9639
rect 23983 9636 23995 9639
rect 24762 9636 24768 9648
rect 23983 9608 24768 9636
rect 23983 9605 23995 9608
rect 23937 9599 23995 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 24946 9596 24952 9648
rect 25004 9636 25010 9648
rect 25004 9608 25452 9636
rect 25004 9596 25010 9608
rect 22327 9571 22385 9577
rect 22327 9568 22339 9571
rect 22112 9540 22339 9568
rect 17402 9500 17408 9512
rect 17236 9472 17408 9500
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9500 17647 9503
rect 18156 9500 18184 9528
rect 17635 9472 18184 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 16390 9392 16396 9444
rect 16448 9432 16454 9444
rect 17604 9432 17632 9463
rect 16448 9404 17632 9432
rect 16448 9392 16454 9404
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12676 9336 13001 9364
rect 12676 9324 12682 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 12989 9327 13047 9333
rect 13170 9324 13176 9376
rect 13228 9324 13234 9376
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 18230 9364 18236 9376
rect 16816 9336 18236 9364
rect 16816 9324 16822 9336
rect 18230 9324 18236 9336
rect 18288 9364 18294 9376
rect 19518 9364 19524 9376
rect 18288 9336 19524 9364
rect 18288 9324 18294 9336
rect 19518 9324 19524 9336
rect 19576 9364 19582 9376
rect 20530 9364 20536 9376
rect 19576 9336 20536 9364
rect 19576 9324 19582 9336
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 22112 9364 22140 9540
rect 22327 9537 22339 9540
rect 22373 9537 22385 9571
rect 22327 9531 22385 9537
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 22189 9503 22247 9509
rect 22189 9469 22201 9503
rect 22235 9500 22247 9503
rect 22572 9500 22600 9531
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 22796 9540 23121 9568
rect 22796 9528 22802 9540
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23707 9571 23765 9577
rect 23707 9568 23719 9571
rect 23109 9531 23167 9537
rect 23492 9540 23719 9568
rect 22922 9500 22928 9512
rect 22235 9472 22508 9500
rect 22572 9472 22928 9500
rect 22235 9469 22247 9472
rect 22189 9463 22247 9469
rect 22480 9444 22508 9472
rect 22922 9460 22928 9472
rect 22980 9500 22986 9512
rect 23492 9509 23520 9540
rect 23707 9537 23719 9540
rect 23753 9537 23765 9571
rect 23707 9531 23765 9537
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9568 24087 9571
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24075 9540 24869 9568
rect 24075 9537 24087 9540
rect 24029 9531 24087 9537
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 24857 9531 24915 9537
rect 25038 9528 25044 9580
rect 25096 9528 25102 9580
rect 25133 9571 25191 9577
rect 25133 9537 25145 9571
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 23017 9503 23075 9509
rect 23017 9500 23029 9503
rect 22980 9472 23029 9500
rect 22980 9460 22986 9472
rect 23017 9469 23029 9472
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 23477 9503 23535 9509
rect 23477 9469 23489 9503
rect 23523 9469 23535 9503
rect 23477 9463 23535 9469
rect 23569 9503 23627 9509
rect 23569 9469 23581 9503
rect 23615 9469 23627 9503
rect 25148 9500 25176 9531
rect 25314 9528 25320 9580
rect 25372 9528 25378 9580
rect 25424 9577 25452 9608
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9568 25467 9571
rect 25682 9568 25688 9580
rect 25455 9540 25688 9568
rect 25455 9537 25467 9540
rect 25409 9531 25467 9537
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 26016 9540 26065 9568
rect 26016 9528 26022 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 25976 9500 26004 9528
rect 25148 9472 26004 9500
rect 23569 9463 23627 9469
rect 22462 9392 22468 9444
rect 22520 9392 22526 9444
rect 22554 9392 22560 9444
rect 22612 9432 22618 9444
rect 23584 9432 23612 9463
rect 26142 9460 26148 9512
rect 26200 9460 26206 9512
rect 25685 9435 25743 9441
rect 25685 9432 25697 9435
rect 22612 9404 23612 9432
rect 24044 9404 25697 9432
rect 22612 9392 22618 9404
rect 24044 9364 24072 9404
rect 25685 9401 25697 9404
rect 25731 9401 25743 9435
rect 25685 9395 25743 9401
rect 22112 9336 24072 9364
rect 24210 9324 24216 9376
rect 24268 9324 24274 9376
rect 1104 9274 30820 9296
rect 1104 9222 4664 9274
rect 4716 9222 4728 9274
rect 4780 9222 4792 9274
rect 4844 9222 4856 9274
rect 4908 9222 4920 9274
rect 4972 9222 12092 9274
rect 12144 9222 12156 9274
rect 12208 9222 12220 9274
rect 12272 9222 12284 9274
rect 12336 9222 12348 9274
rect 12400 9222 19520 9274
rect 19572 9222 19584 9274
rect 19636 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 26948 9274
rect 27000 9222 27012 9274
rect 27064 9222 27076 9274
rect 27128 9222 27140 9274
rect 27192 9222 27204 9274
rect 27256 9222 30820 9274
rect 1104 9200 30820 9222
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 2869 9163 2927 9169
rect 2869 9160 2881 9163
rect 2648 9132 2881 9160
rect 2648 9120 2654 9132
rect 2869 9129 2881 9132
rect 2915 9129 2927 9163
rect 2869 9123 2927 9129
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 3602 9160 3608 9172
rect 3467 9132 3608 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4154 9120 4160 9172
rect 4212 9120 4218 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4890 9160 4896 9172
rect 4396 9132 4896 9160
rect 4396 9120 4402 9132
rect 4890 9120 4896 9132
rect 4948 9160 4954 9172
rect 5166 9160 5172 9172
rect 4948 9132 5172 9160
rect 4948 9120 4954 9132
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9769 9163 9827 9169
rect 9769 9160 9781 9163
rect 9548 9132 9781 9160
rect 9548 9120 9554 9132
rect 9769 9129 9781 9132
rect 9815 9129 9827 9163
rect 9769 9123 9827 9129
rect 12618 9120 12624 9172
rect 12676 9120 12682 9172
rect 13170 9120 13176 9172
rect 13228 9120 13234 9172
rect 14550 9120 14556 9172
rect 14608 9120 14614 9172
rect 14737 9163 14795 9169
rect 14737 9129 14749 9163
rect 14783 9160 14795 9163
rect 14918 9160 14924 9172
rect 14783 9132 14924 9160
rect 14783 9129 14795 9132
rect 14737 9123 14795 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 22922 9120 22928 9172
rect 22980 9120 22986 9172
rect 25038 9120 25044 9172
rect 25096 9160 25102 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 25096 9132 25329 9160
rect 25096 9120 25102 9132
rect 25317 9129 25329 9132
rect 25363 9160 25375 9163
rect 25363 9132 26096 9160
rect 25363 9129 25375 9132
rect 25317 9123 25375 9129
rect 4172 9024 4200 9120
rect 12434 9092 12440 9104
rect 7944 9064 12440 9092
rect 5350 9024 5356 9036
rect 3068 8996 4200 9024
rect 4540 8996 5356 9024
rect 3068 8965 3096 8996
rect 4540 8968 4568 8996
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8956 3387 8959
rect 3418 8956 3424 8968
rect 3375 8928 3424 8956
rect 3375 8925 3387 8928
rect 3329 8919 3387 8925
rect 3418 8916 3424 8928
rect 3476 8956 3482 8968
rect 3476 8928 4016 8956
rect 3476 8916 3482 8928
rect 3988 8900 4016 8928
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 4816 8965 4844 8996
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 6178 9024 6184 9036
rect 5583 8996 6184 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 6178 8984 6184 8996
rect 6236 9024 6242 9036
rect 7944 9033 7972 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 13078 9092 13084 9104
rect 12544 9064 13084 9092
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 6236 8996 7941 9024
rect 6236 8984 6242 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 11330 9024 11336 9036
rect 8352 8996 11336 9024
rect 8352 8984 8358 8996
rect 11330 8984 11336 8996
rect 11388 9024 11394 9036
rect 12544 9024 12572 9064
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 11388 8996 12572 9024
rect 11388 8984 11394 8996
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 3970 8848 3976 8900
rect 4028 8848 4034 8900
rect 4632 8888 4660 8919
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 5132 8928 6929 8956
rect 5132 8916 5138 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 5092 8888 5120 8916
rect 4632 8860 5120 8888
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5261 8891 5319 8897
rect 5261 8888 5273 8891
rect 5224 8860 5273 8888
rect 5224 8848 5230 8860
rect 5261 8857 5273 8860
rect 5307 8857 5319 8891
rect 5261 8851 5319 8857
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 7208 8888 7236 8919
rect 5408 8860 7236 8888
rect 5408 8848 5414 8860
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5442 8820 5448 8832
rect 5040 8792 5448 8820
rect 5040 8780 5046 8792
rect 5442 8780 5448 8792
rect 5500 8820 5506 8832
rect 7392 8820 7420 8919
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9674 8956 9680 8968
rect 9447 8928 9680 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 12443 8959 12501 8965
rect 12443 8925 12455 8959
rect 12489 8956 12501 8959
rect 12544 8956 12572 8996
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 9024 13047 9027
rect 13188 9024 13216 9120
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 15470 9092 15476 9104
rect 13311 9064 15476 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 15470 9052 15476 9064
rect 15528 9052 15534 9104
rect 25406 9092 25412 9104
rect 20916 9064 25412 9092
rect 13035 8996 13216 9024
rect 13035 8993 13047 8996
rect 12989 8987 13047 8993
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 20916 9033 20944 9064
rect 25406 9052 25412 9064
rect 25464 9052 25470 9104
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20864 8996 20913 9024
rect 20864 8984 20870 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 9024 21879 9027
rect 22002 9024 22008 9036
rect 21867 8996 22008 9024
rect 21867 8993 21879 8996
rect 21821 8987 21879 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 26068 9024 26096 9132
rect 26142 9120 26148 9172
rect 26200 9160 26206 9172
rect 26237 9163 26295 9169
rect 26237 9160 26249 9163
rect 26200 9132 26249 9160
rect 26200 9120 26206 9132
rect 26237 9129 26249 9132
rect 26283 9129 26295 9163
rect 26237 9123 26295 9129
rect 26068 8996 26372 9024
rect 12489 8928 12572 8956
rect 12621 8959 12679 8965
rect 12489 8925 12501 8928
rect 12443 8919 12501 8925
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 12710 8956 12716 8968
rect 12667 8928 12716 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 14182 8956 14188 8968
rect 12943 8928 14188 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14366 8956 14372 8968
rect 14323 8928 14372 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15194 8916 15200 8968
rect 15252 8916 15258 8968
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18233 8959 18291 8965
rect 18003 8928 18184 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 7650 8848 7656 8900
rect 7708 8848 7714 8900
rect 9324 8888 9352 8916
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 9324 8860 9597 8888
rect 9585 8857 9597 8860
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 16758 8888 16764 8900
rect 11940 8860 16764 8888
rect 11940 8848 11946 8860
rect 16758 8848 16764 8860
rect 16816 8848 16822 8900
rect 18156 8832 18184 8928
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18414 8956 18420 8968
rect 18279 8928 18420 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18414 8916 18420 8928
rect 18472 8916 18478 8968
rect 21726 8916 21732 8968
rect 21784 8916 21790 8968
rect 22370 8916 22376 8968
rect 22428 8956 22434 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 22428 8928 22569 8956
rect 22428 8916 22434 8928
rect 22557 8925 22569 8928
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 25774 8916 25780 8968
rect 25832 8916 25838 8968
rect 26344 8965 26372 8996
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8925 26019 8959
rect 25961 8919 26019 8925
rect 26053 8959 26111 8965
rect 26053 8925 26065 8959
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26329 8959 26387 8965
rect 26329 8925 26341 8959
rect 26375 8925 26387 8959
rect 26329 8919 26387 8925
rect 22741 8891 22799 8897
rect 22741 8857 22753 8891
rect 22787 8888 22799 8891
rect 22922 8888 22928 8900
rect 22787 8860 22928 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 22922 8848 22928 8860
rect 22980 8848 22986 8900
rect 25866 8848 25872 8900
rect 25924 8888 25930 8900
rect 25976 8888 26004 8919
rect 25924 8860 26004 8888
rect 25924 8848 25930 8860
rect 5500 8792 7420 8820
rect 5500 8780 5506 8792
rect 7558 8780 7564 8832
rect 7616 8820 7622 8832
rect 10502 8820 10508 8832
rect 7616 8792 10508 8820
rect 7616 8780 7622 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 12710 8820 12716 8832
rect 12584 8792 12716 8820
rect 12584 8780 12590 8792
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 15378 8780 15384 8832
rect 15436 8780 15442 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 17221 8823 17279 8829
rect 17221 8820 17233 8823
rect 16632 8792 17233 8820
rect 16632 8780 16638 8792
rect 17221 8789 17233 8792
rect 17267 8789 17279 8823
rect 17221 8783 17279 8789
rect 18138 8780 18144 8832
rect 18196 8780 18202 8832
rect 25130 8780 25136 8832
rect 25188 8820 25194 8832
rect 26068 8820 26096 8919
rect 26421 8823 26479 8829
rect 26421 8820 26433 8823
rect 25188 8792 26433 8820
rect 25188 8780 25194 8792
rect 26421 8789 26433 8792
rect 26467 8789 26479 8823
rect 26421 8783 26479 8789
rect 1104 8730 30820 8752
rect 1104 8678 5324 8730
rect 5376 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 12752 8730
rect 12804 8678 12816 8730
rect 12868 8678 12880 8730
rect 12932 8678 12944 8730
rect 12996 8678 13008 8730
rect 13060 8678 20180 8730
rect 20232 8678 20244 8730
rect 20296 8678 20308 8730
rect 20360 8678 20372 8730
rect 20424 8678 20436 8730
rect 20488 8678 27608 8730
rect 27660 8678 27672 8730
rect 27724 8678 27736 8730
rect 27788 8678 27800 8730
rect 27852 8678 27864 8730
rect 27916 8678 30820 8730
rect 1104 8656 30820 8678
rect 8294 8576 8300 8628
rect 8352 8576 8358 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 8430 8588 10333 8616
rect 8312 8548 8340 8576
rect 7852 8520 8340 8548
rect 8430 8557 8458 8588
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 10778 8576 10784 8628
rect 10836 8576 10842 8628
rect 12526 8576 12532 8628
rect 12584 8576 12590 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 14182 8616 14188 8628
rect 13587 8588 14188 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14921 8619 14979 8625
rect 14921 8585 14933 8619
rect 14967 8616 14979 8619
rect 15194 8616 15200 8628
rect 14967 8588 15200 8616
rect 14967 8585 14979 8588
rect 14921 8579 14979 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15335 8588 17172 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 8430 8551 8493 8557
rect 8430 8520 8447 8551
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7190 8480 7196 8492
rect 6687 8452 7196 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7852 8489 7880 8520
rect 8435 8517 8447 8520
rect 8481 8517 8493 8551
rect 8754 8548 8760 8560
rect 8435 8511 8493 8517
rect 8588 8520 8760 8548
rect 7653 8483 7711 8489
rect 7653 8480 7665 8483
rect 7616 8452 7665 8480
rect 7616 8440 7622 8452
rect 7653 8449 7665 8452
rect 7699 8449 7711 8483
rect 7653 8443 7711 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8110 8440 8116 8492
rect 8168 8440 8174 8492
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8588 8480 8616 8520
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 9490 8548 9496 8560
rect 8864 8520 9496 8548
rect 8864 8489 8892 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 9674 8508 9680 8560
rect 9732 8508 9738 8560
rect 10796 8548 10824 8576
rect 10428 8520 10824 8548
rect 8343 8452 8616 8480
rect 8673 8483 8731 8489
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8673 8449 8685 8483
rect 8719 8480 8731 8483
rect 8849 8483 8907 8489
rect 8719 8452 8800 8480
rect 8719 8449 8731 8452
rect 8673 8443 8731 8449
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 7791 8384 8064 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 7929 8347 7987 8353
rect 7929 8344 7941 8347
rect 6420 8316 7604 8344
rect 6420 8304 6426 8316
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 7101 8279 7159 8285
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7374 8276 7380 8288
rect 7147 8248 7380 8276
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 7576 8276 7604 8316
rect 7760 8316 7941 8344
rect 7760 8276 7788 8316
rect 7929 8313 7941 8316
rect 7975 8313 7987 8347
rect 7929 8307 7987 8313
rect 7576 8248 7788 8276
rect 8036 8276 8064 8384
rect 8404 8384 8585 8412
rect 8404 8276 8432 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8772 8412 8800 8452
rect 8849 8449 8861 8483
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9214 8480 9220 8492
rect 9171 8452 9220 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9692 8480 9720 8508
rect 10428 8489 10456 8520
rect 9447 8452 9720 8480
rect 10229 8483 10287 8489
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 8772 8384 9168 8412
rect 8573 8375 8631 8381
rect 8754 8304 8760 8356
rect 8812 8304 8818 8356
rect 9140 8288 9168 8384
rect 9306 8372 9312 8424
rect 9364 8372 9370 8424
rect 10244 8412 10272 8443
rect 10502 8440 10508 8492
rect 10560 8480 10566 8492
rect 10689 8483 10747 8489
rect 10560 8452 10640 8480
rect 10560 8440 10566 8452
rect 10612 8412 10640 8452
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 10962 8480 10968 8492
rect 10735 8452 10968 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 10962 8440 10968 8452
rect 11020 8480 11026 8492
rect 11330 8480 11336 8492
rect 11020 8452 11336 8480
rect 11020 8440 11026 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 12434 8440 12440 8492
rect 12492 8440 12498 8492
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8480 12679 8483
rect 13630 8480 13636 8492
rect 12667 8452 13636 8480
rect 12667 8449 12679 8452
rect 12621 8443 12679 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15304 8480 15332 8579
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 16235 8551 16293 8557
rect 16235 8548 16247 8551
rect 15528 8520 16247 8548
rect 15528 8508 15534 8520
rect 16235 8517 16247 8520
rect 16281 8517 16293 8551
rect 16235 8511 16293 8517
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 16816 8520 16896 8548
rect 16816 8508 16822 8520
rect 14424 8452 15332 8480
rect 15381 8483 15439 8489
rect 14424 8440 14430 8452
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15427 8452 15761 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15930 8440 15936 8492
rect 15988 8440 15994 8492
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 10870 8412 10876 8424
rect 10244 8384 10548 8412
rect 10612 8384 10876 8412
rect 10520 8353 10548 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8412 14519 8415
rect 14550 8412 14556 8424
rect 14507 8384 14556 8412
rect 14507 8381 14519 8384
rect 14461 8375 14519 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 15838 8412 15844 8424
rect 15611 8384 15844 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 15838 8372 15844 8384
rect 15896 8372 15902 8424
rect 16132 8412 16160 8443
rect 16390 8440 16396 8492
rect 16448 8440 16454 8492
rect 16868 8489 16896 8520
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17144 8424 17172 8588
rect 21726 8576 21732 8628
rect 21784 8576 21790 8628
rect 22281 8619 22339 8625
rect 22281 8585 22293 8619
rect 22327 8585 22339 8619
rect 22281 8579 22339 8585
rect 17313 8551 17371 8557
rect 17313 8517 17325 8551
rect 17359 8548 17371 8551
rect 17954 8548 17960 8560
rect 17359 8520 17960 8548
rect 17359 8517 17371 8520
rect 17313 8511 17371 8517
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 20530 8548 20536 8560
rect 19720 8520 20536 8548
rect 19720 8489 19748 8520
rect 20530 8508 20536 8520
rect 20588 8548 20594 8560
rect 21744 8548 21772 8576
rect 20588 8520 21772 8548
rect 22296 8548 22324 8579
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 23382 8616 23388 8628
rect 22796 8588 23388 8616
rect 22796 8576 22802 8588
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 24578 8576 24584 8628
rect 24636 8576 24642 8628
rect 24762 8576 24768 8628
rect 24820 8616 24826 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24820 8588 24961 8616
rect 24820 8576 24826 8588
rect 24949 8585 24961 8588
rect 24995 8585 25007 8619
rect 25590 8616 25596 8628
rect 24949 8579 25007 8585
rect 25332 8588 25596 8616
rect 25332 8557 25360 8588
rect 25590 8576 25596 8588
rect 25648 8616 25654 8628
rect 25869 8619 25927 8625
rect 25869 8616 25881 8619
rect 25648 8588 25881 8616
rect 25648 8576 25654 8588
rect 25869 8585 25881 8588
rect 25915 8585 25927 8619
rect 25869 8579 25927 8585
rect 25225 8551 25283 8557
rect 25225 8548 25237 8551
rect 22296 8520 25237 8548
rect 20588 8508 20594 8520
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8449 19763 8483
rect 21744 8480 21772 8520
rect 25225 8517 25237 8520
rect 25271 8517 25283 8551
rect 25225 8511 25283 8517
rect 25317 8551 25375 8557
rect 25317 8517 25329 8551
rect 25363 8517 25375 8551
rect 25685 8551 25743 8557
rect 25685 8548 25697 8551
rect 25317 8511 25375 8517
rect 25516 8520 25697 8548
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21744 8452 21833 8480
rect 19705 8443 19763 8449
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22646 8440 22652 8492
rect 22704 8440 22710 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 23707 8452 24532 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 16040 8384 16160 8412
rect 10505 8347 10563 8353
rect 10505 8313 10517 8347
rect 10551 8344 10563 8347
rect 10594 8344 10600 8356
rect 10551 8316 10600 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 11238 8304 11244 8356
rect 11296 8344 11302 8356
rect 16040 8344 16068 8384
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 18138 8372 18144 8424
rect 18196 8372 18202 8424
rect 19886 8372 19892 8424
rect 19944 8372 19950 8424
rect 20806 8372 20812 8424
rect 20864 8372 20870 8424
rect 22370 8372 22376 8424
rect 22428 8372 22434 8424
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23569 8415 23627 8421
rect 23569 8412 23581 8415
rect 23440 8384 23581 8412
rect 23440 8372 23446 8384
rect 23569 8381 23581 8384
rect 23615 8412 23627 8415
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23615 8384 24133 8412
rect 23615 8381 23627 8384
rect 23569 8375 23627 8381
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 17310 8344 17316 8356
rect 11296 8316 17316 8344
rect 11296 8304 11302 8316
rect 17310 8304 17316 8316
rect 17368 8304 17374 8356
rect 18414 8304 18420 8356
rect 18472 8344 18478 8356
rect 24504 8353 24532 8452
rect 25130 8440 25136 8492
rect 25188 8440 25194 8492
rect 25240 8412 25268 8511
rect 25406 8440 25412 8492
rect 25464 8480 25470 8492
rect 25516 8489 25544 8520
rect 25685 8517 25697 8520
rect 25731 8517 25743 8551
rect 26145 8551 26203 8557
rect 26145 8548 26157 8551
rect 25685 8511 25743 8517
rect 25792 8520 26157 8548
rect 25501 8483 25559 8489
rect 25501 8480 25513 8483
rect 25464 8452 25513 8480
rect 25464 8440 25470 8452
rect 25501 8449 25513 8452
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8478 25651 8483
rect 25792 8478 25820 8520
rect 26145 8517 26157 8520
rect 26191 8517 26203 8551
rect 26145 8511 26203 8517
rect 25639 8450 25820 8478
rect 25639 8449 25651 8450
rect 25593 8443 25651 8449
rect 25866 8440 25872 8492
rect 25924 8480 25930 8492
rect 25961 8483 26019 8489
rect 25961 8480 25973 8483
rect 25924 8452 25973 8480
rect 25924 8440 25930 8452
rect 25961 8449 25973 8452
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 26053 8483 26111 8489
rect 26053 8449 26065 8483
rect 26099 8480 26111 8483
rect 26099 8452 26280 8480
rect 26099 8449 26111 8452
rect 26053 8443 26111 8449
rect 25976 8412 26004 8443
rect 25240 8384 26004 8412
rect 24029 8347 24087 8353
rect 18472 8316 19380 8344
rect 18472 8304 18478 8316
rect 8036 8248 8432 8276
rect 8938 8236 8944 8288
rect 8996 8236 9002 8288
rect 9122 8236 9128 8288
rect 9180 8236 9186 8288
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9398 8276 9404 8288
rect 9272 8248 9404 8276
rect 9272 8236 9278 8248
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 16574 8276 16580 8288
rect 14608 8248 16580 8276
rect 14608 8236 14614 8248
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 16758 8236 16764 8288
rect 16816 8236 16822 8288
rect 19352 8276 19380 8316
rect 24029 8313 24041 8347
rect 24075 8344 24087 8347
rect 24489 8347 24547 8353
rect 24075 8316 24440 8344
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 19794 8276 19800 8288
rect 19352 8248 19800 8276
rect 19794 8236 19800 8248
rect 19852 8276 19858 8288
rect 20254 8276 20260 8288
rect 19852 8248 20260 8276
rect 19852 8236 19858 8248
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 22002 8236 22008 8288
rect 22060 8236 22066 8288
rect 24412 8276 24440 8316
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 24670 8344 24676 8356
rect 24535 8316 24676 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 25682 8304 25688 8356
rect 25740 8304 25746 8356
rect 26252 8344 26280 8452
rect 25792 8316 26280 8344
rect 25314 8276 25320 8288
rect 24412 8248 25320 8276
rect 25314 8236 25320 8248
rect 25372 8276 25378 8288
rect 25792 8276 25820 8316
rect 25372 8248 25820 8276
rect 25372 8236 25378 8248
rect 1104 8186 30820 8208
rect 1104 8134 4664 8186
rect 4716 8134 4728 8186
rect 4780 8134 4792 8186
rect 4844 8134 4856 8186
rect 4908 8134 4920 8186
rect 4972 8134 12092 8186
rect 12144 8134 12156 8186
rect 12208 8134 12220 8186
rect 12272 8134 12284 8186
rect 12336 8134 12348 8186
rect 12400 8134 19520 8186
rect 19572 8134 19584 8186
rect 19636 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 26948 8186
rect 27000 8134 27012 8186
rect 27064 8134 27076 8186
rect 27128 8134 27140 8186
rect 27192 8134 27204 8186
rect 27256 8134 30820 8186
rect 1104 8112 30820 8134
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7616 8044 7757 8072
rect 7616 8032 7622 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 8846 8072 8852 8084
rect 8260 8044 8852 8072
rect 8260 8032 8266 8044
rect 8846 8032 8852 8044
rect 8904 8072 8910 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8904 8044 8953 8072
rect 8904 8032 8910 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 10686 8072 10692 8084
rect 9456 8044 10692 8072
rect 9456 8032 9462 8044
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 12434 8072 12440 8084
rect 11287 8044 12440 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 15286 8032 15292 8084
rect 15344 8072 15350 8084
rect 16022 8072 16028 8084
rect 15344 8044 16028 8072
rect 15344 8032 15350 8044
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 17126 8032 17132 8084
rect 17184 8032 17190 8084
rect 17954 8032 17960 8084
rect 18012 8032 18018 8084
rect 18782 8072 18788 8084
rect 18064 8044 18788 8072
rect 4062 7964 4068 8016
rect 4120 8004 4126 8016
rect 4120 7976 5672 8004
rect 4120 7964 4126 7976
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 5350 7896 5356 7948
rect 5408 7896 5414 7948
rect 5644 7945 5672 7976
rect 8110 7964 8116 8016
rect 8168 8004 8174 8016
rect 8754 8004 8760 8016
rect 8168 7976 8760 8004
rect 8168 7964 8174 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 10781 8007 10839 8013
rect 10781 7973 10793 8007
rect 10827 7973 10839 8007
rect 10781 7967 10839 7973
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5718 7936 5724 7948
rect 5675 7908 5724 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7561 7939 7619 7945
rect 6972 7908 7144 7936
rect 6972 7896 6978 7908
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 3988 7800 4016 7831
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 5166 7870 5172 7880
rect 5092 7842 5172 7870
rect 4709 7803 4767 7809
rect 3988 7772 4384 7800
rect 3786 7692 3792 7744
rect 3844 7692 3850 7744
rect 4154 7692 4160 7744
rect 4212 7692 4218 7744
rect 4356 7741 4384 7772
rect 4709 7769 4721 7803
rect 4755 7800 4767 7803
rect 5092 7800 5120 7842
rect 5166 7828 5172 7842
rect 5224 7828 5230 7880
rect 7116 7877 7144 7908
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 9214 7936 9220 7948
rect 7607 7908 9220 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7101 7831 7159 7837
rect 7116 7800 7144 7831
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7852 7877 7880 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 10505 7939 10563 7945
rect 9364 7908 9444 7936
rect 9364 7896 9370 7908
rect 9416 7877 9444 7908
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 10551 7908 10640 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7432 7840 7665 7868
rect 7432 7828 7438 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9490 7828 9496 7880
rect 9548 7828 9554 7880
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 10612 7868 10640 7908
rect 10686 7896 10692 7948
rect 10744 7896 10750 7948
rect 10796 7868 10824 7967
rect 10888 7936 10916 8032
rect 18064 7948 18092 8044
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 19705 8075 19763 8081
rect 19705 8041 19717 8075
rect 19751 8072 19763 8075
rect 19886 8072 19892 8084
rect 19751 8044 19892 8072
rect 19751 8041 19763 8044
rect 19705 8035 19763 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 21361 8075 21419 8081
rect 20364 8044 20944 8072
rect 10888 7908 11100 7936
rect 10459 7840 10548 7868
rect 10612 7840 10824 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 4755 7772 7144 7800
rect 4755 7769 4767 7772
rect 4709 7763 4767 7769
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 9122 7800 9128 7812
rect 7248 7772 9128 7800
rect 7248 7760 7254 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9309 7803 9367 7809
rect 9309 7769 9321 7803
rect 9355 7800 9367 7803
rect 9508 7800 9536 7828
rect 9355 7772 9536 7800
rect 10520 7800 10548 7840
rect 10962 7828 10968 7880
rect 11020 7828 11026 7880
rect 11072 7877 11100 7908
rect 12618 7896 12624 7948
rect 12676 7936 12682 7948
rect 13265 7939 13323 7945
rect 13265 7936 13277 7939
rect 12676 7908 13277 7936
rect 12676 7896 12682 7908
rect 13265 7905 13277 7908
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 15381 7939 15439 7945
rect 15381 7905 15393 7939
rect 15427 7936 15439 7939
rect 16022 7936 16028 7948
rect 15427 7908 16028 7936
rect 15427 7905 15439 7908
rect 15381 7899 15439 7905
rect 16022 7896 16028 7908
rect 16080 7936 16086 7948
rect 17218 7936 17224 7948
rect 16080 7908 17224 7936
rect 16080 7896 16086 7908
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7936 17739 7939
rect 18046 7936 18052 7948
rect 17727 7908 18052 7936
rect 17727 7905 17739 7908
rect 17681 7899 17739 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18248 7908 18552 7936
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11256 7800 11284 7831
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 18248 7877 18276 7908
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7837 18475 7871
rect 18417 7831 18475 7837
rect 10520 7772 11284 7800
rect 11609 7803 11667 7809
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 10520 7744 10548 7772
rect 11609 7769 11621 7803
rect 11655 7800 11667 7803
rect 11974 7800 11980 7812
rect 11655 7772 11980 7800
rect 11655 7769 11667 7772
rect 11609 7763 11667 7769
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 15378 7760 15384 7812
rect 15436 7800 15442 7812
rect 15657 7803 15715 7809
rect 15657 7800 15669 7803
rect 15436 7772 15669 7800
rect 15436 7760 15442 7772
rect 15657 7769 15669 7772
rect 15703 7769 15715 7803
rect 15657 7763 15715 7769
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7701 4399 7735
rect 4341 7695 4399 7701
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 6362 7732 6368 7744
rect 4847 7704 6368 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 9398 7692 9404 7744
rect 9456 7692 9462 7744
rect 10042 7692 10048 7744
rect 10100 7692 10106 7744
rect 10502 7692 10508 7744
rect 10560 7692 10566 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 13814 7732 13820 7744
rect 10836 7704 13820 7732
rect 10836 7692 10842 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 18322 7692 18328 7744
rect 18380 7732 18386 7744
rect 18432 7732 18460 7831
rect 18524 7800 18552 7908
rect 18782 7896 18788 7948
rect 18840 7936 18846 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 18840 7908 19257 7936
rect 18840 7896 18846 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 19794 7936 19800 7948
rect 19245 7899 19303 7905
rect 19352 7908 19800 7936
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7858 18751 7871
rect 19352 7868 19380 7908
rect 19794 7896 19800 7908
rect 19852 7936 19858 7948
rect 19852 7908 20116 7936
rect 19852 7896 19858 7908
rect 20088 7880 20116 7908
rect 20254 7896 20260 7948
rect 20312 7936 20318 7948
rect 20364 7945 20392 8044
rect 20916 8004 20944 8044
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 22002 8072 22008 8084
rect 21407 8044 22008 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 25869 8075 25927 8081
rect 25869 8041 25881 8075
rect 25915 8072 25927 8075
rect 25958 8072 25964 8084
rect 25915 8044 25964 8072
rect 25915 8041 25927 8044
rect 25869 8035 25927 8041
rect 25958 8032 25964 8044
rect 26016 8032 26022 8084
rect 22370 8004 22376 8016
rect 20916 7976 22376 8004
rect 22370 7964 22376 7976
rect 22428 7964 22434 8016
rect 22646 8004 22652 8016
rect 22572 7976 22652 8004
rect 22572 7945 22600 7976
rect 22646 7964 22652 7976
rect 22704 7964 22710 8016
rect 25590 7964 25596 8016
rect 25648 8004 25654 8016
rect 25685 8007 25743 8013
rect 25685 8004 25697 8007
rect 25648 7976 25697 8004
rect 25648 7964 25654 7976
rect 25685 7973 25697 7976
rect 25731 7973 25743 8007
rect 25685 7967 25743 7973
rect 20349 7939 20407 7945
rect 20349 7936 20361 7939
rect 20312 7908 20361 7936
rect 20312 7896 20318 7908
rect 20349 7905 20361 7908
rect 20395 7905 20407 7939
rect 20349 7899 20407 7905
rect 22557 7939 22615 7945
rect 22557 7905 22569 7939
rect 22603 7905 22615 7939
rect 22557 7899 22615 7905
rect 18800 7858 19380 7868
rect 18739 7840 19380 7858
rect 18739 7837 18828 7840
rect 18693 7831 18828 7837
rect 18708 7830 18828 7831
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19484 7840 19625 7868
rect 19484 7828 19490 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19978 7868 19984 7880
rect 19613 7831 19671 7837
rect 19720 7840 19984 7868
rect 19444 7800 19472 7828
rect 18524 7772 19472 7800
rect 19720 7744 19748 7840
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20625 7871 20683 7877
rect 20625 7837 20637 7871
rect 20671 7868 20683 7871
rect 20806 7868 20812 7880
rect 20671 7840 20812 7868
rect 20671 7837 20683 7840
rect 20625 7831 20683 7837
rect 20640 7800 20668 7831
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7868 23995 7871
rect 24670 7868 24676 7880
rect 23983 7840 24676 7868
rect 23983 7837 23995 7840
rect 23937 7831 23995 7837
rect 24670 7828 24676 7840
rect 24728 7828 24734 7880
rect 19996 7772 20668 7800
rect 19996 7744 20024 7772
rect 20714 7760 20720 7812
rect 20772 7800 20778 7812
rect 23753 7803 23811 7809
rect 23753 7800 23765 7803
rect 20772 7772 23765 7800
rect 20772 7760 20778 7772
rect 23753 7769 23765 7772
rect 23799 7769 23811 7803
rect 23753 7763 23811 7769
rect 25038 7760 25044 7812
rect 25096 7800 25102 7812
rect 25406 7800 25412 7812
rect 25096 7772 25412 7800
rect 25096 7760 25102 7772
rect 25406 7760 25412 7772
rect 25464 7760 25470 7812
rect 19702 7732 19708 7744
rect 18380 7704 19708 7732
rect 18380 7692 18386 7704
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 19978 7692 19984 7744
rect 20036 7692 20042 7744
rect 1104 7642 30820 7664
rect 1104 7590 5324 7642
rect 5376 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 12752 7642
rect 12804 7590 12816 7642
rect 12868 7590 12880 7642
rect 12932 7590 12944 7642
rect 12996 7590 13008 7642
rect 13060 7590 20180 7642
rect 20232 7590 20244 7642
rect 20296 7590 20308 7642
rect 20360 7590 20372 7642
rect 20424 7590 20436 7642
rect 20488 7590 27608 7642
rect 27660 7590 27672 7642
rect 27724 7590 27736 7642
rect 27788 7590 27800 7642
rect 27852 7590 27864 7642
rect 27916 7590 30820 7642
rect 1104 7568 30820 7590
rect 3786 7488 3792 7540
rect 3844 7488 3850 7540
rect 5166 7488 5172 7540
rect 5224 7488 5230 7540
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 7377 7531 7435 7537
rect 7377 7528 7389 7531
rect 7248 7500 7389 7528
rect 7248 7488 7254 7500
rect 7377 7497 7389 7500
rect 7423 7497 7435 7531
rect 9398 7528 9404 7540
rect 7377 7491 7435 7497
rect 8496 7500 9404 7528
rect 3697 7463 3755 7469
rect 3697 7429 3709 7463
rect 3743 7460 3755 7463
rect 3804 7460 3832 7488
rect 3743 7432 3832 7460
rect 3743 7429 3755 7432
rect 3697 7423 3755 7429
rect 4154 7420 4160 7472
rect 4212 7420 4218 7472
rect 5736 7392 5764 7488
rect 8496 7401 8524 7500
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10042 7488 10048 7540
rect 10100 7488 10106 7540
rect 10888 7500 13308 7528
rect 8662 7420 8668 7472
rect 8720 7420 8726 7472
rect 8803 7463 8861 7469
rect 8803 7429 8815 7463
rect 8849 7460 8861 7463
rect 10060 7460 10088 7488
rect 8849 7432 10088 7460
rect 8849 7429 8861 7432
rect 8803 7423 8861 7429
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 5736 7364 6653 7392
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 8481 7395 8539 7401
rect 8481 7361 8493 7395
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3384 7296 3433 7324
rect 3384 7284 3390 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3436 7188 3464 7287
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 6328 7296 6377 7324
rect 6328 7284 6334 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 4062 7188 4068 7200
rect 3436 7160 4068 7188
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 8294 7148 8300 7200
rect 8352 7148 8358 7200
rect 8588 7188 8616 7355
rect 8680 7324 8708 7420
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9030 7392 9036 7404
rect 8987 7364 9036 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9030 7352 9036 7364
rect 9088 7392 9094 7404
rect 10778 7392 10784 7404
rect 9088 7364 10784 7392
rect 9088 7352 9094 7364
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10888 7324 10916 7500
rect 13280 7469 13308 7500
rect 15930 7488 15936 7540
rect 15988 7488 15994 7540
rect 16574 7488 16580 7540
rect 16632 7488 16638 7540
rect 18046 7528 18052 7540
rect 17512 7500 18052 7528
rect 13265 7463 13323 7469
rect 13265 7429 13277 7463
rect 13311 7460 13323 7463
rect 13311 7432 15516 7460
rect 13311 7429 13323 7432
rect 13265 7423 13323 7429
rect 15488 7404 15516 7432
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11606 7392 11612 7404
rect 11204 7364 11612 7392
rect 11204 7352 11210 7364
rect 11606 7352 11612 7364
rect 11664 7392 11670 7404
rect 11793 7395 11851 7401
rect 11793 7392 11805 7395
rect 11664 7364 11805 7392
rect 11664 7352 11670 7364
rect 11793 7361 11805 7364
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12069 7395 12127 7401
rect 12069 7392 12081 7395
rect 12032 7364 12081 7392
rect 12032 7352 12038 7364
rect 12069 7361 12081 7364
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 13078 7352 13084 7404
rect 13136 7352 13142 7404
rect 13170 7352 13176 7404
rect 13228 7352 13234 7404
rect 13354 7352 13360 7404
rect 13412 7401 13418 7404
rect 13412 7395 13441 7401
rect 13429 7361 13441 7395
rect 13412 7355 13441 7361
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 13906 7392 13912 7404
rect 13863 7364 13912 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 13412 7352 13418 7355
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 14047 7364 14105 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 14093 7355 14151 7361
rect 14200 7364 14381 7392
rect 8680 7296 10916 7324
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7324 13599 7327
rect 13722 7324 13728 7336
rect 13587 7296 13728 7324
rect 13587 7293 13599 7296
rect 13541 7287 13599 7293
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 14016 7324 14044 7355
rect 14200 7324 14228 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 14660 7364 15393 7392
rect 13924 7296 14044 7324
rect 14108 7296 14228 7324
rect 14277 7327 14335 7333
rect 13924 7256 13952 7296
rect 14108 7268 14136 7296
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14568 7324 14596 7352
rect 14323 7296 14596 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 12728 7228 13952 7256
rect 12728 7200 12756 7228
rect 14090 7216 14096 7268
rect 14148 7216 14154 7268
rect 14660 7256 14688 7364
rect 15381 7361 15393 7364
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15286 7324 15292 7336
rect 14292 7228 14688 7256
rect 14752 7296 15292 7324
rect 8938 7188 8944 7200
rect 8588 7160 8944 7188
rect 8938 7148 8944 7160
rect 8996 7188 9002 7200
rect 12710 7188 12716 7200
rect 8996 7160 12716 7188
rect 8996 7148 9002 7160
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 12802 7148 12808 7200
rect 12860 7148 12866 7200
rect 12894 7148 12900 7200
rect 12952 7148 12958 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13228 7160 13645 7188
rect 13228 7148 13234 7160
rect 13633 7157 13645 7160
rect 13679 7188 13691 7191
rect 14292 7188 14320 7228
rect 13679 7160 14320 7188
rect 14369 7191 14427 7197
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 14458 7188 14464 7200
rect 14415 7160 14464 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 14752 7188 14780 7296
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15396 7324 15424 7355
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 15654 7392 15660 7404
rect 15611 7364 15660 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 15764 7364 15853 7392
rect 15396 7296 15608 7324
rect 15580 7268 15608 7296
rect 15562 7216 15568 7268
rect 15620 7216 15626 7268
rect 14599 7160 14780 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15764 7197 15792 7364
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 15841 7355 15899 7361
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16592 7392 16620 7488
rect 16071 7364 16620 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 17512 7333 17540 7500
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 20070 7528 20076 7540
rect 19720 7500 20076 7528
rect 18064 7432 19472 7460
rect 18064 7401 18092 7432
rect 19444 7404 19472 7432
rect 19720 7404 19748 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 20622 7488 20628 7540
rect 20680 7488 20686 7540
rect 20714 7488 20720 7540
rect 20772 7488 20778 7540
rect 23201 7531 23259 7537
rect 23201 7497 23213 7531
rect 23247 7528 23259 7531
rect 24210 7528 24216 7540
rect 23247 7500 24216 7528
rect 23247 7497 23259 7500
rect 23201 7491 23259 7497
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 24670 7488 24676 7540
rect 24728 7488 24734 7540
rect 25038 7488 25044 7540
rect 25096 7488 25102 7540
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 20732 7460 20760 7488
rect 22370 7460 22376 7472
rect 19904 7432 20760 7460
rect 21928 7432 22376 7460
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7361 18107 7395
rect 18049 7355 18107 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18322 7392 18328 7404
rect 18279 7364 18328 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7293 17555 7327
rect 18524 7324 18552 7355
rect 18782 7352 18788 7404
rect 18840 7392 18846 7404
rect 19061 7395 19119 7401
rect 19061 7392 19073 7395
rect 18840 7364 19073 7392
rect 18840 7352 18846 7364
rect 19061 7361 19073 7364
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19702 7352 19708 7404
rect 19760 7352 19766 7404
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 19812 7324 19840 7352
rect 19904 7333 19932 7432
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 21928 7392 21956 7432
rect 22370 7420 22376 7432
rect 22428 7420 22434 7472
rect 23293 7463 23351 7469
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24688 7460 24716 7488
rect 23339 7432 24716 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 21867 7364 21956 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 18524 7296 19840 7324
rect 17497 7287 17555 7293
rect 19812 7256 19840 7296
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 19996 7324 20024 7355
rect 22002 7352 22008 7404
rect 22060 7392 22066 7404
rect 22097 7395 22155 7401
rect 22097 7392 22109 7395
rect 22060 7364 22109 7392
rect 22060 7352 22066 7364
rect 22097 7361 22109 7364
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 25133 7395 25191 7401
rect 25133 7392 25145 7395
rect 24636 7364 25145 7392
rect 24636 7352 24642 7364
rect 25133 7361 25145 7364
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 20162 7324 20168 7336
rect 19996 7296 20168 7324
rect 19996 7256 20024 7296
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 23014 7324 23020 7336
rect 20809 7287 20867 7293
rect 22756 7296 23020 7324
rect 19812 7228 20024 7256
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15344 7160 15761 7188
rect 15344 7148 15350 7160
rect 15749 7157 15761 7160
rect 15795 7157 15807 7191
rect 15749 7151 15807 7157
rect 17954 7148 17960 7200
rect 18012 7148 18018 7200
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19944 7160 20177 7188
rect 19944 7148 19950 7160
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 20165 7151 20223 7157
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 20824 7188 20852 7287
rect 22756 7188 22784 7296
rect 23014 7284 23020 7296
rect 23072 7284 23078 7336
rect 22833 7259 22891 7265
rect 22833 7225 22845 7259
rect 22879 7256 22891 7259
rect 22922 7256 22928 7268
rect 22879 7228 22928 7256
rect 22879 7225 22891 7228
rect 22833 7219 22891 7225
rect 22922 7216 22928 7228
rect 22980 7256 22986 7268
rect 24949 7259 25007 7265
rect 24949 7256 24961 7259
rect 22980 7228 24961 7256
rect 22980 7216 22986 7228
rect 24949 7225 24961 7228
rect 24995 7225 25007 7259
rect 24949 7219 25007 7225
rect 20312 7160 22784 7188
rect 20312 7148 20318 7160
rect 23658 7148 23664 7200
rect 23716 7148 23722 7200
rect 24964 7188 24992 7219
rect 25225 7191 25283 7197
rect 25225 7188 25237 7191
rect 24964 7160 25237 7188
rect 25225 7157 25237 7160
rect 25271 7157 25283 7191
rect 25225 7151 25283 7157
rect 1104 7098 30820 7120
rect 1104 7046 4664 7098
rect 4716 7046 4728 7098
rect 4780 7046 4792 7098
rect 4844 7046 4856 7098
rect 4908 7046 4920 7098
rect 4972 7046 12092 7098
rect 12144 7046 12156 7098
rect 12208 7046 12220 7098
rect 12272 7046 12284 7098
rect 12336 7046 12348 7098
rect 12400 7046 19520 7098
rect 19572 7046 19584 7098
rect 19636 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 26948 7098
rect 27000 7046 27012 7098
rect 27064 7046 27076 7098
rect 27128 7046 27140 7098
rect 27192 7046 27204 7098
rect 27256 7046 30820 7098
rect 1104 7024 30820 7046
rect 4982 6944 4988 6996
rect 5040 6984 5046 6996
rect 5040 6956 6776 6984
rect 5040 6944 5046 6956
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 4028 6888 6684 6916
rect 4028 6876 4034 6888
rect 6656 6789 6684 6888
rect 6748 6848 6776 6956
rect 9122 6944 9128 6996
rect 9180 6944 9186 6996
rect 10502 6944 10508 6996
rect 10560 6944 10566 6996
rect 12710 6944 12716 6996
rect 12768 6944 12774 6996
rect 13078 6944 13084 6996
rect 13136 6944 13142 6996
rect 13262 6944 13268 6996
rect 13320 6944 13326 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14918 6984 14924 6996
rect 13872 6956 14924 6984
rect 13872 6944 13878 6956
rect 14918 6944 14924 6956
rect 14976 6984 14982 6996
rect 16390 6984 16396 6996
rect 14976 6956 16396 6984
rect 14976 6944 14982 6956
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 20254 6984 20260 6996
rect 16776 6956 20260 6984
rect 8220 6888 8432 6916
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 6748 6820 7665 6848
rect 7653 6817 7665 6820
rect 7699 6848 7711 6851
rect 8220 6848 8248 6888
rect 7699 6820 8248 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 8294 6808 8300 6860
rect 8352 6808 8358 6860
rect 8404 6848 8432 6888
rect 9416 6888 10732 6916
rect 9416 6848 9444 6888
rect 8404 6820 9444 6848
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9539 6820 9873 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9861 6817 9873 6820
rect 9907 6848 9919 6851
rect 10704 6848 10732 6888
rect 11698 6848 11704 6860
rect 9907 6820 10640 6848
rect 10704 6820 11704 6848
rect 9907 6817 9919 6820
rect 9861 6811 9919 6817
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 8312 6780 8340 6808
rect 10612 6792 10640 6820
rect 11698 6808 11704 6820
rect 11756 6848 11762 6860
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 11756 6820 12081 6848
rect 11756 6808 11762 6820
rect 12069 6817 12081 6820
rect 12115 6817 12127 6851
rect 12728 6848 12756 6944
rect 13906 6916 13912 6928
rect 13280 6888 13912 6916
rect 12728 6820 13032 6848
rect 12069 6811 12127 6817
rect 7515 6752 8340 6780
rect 9033 6783 9091 6789
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 9033 6749 9045 6783
rect 9079 6780 9091 6783
rect 9306 6780 9312 6792
rect 9079 6752 9312 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 6472 6712 6500 6743
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9508 6752 10333 6780
rect 6472 6684 7052 6712
rect 6086 6604 6092 6656
rect 6144 6644 6150 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 6144 6616 6285 6644
rect 6144 6604 6150 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 6730 6604 6736 6656
rect 6788 6604 6794 6656
rect 7024 6653 7052 6684
rect 9508 6656 9536 6752
rect 10321 6749 10333 6752
rect 10367 6780 10379 6783
rect 10413 6783 10471 6789
rect 10413 6780 10425 6783
rect 10367 6752 10425 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10413 6749 10425 6752
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12894 6780 12900 6792
rect 12023 6752 12900 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13004 6789 13032 6820
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6780 13231 6783
rect 13280 6780 13308 6888
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14461 6851 14519 6857
rect 14461 6848 14473 6851
rect 13648 6820 14473 6848
rect 13219 6752 13308 6780
rect 13219 6749 13231 6752
rect 13173 6743 13231 6749
rect 13280 6724 13308 6752
rect 13444 6783 13502 6789
rect 13444 6749 13456 6783
rect 13490 6780 13502 6783
rect 13648 6780 13676 6820
rect 14461 6817 14473 6820
rect 14507 6848 14519 6851
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14507 6820 14749 6848
rect 14507 6817 14519 6820
rect 14461 6811 14519 6817
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16776 6848 16804 6956
rect 20254 6944 20260 6956
rect 20312 6944 20318 6996
rect 17954 6876 17960 6928
rect 18012 6876 18018 6928
rect 20088 6888 22094 6916
rect 15896 6820 16804 6848
rect 17405 6851 17463 6857
rect 15896 6808 15902 6820
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 17972 6848 18000 6876
rect 17451 6820 18000 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 18782 6808 18788 6860
rect 18840 6848 18846 6860
rect 20088 6857 20116 6888
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18840 6820 19257 6848
rect 18840 6808 18846 6820
rect 19245 6817 19257 6820
rect 19291 6817 19303 6851
rect 19245 6811 19303 6817
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 21358 6808 21364 6860
rect 21416 6848 21422 6860
rect 21910 6848 21916 6860
rect 21416 6820 21916 6848
rect 21416 6808 21422 6820
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22066 6848 22094 6888
rect 22373 6851 22431 6857
rect 22373 6848 22385 6851
rect 22066 6820 22385 6848
rect 22373 6817 22385 6820
rect 22419 6817 22431 6851
rect 22373 6811 22431 6817
rect 22830 6808 22836 6860
rect 22888 6808 22894 6860
rect 23014 6808 23020 6860
rect 23072 6848 23078 6860
rect 23201 6851 23259 6857
rect 23201 6848 23213 6851
rect 23072 6820 23213 6848
rect 23072 6808 23078 6820
rect 23201 6817 23213 6820
rect 23247 6817 23259 6851
rect 23201 6811 23259 6817
rect 13490 6752 13676 6780
rect 13490 6749 13502 6752
rect 13444 6743 13502 6749
rect 13722 6740 13728 6792
rect 13780 6789 13786 6792
rect 13780 6783 13819 6789
rect 13807 6749 13819 6783
rect 13780 6743 13819 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13955 6752 14105 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 13780 6740 13786 6743
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 11238 6712 11244 6724
rect 10152 6684 11244 6712
rect 7009 6647 7067 6653
rect 7009 6613 7021 6647
rect 7055 6613 7067 6647
rect 7009 6607 7067 6613
rect 7377 6647 7435 6653
rect 7377 6613 7389 6647
rect 7423 6644 7435 6647
rect 7466 6644 7472 6656
rect 7423 6616 7472 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 10152 6653 10180 6684
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11900 6684 12434 6712
rect 10137 6647 10195 6653
rect 10137 6613 10149 6647
rect 10183 6613 10195 6647
rect 10137 6607 10195 6613
rect 10229 6647 10287 6653
rect 10229 6613 10241 6647
rect 10275 6644 10287 6647
rect 10686 6644 10692 6656
rect 10275 6616 10692 6644
rect 10275 6613 10287 6616
rect 10229 6607 10287 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11514 6604 11520 6656
rect 11572 6604 11578 6656
rect 11900 6653 11928 6684
rect 11885 6647 11943 6653
rect 11885 6613 11897 6647
rect 11931 6613 11943 6647
rect 12406 6644 12434 6684
rect 12802 6672 12808 6724
rect 12860 6712 12866 6724
rect 13262 6712 13268 6724
rect 12860 6684 13268 6712
rect 12860 6672 12866 6684
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6681 13599 6715
rect 13541 6675 13599 6681
rect 13446 6644 13452 6656
rect 12406 6616 13452 6644
rect 11885 6607 11943 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 13556 6644 13584 6675
rect 13630 6672 13636 6724
rect 13688 6672 13694 6724
rect 14568 6644 14596 6743
rect 14826 6740 14832 6792
rect 14884 6740 14890 6792
rect 14918 6740 14924 6792
rect 14976 6740 14982 6792
rect 15079 6783 15137 6789
rect 15079 6749 15091 6783
rect 15125 6780 15137 6783
rect 15212 6780 15240 6808
rect 15125 6752 15240 6780
rect 15125 6749 15137 6752
rect 15079 6743 15137 6749
rect 15286 6740 15292 6792
rect 15344 6740 15350 6792
rect 15378 6740 15384 6792
rect 15436 6740 15442 6792
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 15611 6752 15945 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 15933 6743 15991 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 15197 6715 15255 6721
rect 15197 6681 15209 6715
rect 15243 6712 15255 6715
rect 15470 6712 15476 6724
rect 15243 6684 15476 6712
rect 15243 6681 15255 6684
rect 15197 6675 15255 6681
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 16025 6715 16083 6721
rect 16025 6712 16037 6715
rect 15580 6684 16037 6712
rect 15580 6644 15608 6684
rect 16025 6681 16037 6684
rect 16071 6712 16083 6715
rect 17236 6712 17264 6743
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19484 6752 19625 6780
rect 19484 6740 19490 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6749 20039 6783
rect 19981 6743 20039 6749
rect 19996 6712 20024 6743
rect 20162 6740 20168 6792
rect 20220 6740 20226 6792
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6749 22615 6783
rect 22848 6780 22876 6808
rect 23109 6783 23167 6789
rect 23109 6780 23121 6783
rect 22848 6752 23121 6780
rect 22557 6743 22615 6749
rect 23109 6749 23121 6752
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6780 23535 6783
rect 23658 6780 23664 6792
rect 23523 6752 23664 6780
rect 23523 6749 23535 6752
rect 23477 6743 23535 6749
rect 20070 6712 20076 6724
rect 16071 6684 17816 6712
rect 19996 6684 20076 6712
rect 16071 6681 16083 6684
rect 16025 6675 16083 6681
rect 17788 6656 17816 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 22572 6712 22600 6743
rect 23658 6740 23664 6752
rect 23716 6740 23722 6792
rect 22572 6684 23060 6712
rect 13556 6616 15608 6644
rect 16390 6604 16396 6656
rect 16448 6604 16454 6656
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 23032 6653 23060 6684
rect 22649 6647 22707 6653
rect 22649 6644 22661 6647
rect 21416 6616 22661 6644
rect 21416 6604 21422 6616
rect 22649 6613 22661 6616
rect 22695 6613 22707 6647
rect 22649 6607 22707 6613
rect 23017 6647 23075 6653
rect 23017 6613 23029 6647
rect 23063 6644 23075 6647
rect 23566 6644 23572 6656
rect 23063 6616 23572 6644
rect 23063 6613 23075 6616
rect 23017 6607 23075 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 23661 6647 23719 6653
rect 23661 6613 23673 6647
rect 23707 6644 23719 6647
rect 23842 6644 23848 6656
rect 23707 6616 23848 6644
rect 23707 6613 23719 6616
rect 23661 6607 23719 6613
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 1104 6554 30820 6576
rect 1104 6502 5324 6554
rect 5376 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 12752 6554
rect 12804 6502 12816 6554
rect 12868 6502 12880 6554
rect 12932 6502 12944 6554
rect 12996 6502 13008 6554
rect 13060 6502 20180 6554
rect 20232 6502 20244 6554
rect 20296 6502 20308 6554
rect 20360 6502 20372 6554
rect 20424 6502 20436 6554
rect 20488 6502 27608 6554
rect 27660 6502 27672 6554
rect 27724 6502 27736 6554
rect 27788 6502 27800 6554
rect 27852 6502 27864 6554
rect 27916 6502 30820 6554
rect 1104 6480 30820 6502
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9364 6412 9413 6440
rect 9364 6400 9370 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 11514 6400 11520 6452
rect 11572 6400 11578 6452
rect 13722 6440 13728 6452
rect 12406 6412 13728 6440
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 9324 6276 10149 6304
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7524 6208 7604 6236
rect 7524 6196 7530 6208
rect 7576 6168 7604 6208
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9324 6236 9352 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 10612 6304 10640 6400
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 10612 6276 10701 6304
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 11146 6304 11152 6316
rect 10689 6267 10747 6273
rect 10796 6276 11152 6304
rect 8444 6208 9352 6236
rect 10413 6239 10471 6245
rect 8444 6196 8450 6208
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10796 6236 10824 6276
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11256 6313 11284 6400
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6273 11299 6307
rect 11532 6304 11560 6400
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11532 6276 11713 6304
rect 11241 6267 11299 6273
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 10459 6208 10824 6236
rect 10873 6239 10931 6245
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10873 6205 10885 6239
rect 10919 6205 10931 6239
rect 11256 6236 11284 6267
rect 12406 6236 12434 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15436 6412 15577 6440
rect 15436 6400 15442 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 16022 6400 16028 6452
rect 16080 6400 16086 6452
rect 19168 6412 23704 6440
rect 16040 6372 16068 6400
rect 19168 6372 19196 6412
rect 16040 6344 19196 6372
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15562 6304 15568 6316
rect 15519 6276 15568 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6304 16083 6307
rect 16390 6304 16396 6316
rect 16071 6276 16396 6304
rect 16071 6273 16083 6276
rect 16025 6267 16083 6273
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 18046 6264 18052 6316
rect 18104 6264 18110 6316
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6304 18383 6307
rect 18414 6304 18420 6316
rect 18371 6276 18420 6304
rect 18371 6273 18383 6276
rect 18325 6267 18383 6273
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 19168 6313 19196 6344
rect 20162 6332 20168 6384
rect 20220 6332 20226 6384
rect 19153 6307 19211 6313
rect 19153 6273 19165 6307
rect 19199 6273 19211 6307
rect 19153 6267 19211 6273
rect 21358 6264 21364 6316
rect 21416 6264 21422 6316
rect 21836 6313 21864 6412
rect 22554 6332 22560 6384
rect 22612 6332 22618 6384
rect 23676 6313 23704 6412
rect 23842 6400 23848 6452
rect 23900 6440 23906 6452
rect 23900 6412 23980 6440
rect 23900 6400 23906 6412
rect 23952 6381 23980 6412
rect 24670 6400 24676 6452
rect 24728 6440 24734 6452
rect 25409 6443 25467 6449
rect 25409 6440 25421 6443
rect 24728 6412 25421 6440
rect 24728 6400 24734 6412
rect 25409 6409 25421 6412
rect 25455 6409 25467 6443
rect 25409 6403 25467 6409
rect 23937 6375 23995 6381
rect 23937 6341 23949 6375
rect 23983 6341 23995 6375
rect 23937 6335 23995 6341
rect 24394 6332 24400 6384
rect 24452 6332 24458 6384
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 11256 6208 12434 6236
rect 10873 6199 10931 6205
rect 9122 6168 9128 6180
rect 7576 6140 9128 6168
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10888 6100 10916 6199
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 15286 6236 15292 6248
rect 14884 6208 15292 6236
rect 14884 6196 14890 6208
rect 15286 6196 15292 6208
rect 15344 6236 15350 6248
rect 15672 6236 15700 6264
rect 15344 6208 17356 6236
rect 15344 6196 15350 6208
rect 11238 6128 11244 6180
rect 11296 6128 11302 6180
rect 17328 6177 17356 6208
rect 19426 6196 19432 6248
rect 19484 6196 19490 6248
rect 22097 6239 22155 6245
rect 22097 6236 22109 6239
rect 21560 6208 22109 6236
rect 17313 6171 17371 6177
rect 17313 6137 17325 6171
rect 17359 6137 17371 6171
rect 17313 6131 17371 6137
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 21560 6177 21588 6208
rect 22097 6205 22109 6208
rect 22143 6205 22155 6239
rect 24578 6236 24584 6248
rect 22097 6199 22155 6205
rect 23768 6208 24584 6236
rect 20901 6171 20959 6177
rect 20901 6168 20913 6171
rect 20588 6140 20913 6168
rect 20588 6128 20594 6140
rect 20901 6137 20913 6140
rect 20947 6137 20959 6171
rect 20901 6131 20959 6137
rect 21545 6171 21603 6177
rect 21545 6137 21557 6171
rect 21591 6137 21603 6171
rect 21545 6131 21603 6137
rect 23566 6128 23572 6180
rect 23624 6168 23630 6180
rect 23768 6168 23796 6208
rect 24578 6196 24584 6208
rect 24636 6196 24642 6248
rect 23624 6140 23796 6168
rect 23624 6128 23630 6140
rect 9548 6072 10916 6100
rect 9548 6060 9554 6072
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16298 6100 16304 6112
rect 16255 6072 16304 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 1104 6010 30820 6032
rect 1104 5958 4664 6010
rect 4716 5958 4728 6010
rect 4780 5958 4792 6010
rect 4844 5958 4856 6010
rect 4908 5958 4920 6010
rect 4972 5958 12092 6010
rect 12144 5958 12156 6010
rect 12208 5958 12220 6010
rect 12272 5958 12284 6010
rect 12336 5958 12348 6010
rect 12400 5958 19520 6010
rect 19572 5958 19584 6010
rect 19636 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 26948 6010
rect 27000 5958 27012 6010
rect 27064 5958 27076 6010
rect 27128 5958 27140 6010
rect 27192 5958 27204 6010
rect 27256 5958 30820 6010
rect 1104 5936 30820 5958
rect 5984 5899 6042 5905
rect 5984 5865 5996 5899
rect 6030 5896 6042 5899
rect 6086 5896 6092 5908
rect 6030 5868 6092 5896
rect 6030 5865 6042 5868
rect 5984 5859 6042 5865
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 9490 5856 9496 5908
rect 9548 5856 9554 5908
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 12805 5899 12863 5905
rect 11296 5868 12434 5896
rect 11296 5856 11302 5868
rect 4062 5720 4068 5772
rect 4120 5760 4126 5772
rect 5721 5763 5779 5769
rect 5721 5760 5733 5763
rect 4120 5732 5733 5760
rect 4120 5720 4126 5732
rect 5721 5729 5733 5732
rect 5767 5760 5779 5763
rect 7006 5760 7012 5772
rect 5767 5732 7012 5760
rect 5767 5729 5779 5732
rect 5721 5723 5779 5729
rect 7006 5720 7012 5732
rect 7064 5760 7070 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 7064 5732 10517 5760
rect 7064 5720 7070 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11514 5760 11520 5772
rect 10827 5732 11520 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12406 5760 12434 5868
rect 12805 5865 12817 5899
rect 12851 5896 12863 5899
rect 13354 5896 13360 5908
rect 12851 5868 13360 5896
rect 12851 5865 12863 5868
rect 12805 5859 12863 5865
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 13817 5899 13875 5905
rect 13817 5865 13829 5899
rect 13863 5896 13875 5899
rect 14274 5896 14280 5908
rect 13863 5868 14280 5896
rect 13863 5865 13875 5868
rect 13817 5859 13875 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 17770 5896 17776 5908
rect 15212 5868 17776 5896
rect 13446 5788 13452 5840
rect 13504 5828 13510 5840
rect 13633 5831 13691 5837
rect 13633 5828 13645 5831
rect 13504 5800 13645 5828
rect 13504 5788 13510 5800
rect 13633 5797 13645 5800
rect 13679 5797 13691 5831
rect 14292 5828 14320 5856
rect 14292 5800 14596 5828
rect 13633 5791 13691 5797
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12406 5732 12633 5760
rect 12621 5729 12633 5732
rect 12667 5760 12679 5763
rect 12667 5732 14320 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5692 9091 5695
rect 9122 5692 9128 5704
rect 9079 5664 9128 5692
rect 9079 5661 9091 5664
rect 9033 5655 9091 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 14090 5652 14096 5704
rect 14148 5652 14154 5704
rect 14292 5701 14320 5732
rect 14568 5701 14596 5800
rect 15212 5701 15240 5868
rect 17770 5856 17776 5868
rect 17828 5856 17834 5908
rect 19426 5856 19432 5908
rect 19484 5856 19490 5908
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 20257 5899 20315 5905
rect 20257 5896 20269 5899
rect 20220 5868 20269 5896
rect 20220 5856 20226 5868
rect 20257 5865 20269 5868
rect 20303 5865 20315 5899
rect 20257 5859 20315 5865
rect 22465 5899 22523 5905
rect 22465 5865 22477 5899
rect 22511 5896 22523 5899
rect 22554 5896 22560 5908
rect 22511 5868 22560 5896
rect 22511 5865 22523 5868
rect 22465 5859 22523 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 23569 5899 23627 5905
rect 23569 5865 23581 5899
rect 23615 5896 23627 5899
rect 24394 5896 24400 5908
rect 23615 5868 24400 5896
rect 23615 5865 23627 5868
rect 23569 5859 23627 5865
rect 24394 5856 24400 5868
rect 24452 5856 24458 5908
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 16022 5720 16028 5772
rect 16080 5720 16086 5772
rect 16298 5720 16304 5772
rect 16356 5720 16362 5772
rect 18248 5732 20208 5760
rect 18248 5704 18276 5732
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 18141 5695 18199 5701
rect 18141 5661 18153 5695
rect 18187 5692 18199 5695
rect 18230 5692 18236 5704
rect 18187 5664 18236 5692
rect 18187 5661 18199 5664
rect 18141 5655 18199 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19886 5692 19892 5704
rect 19659 5664 19892 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 20180 5701 20208 5732
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 22373 5695 22431 5701
rect 22373 5692 22385 5695
rect 20211 5664 22385 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 22373 5661 22385 5664
rect 22419 5692 22431 5695
rect 23477 5695 23535 5701
rect 23477 5692 23489 5695
rect 22419 5664 23489 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 23477 5661 23489 5664
rect 23523 5661 23535 5695
rect 23477 5655 23535 5661
rect 6730 5584 6736 5636
rect 6788 5584 6794 5636
rect 11514 5584 11520 5636
rect 11572 5584 11578 5636
rect 13262 5584 13268 5636
rect 13320 5624 13326 5636
rect 13357 5627 13415 5633
rect 13357 5624 13369 5627
rect 13320 5596 13369 5624
rect 13320 5584 13326 5596
rect 13357 5593 13369 5596
rect 13403 5593 13415 5627
rect 18049 5627 18107 5633
rect 18049 5624 18061 5627
rect 17526 5596 18061 5624
rect 13357 5587 13415 5593
rect 18049 5593 18061 5596
rect 18095 5593 18107 5627
rect 18049 5587 18107 5593
rect 12250 5516 12256 5568
rect 12308 5556 12314 5568
rect 13446 5556 13452 5568
rect 12308 5528 13452 5556
rect 12308 5516 12314 5528
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 14734 5516 14740 5568
rect 14792 5516 14798 5568
rect 14826 5516 14832 5568
rect 14884 5516 14890 5568
rect 1104 5466 30820 5488
rect 1104 5414 5324 5466
rect 5376 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 12752 5466
rect 12804 5414 12816 5466
rect 12868 5414 12880 5466
rect 12932 5414 12944 5466
rect 12996 5414 13008 5466
rect 13060 5414 20180 5466
rect 20232 5414 20244 5466
rect 20296 5414 20308 5466
rect 20360 5414 20372 5466
rect 20424 5414 20436 5466
rect 20488 5414 27608 5466
rect 27660 5414 27672 5466
rect 27724 5414 27736 5466
rect 27788 5414 27800 5466
rect 27852 5414 27864 5466
rect 27916 5414 30820 5466
rect 1104 5392 30820 5414
rect 11514 5312 11520 5364
rect 11572 5352 11578 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11572 5324 11621 5352
rect 11572 5312 11578 5324
rect 11609 5321 11621 5324
rect 11655 5321 11667 5355
rect 11609 5315 11667 5321
rect 12526 5312 12532 5364
rect 12584 5352 12590 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 12584 5324 12633 5352
rect 12584 5312 12590 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 12621 5315 12679 5321
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13630 5352 13636 5364
rect 13035 5324 13636 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11882 5216 11888 5228
rect 11563 5188 11888 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12636 5216 12664 5315
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14148 5324 14289 5352
rect 14148 5312 14154 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 13446 5244 13452 5296
rect 13504 5284 13510 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 13504 5256 13829 5284
rect 13504 5244 13510 5256
rect 13817 5253 13829 5256
rect 13863 5253 13875 5287
rect 13817 5247 13875 5253
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12636 5188 13185 5216
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 14826 5216 14832 5228
rect 13403 5188 14832 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 13262 5148 13268 5160
rect 12391 5120 13268 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 13262 5108 13268 5120
rect 13320 5148 13326 5160
rect 13320 5120 14136 5148
rect 13320 5108 13326 5120
rect 14108 5089 14136 5120
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 14093 5083 14151 5089
rect 14093 5049 14105 5083
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 1104 4922 30820 4944
rect 1104 4870 4664 4922
rect 4716 4870 4728 4922
rect 4780 4870 4792 4922
rect 4844 4870 4856 4922
rect 4908 4870 4920 4922
rect 4972 4870 12092 4922
rect 12144 4870 12156 4922
rect 12208 4870 12220 4922
rect 12272 4870 12284 4922
rect 12336 4870 12348 4922
rect 12400 4870 19520 4922
rect 19572 4870 19584 4922
rect 19636 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 26948 4922
rect 27000 4870 27012 4922
rect 27064 4870 27076 4922
rect 27128 4870 27140 4922
rect 27192 4870 27204 4922
rect 27256 4870 30820 4922
rect 1104 4848 30820 4870
rect 1104 4378 30820 4400
rect 1104 4326 5324 4378
rect 5376 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 12752 4378
rect 12804 4326 12816 4378
rect 12868 4326 12880 4378
rect 12932 4326 12944 4378
rect 12996 4326 13008 4378
rect 13060 4326 20180 4378
rect 20232 4326 20244 4378
rect 20296 4326 20308 4378
rect 20360 4326 20372 4378
rect 20424 4326 20436 4378
rect 20488 4326 27608 4378
rect 27660 4326 27672 4378
rect 27724 4326 27736 4378
rect 27788 4326 27800 4378
rect 27852 4326 27864 4378
rect 27916 4326 30820 4378
rect 1104 4304 30820 4326
rect 14826 4088 14832 4140
rect 14884 4128 14890 4140
rect 16114 4128 16120 4140
rect 14884 4100 16120 4128
rect 14884 4088 14890 4100
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 17402 4088 17408 4140
rect 17460 4128 17466 4140
rect 18138 4128 18144 4140
rect 17460 4100 18144 4128
rect 17460 4088 17466 4100
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 1104 3834 30820 3856
rect 1104 3782 4664 3834
rect 4716 3782 4728 3834
rect 4780 3782 4792 3834
rect 4844 3782 4856 3834
rect 4908 3782 4920 3834
rect 4972 3782 12092 3834
rect 12144 3782 12156 3834
rect 12208 3782 12220 3834
rect 12272 3782 12284 3834
rect 12336 3782 12348 3834
rect 12400 3782 19520 3834
rect 19572 3782 19584 3834
rect 19636 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 26948 3834
rect 27000 3782 27012 3834
rect 27064 3782 27076 3834
rect 27128 3782 27140 3834
rect 27192 3782 27204 3834
rect 27256 3782 30820 3834
rect 1104 3760 30820 3782
rect 1104 3290 30820 3312
rect 1104 3238 5324 3290
rect 5376 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 12752 3290
rect 12804 3238 12816 3290
rect 12868 3238 12880 3290
rect 12932 3238 12944 3290
rect 12996 3238 13008 3290
rect 13060 3238 20180 3290
rect 20232 3238 20244 3290
rect 20296 3238 20308 3290
rect 20360 3238 20372 3290
rect 20424 3238 20436 3290
rect 20488 3238 27608 3290
rect 27660 3238 27672 3290
rect 27724 3238 27736 3290
rect 27788 3238 27800 3290
rect 27852 3238 27864 3290
rect 27916 3238 30820 3290
rect 1104 3216 30820 3238
rect 1104 2746 30820 2768
rect 1104 2694 4664 2746
rect 4716 2694 4728 2746
rect 4780 2694 4792 2746
rect 4844 2694 4856 2746
rect 4908 2694 4920 2746
rect 4972 2694 12092 2746
rect 12144 2694 12156 2746
rect 12208 2694 12220 2746
rect 12272 2694 12284 2746
rect 12336 2694 12348 2746
rect 12400 2694 19520 2746
rect 19572 2694 19584 2746
rect 19636 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 26948 2746
rect 27000 2694 27012 2746
rect 27064 2694 27076 2746
rect 27128 2694 27140 2746
rect 27192 2694 27204 2746
rect 27256 2694 30820 2746
rect 1104 2672 30820 2694
rect 1104 2202 30820 2224
rect 1104 2150 5324 2202
rect 5376 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 12752 2202
rect 12804 2150 12816 2202
rect 12868 2150 12880 2202
rect 12932 2150 12944 2202
rect 12996 2150 13008 2202
rect 13060 2150 20180 2202
rect 20232 2150 20244 2202
rect 20296 2150 20308 2202
rect 20360 2150 20372 2202
rect 20424 2150 20436 2202
rect 20488 2150 27608 2202
rect 27660 2150 27672 2202
rect 27724 2150 27736 2202
rect 27788 2150 27800 2202
rect 27852 2150 27864 2202
rect 27916 2150 30820 2202
rect 1104 2128 30820 2150
<< via1 >>
rect 5324 29350 5376 29402
rect 5388 29350 5440 29402
rect 5452 29350 5504 29402
rect 5516 29350 5568 29402
rect 5580 29350 5632 29402
rect 12752 29350 12804 29402
rect 12816 29350 12868 29402
rect 12880 29350 12932 29402
rect 12944 29350 12996 29402
rect 13008 29350 13060 29402
rect 20180 29350 20232 29402
rect 20244 29350 20296 29402
rect 20308 29350 20360 29402
rect 20372 29350 20424 29402
rect 20436 29350 20488 29402
rect 27608 29350 27660 29402
rect 27672 29350 27724 29402
rect 27736 29350 27788 29402
rect 27800 29350 27852 29402
rect 27864 29350 27916 29402
rect 13084 29248 13136 29300
rect 15476 29248 15528 29300
rect 18144 29248 18196 29300
rect 13360 29112 13412 29164
rect 16396 29112 16448 29164
rect 18052 29112 18104 29164
rect 4664 28806 4716 28858
rect 4728 28806 4780 28858
rect 4792 28806 4844 28858
rect 4856 28806 4908 28858
rect 4920 28806 4972 28858
rect 12092 28806 12144 28858
rect 12156 28806 12208 28858
rect 12220 28806 12272 28858
rect 12284 28806 12336 28858
rect 12348 28806 12400 28858
rect 19520 28806 19572 28858
rect 19584 28806 19636 28858
rect 19648 28806 19700 28858
rect 19712 28806 19764 28858
rect 19776 28806 19828 28858
rect 26948 28806 27000 28858
rect 27012 28806 27064 28858
rect 27076 28806 27128 28858
rect 27140 28806 27192 28858
rect 27204 28806 27256 28858
rect 5324 28262 5376 28314
rect 5388 28262 5440 28314
rect 5452 28262 5504 28314
rect 5516 28262 5568 28314
rect 5580 28262 5632 28314
rect 12752 28262 12804 28314
rect 12816 28262 12868 28314
rect 12880 28262 12932 28314
rect 12944 28262 12996 28314
rect 13008 28262 13060 28314
rect 20180 28262 20232 28314
rect 20244 28262 20296 28314
rect 20308 28262 20360 28314
rect 20372 28262 20424 28314
rect 20436 28262 20488 28314
rect 27608 28262 27660 28314
rect 27672 28262 27724 28314
rect 27736 28262 27788 28314
rect 27800 28262 27852 28314
rect 27864 28262 27916 28314
rect 4664 27718 4716 27770
rect 4728 27718 4780 27770
rect 4792 27718 4844 27770
rect 4856 27718 4908 27770
rect 4920 27718 4972 27770
rect 12092 27718 12144 27770
rect 12156 27718 12208 27770
rect 12220 27718 12272 27770
rect 12284 27718 12336 27770
rect 12348 27718 12400 27770
rect 19520 27718 19572 27770
rect 19584 27718 19636 27770
rect 19648 27718 19700 27770
rect 19712 27718 19764 27770
rect 19776 27718 19828 27770
rect 26948 27718 27000 27770
rect 27012 27718 27064 27770
rect 27076 27718 27128 27770
rect 27140 27718 27192 27770
rect 27204 27718 27256 27770
rect 5324 27174 5376 27226
rect 5388 27174 5440 27226
rect 5452 27174 5504 27226
rect 5516 27174 5568 27226
rect 5580 27174 5632 27226
rect 12752 27174 12804 27226
rect 12816 27174 12868 27226
rect 12880 27174 12932 27226
rect 12944 27174 12996 27226
rect 13008 27174 13060 27226
rect 20180 27174 20232 27226
rect 20244 27174 20296 27226
rect 20308 27174 20360 27226
rect 20372 27174 20424 27226
rect 20436 27174 20488 27226
rect 27608 27174 27660 27226
rect 27672 27174 27724 27226
rect 27736 27174 27788 27226
rect 27800 27174 27852 27226
rect 27864 27174 27916 27226
rect 14556 26979 14608 26988
rect 14556 26945 14565 26979
rect 14565 26945 14599 26979
rect 14599 26945 14608 26979
rect 14556 26936 14608 26945
rect 15200 26936 15252 26988
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 18696 26911 18748 26920
rect 18696 26877 18705 26911
rect 18705 26877 18739 26911
rect 18739 26877 18748 26911
rect 18696 26868 18748 26877
rect 19892 26800 19944 26852
rect 14648 26775 14700 26784
rect 14648 26741 14657 26775
rect 14657 26741 14691 26775
rect 14691 26741 14700 26775
rect 14648 26732 14700 26741
rect 15384 26732 15436 26784
rect 17132 26775 17184 26784
rect 17132 26741 17141 26775
rect 17141 26741 17175 26775
rect 17175 26741 17184 26775
rect 17132 26732 17184 26741
rect 4664 26630 4716 26682
rect 4728 26630 4780 26682
rect 4792 26630 4844 26682
rect 4856 26630 4908 26682
rect 4920 26630 4972 26682
rect 12092 26630 12144 26682
rect 12156 26630 12208 26682
rect 12220 26630 12272 26682
rect 12284 26630 12336 26682
rect 12348 26630 12400 26682
rect 19520 26630 19572 26682
rect 19584 26630 19636 26682
rect 19648 26630 19700 26682
rect 19712 26630 19764 26682
rect 19776 26630 19828 26682
rect 26948 26630 27000 26682
rect 27012 26630 27064 26682
rect 27076 26630 27128 26682
rect 27140 26630 27192 26682
rect 27204 26630 27256 26682
rect 17132 26528 17184 26580
rect 19892 26571 19944 26580
rect 19892 26537 19901 26571
rect 19901 26537 19935 26571
rect 19935 26537 19944 26571
rect 19892 26528 19944 26537
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 14372 26324 14424 26376
rect 14740 26299 14792 26308
rect 14740 26265 14749 26299
rect 14749 26265 14783 26299
rect 14783 26265 14792 26299
rect 14740 26256 14792 26265
rect 16212 26367 16264 26376
rect 16212 26333 16221 26367
rect 16221 26333 16255 26367
rect 16255 26333 16264 26367
rect 16212 26324 16264 26333
rect 16764 26324 16816 26376
rect 15200 26231 15252 26240
rect 15200 26197 15209 26231
rect 15209 26197 15243 26231
rect 15243 26197 15252 26231
rect 15200 26188 15252 26197
rect 15568 26231 15620 26240
rect 15568 26197 15577 26231
rect 15577 26197 15611 26231
rect 15611 26197 15620 26231
rect 15568 26188 15620 26197
rect 16948 26231 17000 26240
rect 16948 26197 16957 26231
rect 16957 26197 16991 26231
rect 16991 26197 17000 26231
rect 16948 26188 17000 26197
rect 5324 26086 5376 26138
rect 5388 26086 5440 26138
rect 5452 26086 5504 26138
rect 5516 26086 5568 26138
rect 5580 26086 5632 26138
rect 12752 26086 12804 26138
rect 12816 26086 12868 26138
rect 12880 26086 12932 26138
rect 12944 26086 12996 26138
rect 13008 26086 13060 26138
rect 20180 26086 20232 26138
rect 20244 26086 20296 26138
rect 20308 26086 20360 26138
rect 20372 26086 20424 26138
rect 20436 26086 20488 26138
rect 27608 26086 27660 26138
rect 27672 26086 27724 26138
rect 27736 26086 27788 26138
rect 27800 26086 27852 26138
rect 27864 26086 27916 26138
rect 14096 25984 14148 26036
rect 14556 26027 14608 26036
rect 14556 25993 14565 26027
rect 14565 25993 14599 26027
rect 14599 25993 14608 26027
rect 14556 25984 14608 25993
rect 14740 25984 14792 26036
rect 16212 26027 16264 26036
rect 16212 25993 16221 26027
rect 16221 25993 16255 26027
rect 16255 25993 16264 26027
rect 16212 25984 16264 25993
rect 18696 25984 18748 26036
rect 14648 25916 14700 25968
rect 12808 25848 12860 25900
rect 14372 25848 14424 25900
rect 16948 25959 17000 25968
rect 10876 25780 10928 25832
rect 15384 25848 15436 25900
rect 16948 25925 16982 25959
rect 16982 25925 17000 25959
rect 16948 25916 17000 25925
rect 16764 25848 16816 25900
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 18512 25687 18564 25696
rect 18512 25653 18521 25687
rect 18521 25653 18555 25687
rect 18555 25653 18564 25687
rect 18512 25644 18564 25653
rect 19892 25644 19944 25696
rect 4664 25542 4716 25594
rect 4728 25542 4780 25594
rect 4792 25542 4844 25594
rect 4856 25542 4908 25594
rect 4920 25542 4972 25594
rect 12092 25542 12144 25594
rect 12156 25542 12208 25594
rect 12220 25542 12272 25594
rect 12284 25542 12336 25594
rect 12348 25542 12400 25594
rect 19520 25542 19572 25594
rect 19584 25542 19636 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 26948 25542 27000 25594
rect 27012 25542 27064 25594
rect 27076 25542 27128 25594
rect 27140 25542 27192 25594
rect 27204 25542 27256 25594
rect 12808 25483 12860 25492
rect 12808 25449 12817 25483
rect 12817 25449 12851 25483
rect 12851 25449 12860 25483
rect 12808 25440 12860 25449
rect 12992 25440 13044 25492
rect 10876 25304 10928 25356
rect 14372 25440 14424 25492
rect 15476 25440 15528 25492
rect 18512 25440 18564 25492
rect 15200 25236 15252 25288
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 10968 25168 11020 25220
rect 11888 25168 11940 25220
rect 8484 25100 8536 25152
rect 9404 25143 9456 25152
rect 9404 25109 9413 25143
rect 9413 25109 9447 25143
rect 9447 25109 9456 25143
rect 9404 25100 9456 25109
rect 12348 25143 12400 25152
rect 12348 25109 12357 25143
rect 12357 25109 12391 25143
rect 12391 25109 12400 25143
rect 12348 25100 12400 25109
rect 20628 25279 20680 25288
rect 20628 25245 20637 25279
rect 20637 25245 20671 25279
rect 20671 25245 20680 25279
rect 20628 25236 20680 25245
rect 17960 25100 18012 25152
rect 18788 25100 18840 25152
rect 5324 24998 5376 25050
rect 5388 24998 5440 25050
rect 5452 24998 5504 25050
rect 5516 24998 5568 25050
rect 5580 24998 5632 25050
rect 12752 24998 12804 25050
rect 12816 24998 12868 25050
rect 12880 24998 12932 25050
rect 12944 24998 12996 25050
rect 13008 24998 13060 25050
rect 20180 24998 20232 25050
rect 20244 24998 20296 25050
rect 20308 24998 20360 25050
rect 20372 24998 20424 25050
rect 20436 24998 20488 25050
rect 27608 24998 27660 25050
rect 27672 24998 27724 25050
rect 27736 24998 27788 25050
rect 27800 24998 27852 25050
rect 27864 24998 27916 25050
rect 9404 24828 9456 24880
rect 8392 24760 8444 24812
rect 10876 24896 10928 24948
rect 10968 24939 11020 24948
rect 10968 24905 10977 24939
rect 10977 24905 11011 24939
rect 11011 24905 11020 24939
rect 10968 24896 11020 24905
rect 11888 24896 11940 24948
rect 6644 24735 6696 24744
rect 6644 24701 6653 24735
rect 6653 24701 6687 24735
rect 6687 24701 6696 24735
rect 6644 24692 6696 24701
rect 9312 24692 9364 24744
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10324 24735 10376 24744
rect 10324 24701 10333 24735
rect 10333 24701 10367 24735
rect 10367 24701 10376 24735
rect 10324 24692 10376 24701
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 17960 24828 18012 24880
rect 10416 24624 10468 24676
rect 6460 24556 6512 24608
rect 7932 24556 7984 24608
rect 9680 24556 9732 24608
rect 11060 24760 11112 24812
rect 12348 24760 12400 24812
rect 15476 24760 15528 24812
rect 16764 24760 16816 24812
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 12440 24556 12492 24608
rect 13084 24735 13136 24744
rect 13084 24701 13093 24735
rect 13093 24701 13127 24735
rect 13127 24701 13136 24735
rect 13084 24692 13136 24701
rect 14188 24624 14240 24676
rect 18512 24624 18564 24676
rect 14372 24556 14424 24608
rect 18144 24599 18196 24608
rect 18144 24565 18153 24599
rect 18153 24565 18187 24599
rect 18187 24565 18196 24599
rect 18144 24556 18196 24565
rect 18880 24599 18932 24608
rect 18880 24565 18889 24599
rect 18889 24565 18923 24599
rect 18923 24565 18932 24599
rect 18880 24556 18932 24565
rect 4664 24454 4716 24506
rect 4728 24454 4780 24506
rect 4792 24454 4844 24506
rect 4856 24454 4908 24506
rect 4920 24454 4972 24506
rect 12092 24454 12144 24506
rect 12156 24454 12208 24506
rect 12220 24454 12272 24506
rect 12284 24454 12336 24506
rect 12348 24454 12400 24506
rect 19520 24454 19572 24506
rect 19584 24454 19636 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 26948 24454 27000 24506
rect 27012 24454 27064 24506
rect 27076 24454 27128 24506
rect 27140 24454 27192 24506
rect 27204 24454 27256 24506
rect 6644 24352 6696 24404
rect 8392 24395 8444 24404
rect 8392 24361 8401 24395
rect 8401 24361 8435 24395
rect 8435 24361 8444 24395
rect 8392 24352 8444 24361
rect 10048 24352 10100 24404
rect 8484 24284 8536 24336
rect 6460 24259 6512 24268
rect 6460 24225 6469 24259
rect 6469 24225 6503 24259
rect 6503 24225 6512 24259
rect 6460 24216 6512 24225
rect 8300 24216 8352 24268
rect 10324 24216 10376 24268
rect 12440 24284 12492 24336
rect 4436 24123 4488 24132
rect 4436 24089 4445 24123
rect 4445 24089 4479 24123
rect 4479 24089 4488 24123
rect 4436 24080 4488 24089
rect 5724 24080 5776 24132
rect 6184 24123 6236 24132
rect 6184 24089 6193 24123
rect 6193 24089 6227 24123
rect 6227 24089 6236 24123
rect 6184 24080 6236 24089
rect 6920 24123 6972 24132
rect 6920 24089 6929 24123
rect 6929 24089 6963 24123
rect 6963 24089 6972 24123
rect 6920 24080 6972 24089
rect 7104 24191 7156 24200
rect 7104 24157 7113 24191
rect 7113 24157 7147 24191
rect 7147 24157 7156 24191
rect 7104 24148 7156 24157
rect 7196 24148 7248 24200
rect 7932 24148 7984 24200
rect 9220 24191 9272 24200
rect 9220 24157 9229 24191
rect 9229 24157 9263 24191
rect 9263 24157 9272 24191
rect 9220 24148 9272 24157
rect 14372 24216 14424 24268
rect 18052 24352 18104 24404
rect 18512 24352 18564 24404
rect 19064 24352 19116 24404
rect 15476 24216 15528 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 18788 24327 18840 24336
rect 18788 24293 18797 24327
rect 18797 24293 18831 24327
rect 18831 24293 18840 24327
rect 18788 24284 18840 24293
rect 8392 24080 8444 24132
rect 9036 24080 9088 24132
rect 9128 24123 9180 24132
rect 9128 24089 9137 24123
rect 9137 24089 9171 24123
rect 9171 24089 9180 24123
rect 9128 24080 9180 24089
rect 8116 24012 8168 24064
rect 14188 24148 14240 24200
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 16764 24148 16816 24200
rect 19248 24148 19300 24200
rect 10692 24123 10744 24132
rect 10692 24089 10701 24123
rect 10701 24089 10735 24123
rect 10735 24089 10744 24123
rect 10692 24080 10744 24089
rect 11060 24012 11112 24064
rect 11980 24012 12032 24064
rect 13084 24012 13136 24064
rect 15568 24080 15620 24132
rect 18144 24123 18196 24132
rect 18144 24089 18162 24123
rect 18162 24089 18196 24123
rect 18144 24080 18196 24089
rect 16304 24055 16356 24064
rect 16304 24021 16313 24055
rect 16313 24021 16347 24055
rect 16347 24021 16356 24055
rect 16304 24012 16356 24021
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 5324 23910 5376 23962
rect 5388 23910 5440 23962
rect 5452 23910 5504 23962
rect 5516 23910 5568 23962
rect 5580 23910 5632 23962
rect 12752 23910 12804 23962
rect 12816 23910 12868 23962
rect 12880 23910 12932 23962
rect 12944 23910 12996 23962
rect 13008 23910 13060 23962
rect 20180 23910 20232 23962
rect 20244 23910 20296 23962
rect 20308 23910 20360 23962
rect 20372 23910 20424 23962
rect 20436 23910 20488 23962
rect 27608 23910 27660 23962
rect 27672 23910 27724 23962
rect 27736 23910 27788 23962
rect 27800 23910 27852 23962
rect 27864 23910 27916 23962
rect 5724 23808 5776 23860
rect 6184 23808 6236 23860
rect 6552 23715 6604 23724
rect 6552 23681 6561 23715
rect 6561 23681 6595 23715
rect 6595 23681 6604 23715
rect 6552 23672 6604 23681
rect 7104 23740 7156 23792
rect 7012 23672 7064 23724
rect 8392 23740 8444 23792
rect 10692 23808 10744 23860
rect 10784 23740 10836 23792
rect 14188 23808 14240 23860
rect 14280 23808 14332 23860
rect 15568 23851 15620 23860
rect 15568 23817 15577 23851
rect 15577 23817 15611 23851
rect 15611 23817 15620 23851
rect 15568 23808 15620 23817
rect 16856 23808 16908 23860
rect 18880 23808 18932 23860
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 9036 23672 9088 23724
rect 11060 23672 11112 23724
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 13636 23672 13688 23724
rect 14556 23672 14608 23724
rect 14740 23672 14792 23724
rect 16304 23740 16356 23792
rect 15476 23715 15528 23724
rect 15476 23681 15485 23715
rect 15485 23681 15519 23715
rect 15519 23681 15528 23715
rect 15476 23672 15528 23681
rect 10508 23604 10560 23656
rect 10416 23536 10468 23588
rect 11152 23536 11204 23588
rect 14372 23604 14424 23656
rect 25412 23740 25464 23792
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 16028 23604 16080 23656
rect 7840 23468 7892 23520
rect 8208 23511 8260 23520
rect 8208 23477 8217 23511
rect 8217 23477 8251 23511
rect 8251 23477 8260 23511
rect 8208 23468 8260 23477
rect 13728 23468 13780 23520
rect 14832 23468 14884 23520
rect 24492 23647 24544 23656
rect 24492 23613 24501 23647
rect 24501 23613 24535 23647
rect 24535 23613 24544 23647
rect 24492 23604 24544 23613
rect 24860 23604 24912 23656
rect 24400 23536 24452 23588
rect 19248 23468 19300 23520
rect 19432 23468 19484 23520
rect 20536 23468 20588 23520
rect 23480 23468 23532 23520
rect 27436 23468 27488 23520
rect 4664 23366 4716 23418
rect 4728 23366 4780 23418
rect 4792 23366 4844 23418
rect 4856 23366 4908 23418
rect 4920 23366 4972 23418
rect 12092 23366 12144 23418
rect 12156 23366 12208 23418
rect 12220 23366 12272 23418
rect 12284 23366 12336 23418
rect 12348 23366 12400 23418
rect 19520 23366 19572 23418
rect 19584 23366 19636 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 26948 23366 27000 23418
rect 27012 23366 27064 23418
rect 27076 23366 27128 23418
rect 27140 23366 27192 23418
rect 27204 23366 27256 23418
rect 6552 23264 6604 23316
rect 6644 23171 6696 23180
rect 6644 23137 6653 23171
rect 6653 23137 6687 23171
rect 6687 23137 6696 23171
rect 6644 23128 6696 23137
rect 7104 23128 7156 23180
rect 7840 23239 7892 23248
rect 7840 23205 7849 23239
rect 7849 23205 7883 23239
rect 7883 23205 7892 23239
rect 7840 23196 7892 23205
rect 8024 23196 8076 23248
rect 9588 23264 9640 23316
rect 11060 23264 11112 23316
rect 12256 23264 12308 23316
rect 13544 23264 13596 23316
rect 24860 23264 24912 23316
rect 25412 23307 25464 23316
rect 25412 23273 25421 23307
rect 25421 23273 25455 23307
rect 25455 23273 25464 23307
rect 25412 23264 25464 23273
rect 27436 23264 27488 23316
rect 11152 23196 11204 23248
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 12440 23128 12492 23180
rect 13268 23196 13320 23248
rect 13636 23196 13688 23248
rect 19340 23128 19392 23180
rect 19984 23128 20036 23180
rect 20628 23128 20680 23180
rect 23940 23128 23992 23180
rect 24492 23128 24544 23180
rect 7932 23103 7984 23112
rect 7932 23069 7953 23103
rect 7953 23069 7984 23103
rect 7932 23060 7984 23069
rect 8208 23060 8260 23112
rect 9220 23060 9272 23112
rect 11980 23103 12032 23112
rect 11980 23069 11989 23103
rect 11989 23069 12023 23103
rect 12023 23069 12032 23103
rect 11980 23060 12032 23069
rect 6552 22924 6604 22976
rect 7012 22924 7064 22976
rect 7472 22967 7524 22976
rect 7472 22933 7481 22967
rect 7481 22933 7515 22967
rect 7515 22933 7524 22967
rect 7472 22924 7524 22933
rect 7748 22924 7800 22976
rect 7840 22924 7892 22976
rect 8484 22924 8536 22976
rect 11888 22992 11940 23044
rect 15660 23060 15712 23112
rect 16028 22992 16080 23044
rect 20536 22992 20588 23044
rect 9312 22967 9364 22976
rect 9312 22933 9339 22967
rect 9339 22933 9364 22967
rect 9312 22924 9364 22933
rect 10508 22924 10560 22976
rect 11612 22924 11664 22976
rect 12256 22924 12308 22976
rect 13176 22967 13228 22976
rect 13176 22933 13185 22967
rect 13185 22933 13219 22967
rect 13219 22933 13228 22967
rect 13176 22924 13228 22933
rect 14924 22967 14976 22976
rect 14924 22933 14933 22967
rect 14933 22933 14967 22967
rect 14967 22933 14976 22967
rect 14924 22924 14976 22933
rect 15752 22924 15804 22976
rect 21916 22924 21968 22976
rect 25136 23103 25188 23112
rect 25136 23069 25145 23103
rect 25145 23069 25179 23103
rect 25179 23069 25188 23103
rect 25136 23060 25188 23069
rect 27988 23060 28040 23112
rect 22744 23035 22796 23044
rect 22744 23001 22753 23035
rect 22753 23001 22787 23035
rect 22787 23001 22796 23035
rect 22744 22992 22796 23001
rect 23480 22992 23532 23044
rect 24400 22992 24452 23044
rect 25228 22992 25280 23044
rect 24216 22967 24268 22976
rect 24216 22933 24225 22967
rect 24225 22933 24259 22967
rect 24259 22933 24268 22967
rect 24216 22924 24268 22933
rect 28908 22924 28960 22976
rect 5324 22822 5376 22874
rect 5388 22822 5440 22874
rect 5452 22822 5504 22874
rect 5516 22822 5568 22874
rect 5580 22822 5632 22874
rect 12752 22822 12804 22874
rect 12816 22822 12868 22874
rect 12880 22822 12932 22874
rect 12944 22822 12996 22874
rect 13008 22822 13060 22874
rect 20180 22822 20232 22874
rect 20244 22822 20296 22874
rect 20308 22822 20360 22874
rect 20372 22822 20424 22874
rect 20436 22822 20488 22874
rect 27608 22822 27660 22874
rect 27672 22822 27724 22874
rect 27736 22822 27788 22874
rect 27800 22822 27852 22874
rect 27864 22822 27916 22874
rect 4436 22763 4488 22772
rect 4436 22729 4445 22763
rect 4445 22729 4479 22763
rect 4479 22729 4488 22763
rect 4436 22720 4488 22729
rect 5172 22652 5224 22704
rect 4160 22559 4212 22568
rect 4160 22525 4169 22559
rect 4169 22525 4203 22559
rect 4203 22525 4212 22559
rect 4160 22516 4212 22525
rect 6092 22652 6144 22704
rect 6644 22763 6696 22772
rect 6644 22729 6653 22763
rect 6653 22729 6687 22763
rect 6687 22729 6696 22763
rect 6644 22720 6696 22729
rect 6920 22720 6972 22772
rect 7656 22720 7708 22772
rect 9128 22720 9180 22772
rect 10508 22763 10560 22772
rect 10508 22729 10517 22763
rect 10517 22729 10551 22763
rect 10551 22729 10560 22763
rect 10508 22720 10560 22729
rect 5908 22627 5960 22636
rect 5908 22593 5917 22627
rect 5917 22593 5951 22627
rect 5951 22593 5960 22627
rect 5908 22584 5960 22593
rect 4988 22380 5040 22432
rect 5080 22380 5132 22432
rect 6920 22584 6972 22636
rect 7196 22584 7248 22636
rect 6552 22559 6604 22568
rect 6552 22525 6570 22559
rect 6570 22525 6604 22559
rect 6552 22516 6604 22525
rect 7748 22584 7800 22636
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 8484 22627 8536 22636
rect 8484 22593 8494 22627
rect 8494 22593 8528 22627
rect 8528 22593 8536 22627
rect 8484 22584 8536 22593
rect 8576 22584 8628 22636
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 8760 22627 8812 22636
rect 8760 22593 8769 22627
rect 8769 22593 8803 22627
rect 8803 22593 8812 22627
rect 8760 22584 8812 22593
rect 10784 22763 10836 22772
rect 10784 22729 10793 22763
rect 10793 22729 10827 22763
rect 10827 22729 10836 22763
rect 10784 22720 10836 22729
rect 11980 22720 12032 22772
rect 12256 22720 12308 22772
rect 9680 22584 9732 22636
rect 8024 22516 8076 22568
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 11060 22627 11112 22636
rect 11060 22593 11069 22627
rect 11069 22593 11103 22627
rect 11103 22593 11112 22627
rect 11060 22584 11112 22593
rect 11428 22652 11480 22704
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 11796 22627 11848 22636
rect 11796 22593 11805 22627
rect 11805 22593 11839 22627
rect 11839 22593 11848 22627
rect 11796 22584 11848 22593
rect 11980 22627 12032 22636
rect 12348 22695 12400 22704
rect 12348 22661 12357 22695
rect 12357 22661 12391 22695
rect 12391 22661 12400 22695
rect 12348 22652 12400 22661
rect 14924 22720 14976 22772
rect 17868 22720 17920 22772
rect 11980 22593 12015 22627
rect 12015 22593 12032 22627
rect 11980 22584 12032 22593
rect 7472 22423 7524 22432
rect 7472 22389 7481 22423
rect 7481 22389 7515 22423
rect 7515 22389 7524 22423
rect 7472 22380 7524 22389
rect 9864 22448 9916 22500
rect 15752 22652 15804 22704
rect 20812 22720 20864 22772
rect 21916 22720 21968 22772
rect 22744 22720 22796 22772
rect 11796 22448 11848 22500
rect 12256 22448 12308 22500
rect 13268 22584 13320 22636
rect 13544 22584 13596 22636
rect 14372 22584 14424 22636
rect 18052 22584 18104 22636
rect 15200 22516 15252 22568
rect 12532 22448 12584 22500
rect 16948 22559 17000 22568
rect 16948 22525 16957 22559
rect 16957 22525 16991 22559
rect 16991 22525 17000 22559
rect 16948 22516 17000 22525
rect 10692 22380 10744 22432
rect 10968 22380 11020 22432
rect 13268 22380 13320 22432
rect 16764 22380 16816 22432
rect 17960 22380 18012 22432
rect 18972 22423 19024 22432
rect 18972 22389 18981 22423
rect 18981 22389 19015 22423
rect 19015 22389 19024 22423
rect 18972 22380 19024 22389
rect 21180 22559 21232 22568
rect 21180 22525 21189 22559
rect 21189 22525 21223 22559
rect 21223 22525 21232 22559
rect 21180 22516 21232 22525
rect 25136 22763 25188 22772
rect 25136 22729 25145 22763
rect 25145 22729 25179 22763
rect 25179 22729 25188 22763
rect 25136 22720 25188 22729
rect 27528 22720 27580 22772
rect 28908 22720 28960 22772
rect 24216 22652 24268 22704
rect 24768 22652 24820 22704
rect 25044 22584 25096 22636
rect 25504 22627 25556 22636
rect 25504 22593 25513 22627
rect 25513 22593 25547 22627
rect 25547 22593 25556 22627
rect 25504 22584 25556 22593
rect 25412 22516 25464 22568
rect 28172 22627 28224 22636
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 28172 22584 28224 22593
rect 20168 22448 20220 22500
rect 24768 22448 24820 22500
rect 19432 22380 19484 22432
rect 19892 22380 19944 22432
rect 22100 22380 22152 22432
rect 26056 22380 26108 22432
rect 27344 22380 27396 22432
rect 28816 22448 28868 22500
rect 28632 22423 28684 22432
rect 28632 22389 28641 22423
rect 28641 22389 28675 22423
rect 28675 22389 28684 22423
rect 28632 22380 28684 22389
rect 29092 22423 29144 22432
rect 29092 22389 29101 22423
rect 29101 22389 29135 22423
rect 29135 22389 29144 22423
rect 29092 22380 29144 22389
rect 29276 22423 29328 22432
rect 29276 22389 29285 22423
rect 29285 22389 29319 22423
rect 29319 22389 29328 22423
rect 29276 22380 29328 22389
rect 4664 22278 4716 22330
rect 4728 22278 4780 22330
rect 4792 22278 4844 22330
rect 4856 22278 4908 22330
rect 4920 22278 4972 22330
rect 12092 22278 12144 22330
rect 12156 22278 12208 22330
rect 12220 22278 12272 22330
rect 12284 22278 12336 22330
rect 12348 22278 12400 22330
rect 19520 22278 19572 22330
rect 19584 22278 19636 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 26948 22278 27000 22330
rect 27012 22278 27064 22330
rect 27076 22278 27128 22330
rect 27140 22278 27192 22330
rect 27204 22278 27256 22330
rect 4160 22219 4212 22228
rect 4160 22185 4169 22219
rect 4169 22185 4203 22219
rect 4203 22185 4212 22219
rect 4160 22176 4212 22185
rect 4988 22176 5040 22228
rect 5908 22176 5960 22228
rect 6736 22176 6788 22228
rect 8576 22176 8628 22228
rect 8668 22176 8720 22228
rect 11704 22176 11756 22228
rect 4436 22040 4488 22092
rect 4344 22015 4396 22024
rect 4344 21981 4353 22015
rect 4353 21981 4387 22015
rect 4387 21981 4396 22015
rect 4344 21972 4396 21981
rect 5172 22040 5224 22092
rect 7196 22040 7248 22092
rect 9312 22040 9364 22092
rect 4988 21972 5040 22024
rect 9220 21972 9272 22024
rect 9864 22108 9916 22160
rect 10968 22108 11020 22160
rect 11060 22040 11112 22092
rect 13636 22176 13688 22228
rect 15660 22219 15712 22228
rect 15660 22185 15669 22219
rect 15669 22185 15703 22219
rect 15703 22185 15712 22219
rect 15660 22176 15712 22185
rect 16948 22219 17000 22228
rect 16948 22185 16957 22219
rect 16957 22185 16991 22219
rect 16991 22185 17000 22219
rect 16948 22176 17000 22185
rect 18052 22176 18104 22228
rect 4436 21836 4488 21888
rect 4528 21879 4580 21888
rect 4528 21845 4537 21879
rect 4537 21845 4571 21879
rect 4571 21845 4580 21879
rect 4528 21836 4580 21845
rect 4620 21836 4672 21888
rect 10048 21972 10100 22024
rect 12532 21972 12584 22024
rect 11428 21904 11480 21956
rect 11704 21904 11756 21956
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9496 21879 9548 21888
rect 9496 21845 9505 21879
rect 9505 21845 9539 21879
rect 9539 21845 9548 21879
rect 9496 21836 9548 21845
rect 9864 21836 9916 21888
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 13084 21904 13136 21956
rect 14004 21972 14056 22024
rect 14832 21972 14884 22024
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 17868 22108 17920 22160
rect 17776 22083 17828 22092
rect 17776 22049 17785 22083
rect 17785 22049 17819 22083
rect 17819 22049 17828 22083
rect 17776 22040 17828 22049
rect 18696 22040 18748 22092
rect 21180 22176 21232 22228
rect 25044 22176 25096 22228
rect 20536 22108 20588 22160
rect 21916 22108 21968 22160
rect 17960 21972 18012 22024
rect 13176 21836 13228 21888
rect 13544 21879 13596 21888
rect 13544 21845 13553 21879
rect 13553 21845 13587 21879
rect 13587 21845 13596 21879
rect 15292 21947 15344 21956
rect 15292 21913 15301 21947
rect 15301 21913 15335 21947
rect 15335 21913 15344 21947
rect 15292 21904 15344 21913
rect 16764 21904 16816 21956
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 19248 21972 19300 22024
rect 19616 21972 19668 22024
rect 19800 22015 19852 22024
rect 19800 21981 19809 22015
rect 19809 21981 19843 22015
rect 19843 21981 19852 22015
rect 19800 21972 19852 21981
rect 20168 21972 20220 22024
rect 25504 22108 25556 22160
rect 27436 22176 27488 22228
rect 27896 22219 27948 22228
rect 27896 22185 27905 22219
rect 27905 22185 27939 22219
rect 27939 22185 27948 22219
rect 27896 22176 27948 22185
rect 26240 22040 26292 22092
rect 18512 21904 18564 21956
rect 13544 21836 13596 21845
rect 13820 21879 13872 21888
rect 13820 21845 13829 21879
rect 13829 21845 13863 21879
rect 13863 21845 13872 21879
rect 13820 21836 13872 21845
rect 14556 21836 14608 21888
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 19800 21836 19852 21888
rect 20812 21836 20864 21888
rect 22100 22015 22152 22024
rect 22100 21981 22109 22015
rect 22109 21981 22143 22015
rect 22143 21981 22152 22015
rect 22100 21972 22152 21981
rect 21180 21947 21232 21956
rect 21180 21913 21189 21947
rect 21189 21913 21223 21947
rect 21223 21913 21232 21947
rect 21180 21904 21232 21913
rect 21548 21904 21600 21956
rect 21824 21947 21876 21956
rect 21824 21913 21833 21947
rect 21833 21913 21867 21947
rect 21867 21913 21876 21947
rect 21824 21904 21876 21913
rect 22560 21904 22612 21956
rect 22192 21879 22244 21888
rect 22192 21845 22201 21879
rect 22201 21845 22235 21879
rect 22235 21845 22244 21879
rect 22192 21836 22244 21845
rect 22284 21836 22336 21888
rect 22836 21904 22888 21956
rect 24032 21972 24084 22024
rect 25320 21904 25372 21956
rect 24400 21836 24452 21888
rect 26332 22015 26384 22024
rect 26332 21981 26354 22015
rect 26354 21981 26384 22015
rect 26332 21972 26384 21981
rect 26884 22015 26936 22024
rect 26884 21981 26893 22015
rect 26893 21981 26927 22015
rect 26927 21981 26936 22015
rect 26884 21972 26936 21981
rect 27252 21972 27304 22024
rect 26240 21947 26292 21956
rect 26240 21913 26249 21947
rect 26249 21913 26283 21947
rect 26283 21913 26292 21947
rect 26240 21904 26292 21913
rect 28172 22108 28224 22160
rect 28816 22108 28868 22160
rect 28632 22015 28684 22024
rect 28632 21981 28641 22015
rect 28641 21981 28675 22015
rect 28675 21981 28684 22015
rect 28632 21972 28684 21981
rect 28816 22015 28868 22024
rect 28816 21981 28825 22015
rect 28825 21981 28859 22015
rect 28859 21981 28868 22015
rect 28816 21972 28868 21981
rect 29092 22015 29144 22024
rect 29092 21981 29101 22015
rect 29101 21981 29135 22015
rect 29135 21981 29144 22015
rect 29092 21972 29144 21981
rect 29276 21947 29328 21956
rect 29276 21913 29285 21947
rect 29285 21913 29319 21947
rect 29319 21913 29328 21947
rect 29276 21904 29328 21913
rect 26884 21836 26936 21888
rect 28080 21836 28132 21888
rect 29368 21836 29420 21888
rect 5324 21734 5376 21786
rect 5388 21734 5440 21786
rect 5452 21734 5504 21786
rect 5516 21734 5568 21786
rect 5580 21734 5632 21786
rect 12752 21734 12804 21786
rect 12816 21734 12868 21786
rect 12880 21734 12932 21786
rect 12944 21734 12996 21786
rect 13008 21734 13060 21786
rect 20180 21734 20232 21786
rect 20244 21734 20296 21786
rect 20308 21734 20360 21786
rect 20372 21734 20424 21786
rect 20436 21734 20488 21786
rect 27608 21734 27660 21786
rect 27672 21734 27724 21786
rect 27736 21734 27788 21786
rect 27800 21734 27852 21786
rect 27864 21734 27916 21786
rect 4344 21632 4396 21684
rect 6828 21632 6880 21684
rect 7104 21632 7156 21684
rect 7656 21632 7708 21684
rect 9220 21632 9272 21684
rect 4528 21564 4580 21616
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 4988 21564 5040 21616
rect 5540 21496 5592 21548
rect 8208 21564 8260 21616
rect 9772 21632 9824 21684
rect 10600 21632 10652 21684
rect 13268 21632 13320 21684
rect 15292 21632 15344 21684
rect 17684 21632 17736 21684
rect 6092 21496 6144 21548
rect 6552 21539 6604 21548
rect 6552 21505 6561 21539
rect 6561 21505 6595 21539
rect 6595 21505 6604 21539
rect 6552 21496 6604 21505
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 11980 21564 12032 21616
rect 16764 21564 16816 21616
rect 18512 21632 18564 21684
rect 18604 21632 18656 21684
rect 19064 21632 19116 21684
rect 19984 21632 20036 21684
rect 10416 21539 10468 21548
rect 10416 21505 10425 21539
rect 10425 21505 10459 21539
rect 10459 21505 10468 21539
rect 10416 21496 10468 21505
rect 10508 21539 10560 21548
rect 10508 21505 10517 21539
rect 10517 21505 10551 21539
rect 10551 21505 10560 21539
rect 10508 21496 10560 21505
rect 10692 21539 10744 21548
rect 10692 21505 10700 21539
rect 10700 21505 10734 21539
rect 10734 21505 10744 21539
rect 10692 21496 10744 21505
rect 10784 21539 10836 21548
rect 10784 21505 10793 21539
rect 10793 21505 10827 21539
rect 10827 21505 10836 21539
rect 10784 21496 10836 21505
rect 12624 21496 12676 21548
rect 9864 21428 9916 21480
rect 11060 21360 11112 21412
rect 13728 21496 13780 21548
rect 14832 21496 14884 21548
rect 17868 21607 17920 21616
rect 17868 21573 17877 21607
rect 17877 21573 17911 21607
rect 17911 21573 17920 21607
rect 17868 21564 17920 21573
rect 21180 21632 21232 21684
rect 22560 21632 22612 21684
rect 24400 21632 24452 21684
rect 26148 21632 26200 21684
rect 20168 21564 20220 21616
rect 940 21292 992 21344
rect 4436 21292 4488 21344
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 6828 21292 6880 21344
rect 8484 21292 8536 21344
rect 9680 21292 9732 21344
rect 10048 21292 10100 21344
rect 13176 21292 13228 21344
rect 15016 21471 15068 21480
rect 15016 21437 15025 21471
rect 15025 21437 15059 21471
rect 15059 21437 15068 21471
rect 15016 21428 15068 21437
rect 15200 21428 15252 21480
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 18788 21496 18840 21548
rect 19892 21496 19944 21548
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 14280 21292 14332 21344
rect 14464 21335 14516 21344
rect 14464 21301 14473 21335
rect 14473 21301 14507 21335
rect 14507 21301 14516 21335
rect 14464 21292 14516 21301
rect 16580 21292 16632 21344
rect 18052 21428 18104 21480
rect 18328 21360 18380 21412
rect 19340 21360 19392 21412
rect 18604 21292 18656 21344
rect 20444 21292 20496 21344
rect 20812 21428 20864 21480
rect 21548 21539 21600 21548
rect 21548 21505 21557 21539
rect 21557 21505 21591 21539
rect 21591 21505 21600 21539
rect 21548 21496 21600 21505
rect 22836 21496 22888 21548
rect 23020 21496 23072 21548
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 24216 21564 24268 21616
rect 26792 21564 26844 21616
rect 27988 21564 28040 21616
rect 22284 21428 22336 21480
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 24032 21428 24084 21480
rect 25320 21428 25372 21480
rect 25872 21539 25924 21548
rect 25872 21505 25881 21539
rect 25881 21505 25915 21539
rect 25915 21505 25924 21539
rect 25872 21496 25924 21505
rect 26424 21496 26476 21548
rect 26976 21496 27028 21548
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 20628 21292 20680 21344
rect 26884 21428 26936 21480
rect 26608 21403 26660 21412
rect 26608 21369 26617 21403
rect 26617 21369 26651 21403
rect 26651 21369 26660 21403
rect 26608 21360 26660 21369
rect 26976 21335 27028 21344
rect 26976 21301 26985 21335
rect 26985 21301 27019 21335
rect 27019 21301 27028 21335
rect 26976 21292 27028 21301
rect 27252 21335 27304 21344
rect 27252 21301 27261 21335
rect 27261 21301 27295 21335
rect 27295 21301 27304 21335
rect 27252 21292 27304 21301
rect 4664 21190 4716 21242
rect 4728 21190 4780 21242
rect 4792 21190 4844 21242
rect 4856 21190 4908 21242
rect 4920 21190 4972 21242
rect 12092 21190 12144 21242
rect 12156 21190 12208 21242
rect 12220 21190 12272 21242
rect 12284 21190 12336 21242
rect 12348 21190 12400 21242
rect 19520 21190 19572 21242
rect 19584 21190 19636 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 26948 21190 27000 21242
rect 27012 21190 27064 21242
rect 27076 21190 27128 21242
rect 27140 21190 27192 21242
rect 27204 21190 27256 21242
rect 5080 21088 5132 21140
rect 6552 21088 6604 21140
rect 8576 21088 8628 21140
rect 9496 21088 9548 21140
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 6092 21020 6144 21072
rect 6828 21020 6880 21072
rect 4160 20884 4212 20936
rect 4252 20884 4304 20936
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5540 20927 5592 20936
rect 5540 20893 5569 20927
rect 5569 20893 5592 20927
rect 7012 20995 7064 21004
rect 7012 20961 7021 20995
rect 7021 20961 7055 20995
rect 7055 20961 7064 20995
rect 7012 20952 7064 20961
rect 5540 20884 5592 20893
rect 6460 20927 6512 20936
rect 6460 20893 6469 20927
rect 6469 20893 6503 20927
rect 6503 20893 6512 20927
rect 6460 20884 6512 20893
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 7564 20995 7616 21004
rect 7564 20961 7573 20995
rect 7573 20961 7607 20995
rect 7607 20961 7616 20995
rect 7564 20952 7616 20961
rect 9680 20952 9732 21004
rect 9956 21088 10008 21140
rect 10508 21131 10560 21140
rect 10508 21097 10517 21131
rect 10517 21097 10551 21131
rect 10551 21097 10560 21131
rect 10508 21088 10560 21097
rect 10784 21088 10836 21140
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 12440 21088 12492 21140
rect 15016 21088 15068 21140
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 6644 20748 6696 20800
rect 6920 20816 6972 20868
rect 7656 20748 7708 20800
rect 8208 20748 8260 20800
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 10416 21020 10468 21072
rect 12624 21063 12676 21072
rect 12624 21029 12633 21063
rect 12633 21029 12667 21063
rect 12667 21029 12676 21063
rect 12624 21020 12676 21029
rect 16396 21088 16448 21140
rect 19432 21131 19484 21140
rect 19432 21097 19441 21131
rect 19441 21097 19475 21131
rect 19475 21097 19484 21131
rect 19432 21088 19484 21097
rect 20352 21088 20404 21140
rect 23112 21088 23164 21140
rect 18696 21063 18748 21072
rect 18696 21029 18705 21063
rect 18705 21029 18739 21063
rect 18739 21029 18748 21063
rect 18696 21020 18748 21029
rect 10968 20952 11020 21004
rect 11520 20884 11572 20936
rect 11796 20927 11848 20936
rect 11796 20893 11805 20927
rect 11805 20893 11839 20927
rect 11839 20893 11848 20927
rect 11796 20884 11848 20893
rect 13084 20884 13136 20936
rect 9312 20816 9364 20868
rect 9588 20748 9640 20800
rect 9680 20791 9732 20800
rect 9680 20757 9705 20791
rect 9705 20757 9732 20791
rect 9864 20816 9916 20868
rect 10140 20816 10192 20868
rect 10968 20859 11020 20868
rect 10968 20825 10977 20859
rect 10977 20825 11011 20859
rect 11011 20825 11020 20859
rect 10968 20816 11020 20825
rect 11060 20859 11112 20868
rect 11060 20825 11069 20859
rect 11069 20825 11103 20859
rect 11103 20825 11112 20859
rect 11060 20816 11112 20825
rect 11152 20859 11204 20868
rect 11152 20825 11187 20859
rect 11187 20825 11204 20859
rect 11152 20816 11204 20825
rect 11612 20859 11664 20868
rect 11612 20825 11621 20859
rect 11621 20825 11655 20859
rect 11655 20825 11664 20859
rect 11612 20816 11664 20825
rect 12440 20816 12492 20868
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 15660 20995 15712 21004
rect 15660 20961 15669 20995
rect 15669 20961 15703 20995
rect 15703 20961 15712 20995
rect 15660 20952 15712 20961
rect 16672 20952 16724 21004
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 15292 20884 15344 20936
rect 14280 20859 14332 20868
rect 14280 20825 14289 20859
rect 14289 20825 14323 20859
rect 14323 20825 14332 20859
rect 14280 20816 14332 20825
rect 15936 20859 15988 20868
rect 15936 20825 15945 20859
rect 15945 20825 15979 20859
rect 15979 20825 15988 20859
rect 15936 20816 15988 20825
rect 16580 20816 16632 20868
rect 18788 20927 18840 20936
rect 18788 20893 18797 20927
rect 18797 20893 18831 20927
rect 18831 20893 18840 20927
rect 18788 20884 18840 20893
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 19340 20884 19392 20936
rect 9680 20748 9732 20757
rect 12072 20748 12124 20800
rect 13728 20748 13780 20800
rect 14188 20748 14240 20800
rect 15016 20748 15068 20800
rect 16764 20748 16816 20800
rect 18972 20816 19024 20868
rect 22284 21063 22336 21072
rect 22284 21029 22293 21063
rect 22293 21029 22327 21063
rect 22327 21029 22336 21063
rect 22284 21020 22336 21029
rect 22836 21020 22888 21072
rect 23020 21063 23072 21072
rect 23020 21029 23029 21063
rect 23029 21029 23063 21063
rect 23063 21029 23072 21063
rect 23020 21020 23072 21029
rect 26700 21088 26752 21140
rect 26792 21088 26844 21140
rect 27528 21088 27580 21140
rect 19616 20952 19668 21004
rect 20720 20995 20772 21004
rect 20720 20961 20729 20995
rect 20729 20961 20763 20995
rect 20763 20961 20772 20995
rect 20720 20952 20772 20961
rect 20812 20952 20864 21004
rect 22192 20884 22244 20936
rect 17960 20748 18012 20800
rect 19892 20748 19944 20800
rect 20996 20816 21048 20868
rect 21916 20859 21968 20868
rect 21916 20825 21925 20859
rect 21925 20825 21959 20859
rect 21959 20825 21968 20859
rect 21916 20816 21968 20825
rect 20076 20748 20128 20800
rect 25504 20952 25556 21004
rect 26608 20952 26660 21004
rect 27160 20952 27212 21004
rect 24124 20816 24176 20868
rect 26792 20927 26844 20936
rect 26792 20893 26801 20927
rect 26801 20893 26835 20927
rect 26835 20893 26844 20927
rect 26792 20884 26844 20893
rect 27160 20816 27212 20868
rect 27988 21020 28040 21072
rect 28632 21020 28684 21072
rect 28448 20884 28500 20936
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 29368 20884 29420 20936
rect 29644 20748 29696 20800
rect 5324 20646 5376 20698
rect 5388 20646 5440 20698
rect 5452 20646 5504 20698
rect 5516 20646 5568 20698
rect 5580 20646 5632 20698
rect 12752 20646 12804 20698
rect 12816 20646 12868 20698
rect 12880 20646 12932 20698
rect 12944 20646 12996 20698
rect 13008 20646 13060 20698
rect 20180 20646 20232 20698
rect 20244 20646 20296 20698
rect 20308 20646 20360 20698
rect 20372 20646 20424 20698
rect 20436 20646 20488 20698
rect 27608 20646 27660 20698
rect 27672 20646 27724 20698
rect 27736 20646 27788 20698
rect 27800 20646 27852 20698
rect 27864 20646 27916 20698
rect 4252 20587 4304 20596
rect 4252 20553 4261 20587
rect 4261 20553 4295 20587
rect 4295 20553 4304 20587
rect 4252 20544 4304 20553
rect 4528 20544 4580 20596
rect 5080 20544 5132 20596
rect 4620 20476 4672 20528
rect 5172 20476 5224 20528
rect 3884 20408 3936 20460
rect 4252 20408 4304 20460
rect 2504 20383 2556 20392
rect 2504 20349 2513 20383
rect 2513 20349 2547 20383
rect 2547 20349 2556 20383
rect 2504 20340 2556 20349
rect 2780 20383 2832 20392
rect 2780 20349 2789 20383
rect 2789 20349 2823 20383
rect 2823 20349 2832 20383
rect 2780 20340 2832 20349
rect 4160 20340 4212 20392
rect 5080 20340 5132 20392
rect 5540 20451 5592 20460
rect 5540 20417 5549 20451
rect 5549 20417 5583 20451
rect 5583 20417 5592 20451
rect 5540 20408 5592 20417
rect 7012 20544 7064 20596
rect 7564 20587 7616 20596
rect 7564 20553 7573 20587
rect 7573 20553 7607 20587
rect 7607 20553 7616 20587
rect 7564 20544 7616 20553
rect 9864 20544 9916 20596
rect 10968 20544 11020 20596
rect 11520 20587 11572 20596
rect 11520 20553 11529 20587
rect 11529 20553 11563 20587
rect 11563 20553 11572 20587
rect 11520 20544 11572 20553
rect 11796 20544 11848 20596
rect 11888 20544 11940 20596
rect 6460 20408 6512 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 8760 20476 8812 20528
rect 11612 20408 11664 20460
rect 11244 20340 11296 20392
rect 11060 20272 11112 20324
rect 4344 20247 4396 20256
rect 4344 20213 4353 20247
rect 4353 20213 4387 20247
rect 4387 20213 4396 20247
rect 4344 20204 4396 20213
rect 5356 20204 5408 20256
rect 8024 20204 8076 20256
rect 12072 20408 12124 20460
rect 12440 20544 12492 20596
rect 13084 20544 13136 20596
rect 13728 20544 13780 20596
rect 12440 20408 12492 20460
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 15660 20544 15712 20596
rect 15936 20544 15988 20596
rect 14464 20476 14516 20528
rect 16028 20476 16080 20528
rect 15568 20408 15620 20460
rect 19984 20544 20036 20596
rect 20720 20544 20772 20596
rect 21824 20544 21876 20596
rect 22100 20544 22152 20596
rect 22836 20587 22888 20596
rect 22836 20553 22845 20587
rect 22845 20553 22879 20587
rect 22879 20553 22888 20587
rect 22836 20544 22888 20553
rect 26792 20544 26844 20596
rect 27344 20544 27396 20596
rect 28632 20544 28684 20596
rect 28816 20544 28868 20596
rect 19340 20476 19392 20528
rect 14280 20340 14332 20392
rect 15200 20272 15252 20324
rect 16764 20408 16816 20460
rect 18880 20408 18932 20460
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 17776 20340 17828 20392
rect 18788 20383 18840 20392
rect 18788 20349 18797 20383
rect 18797 20349 18831 20383
rect 18831 20349 18840 20383
rect 18788 20340 18840 20349
rect 21088 20383 21140 20392
rect 21088 20349 21097 20383
rect 21097 20349 21131 20383
rect 21131 20349 21140 20383
rect 21088 20340 21140 20349
rect 21456 20340 21508 20392
rect 17408 20272 17460 20324
rect 18696 20272 18748 20324
rect 23020 20408 23072 20460
rect 23388 20408 23440 20460
rect 25044 20476 25096 20528
rect 25228 20476 25280 20528
rect 26700 20476 26752 20528
rect 29000 20476 29052 20528
rect 22928 20383 22980 20392
rect 22928 20349 22937 20383
rect 22937 20349 22971 20383
rect 22971 20349 22980 20383
rect 22928 20340 22980 20349
rect 23480 20340 23532 20392
rect 23848 20272 23900 20324
rect 29460 20451 29512 20460
rect 28540 20340 28592 20392
rect 12348 20204 12400 20256
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 13636 20247 13688 20256
rect 13636 20213 13645 20247
rect 13645 20213 13679 20247
rect 13679 20213 13688 20247
rect 13636 20204 13688 20213
rect 14004 20204 14056 20256
rect 19432 20204 19484 20256
rect 22836 20204 22888 20256
rect 24952 20247 25004 20256
rect 24952 20213 24961 20247
rect 24961 20213 24995 20247
rect 24995 20213 25004 20247
rect 24952 20204 25004 20213
rect 28172 20204 28224 20256
rect 29460 20417 29469 20451
rect 29469 20417 29503 20451
rect 29503 20417 29512 20451
rect 29460 20408 29512 20417
rect 29000 20272 29052 20324
rect 29092 20272 29144 20324
rect 28908 20204 28960 20256
rect 30104 20408 30156 20460
rect 29552 20340 29604 20392
rect 30288 20247 30340 20256
rect 30288 20213 30297 20247
rect 30297 20213 30331 20247
rect 30331 20213 30340 20247
rect 30288 20204 30340 20213
rect 4664 20102 4716 20154
rect 4728 20102 4780 20154
rect 4792 20102 4844 20154
rect 4856 20102 4908 20154
rect 4920 20102 4972 20154
rect 12092 20102 12144 20154
rect 12156 20102 12208 20154
rect 12220 20102 12272 20154
rect 12284 20102 12336 20154
rect 12348 20102 12400 20154
rect 19520 20102 19572 20154
rect 19584 20102 19636 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 26948 20102 27000 20154
rect 27012 20102 27064 20154
rect 27076 20102 27128 20154
rect 27140 20102 27192 20154
rect 27204 20102 27256 20154
rect 2780 20000 2832 20052
rect 3884 20043 3936 20052
rect 3884 20009 3893 20043
rect 3893 20009 3927 20043
rect 3927 20009 3936 20043
rect 3884 20000 3936 20009
rect 4344 20000 4396 20052
rect 7932 20000 7984 20052
rect 3700 19796 3752 19848
rect 4988 19864 5040 19916
rect 5356 19864 5408 19916
rect 7380 19864 7432 19916
rect 940 19660 992 19712
rect 4712 19703 4764 19712
rect 4712 19669 4721 19703
rect 4721 19669 4755 19703
rect 4755 19669 4764 19703
rect 4712 19660 4764 19669
rect 4896 19660 4948 19712
rect 5540 19796 5592 19848
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 7472 19660 7524 19712
rect 8024 19796 8076 19848
rect 7840 19771 7892 19780
rect 7840 19737 7849 19771
rect 7849 19737 7883 19771
rect 7883 19737 7892 19771
rect 7840 19728 7892 19737
rect 9036 19796 9088 19848
rect 9312 19864 9364 19916
rect 9772 19864 9824 19916
rect 10324 19864 10376 19916
rect 11152 20043 11204 20052
rect 11152 20009 11161 20043
rect 11161 20009 11195 20043
rect 11195 20009 11204 20043
rect 11152 20000 11204 20009
rect 11060 19975 11112 19984
rect 11060 19941 11069 19975
rect 11069 19941 11103 19975
rect 11103 19941 11112 19975
rect 11060 19932 11112 19941
rect 12532 20000 12584 20052
rect 13360 20000 13412 20052
rect 11612 19907 11664 19916
rect 11612 19873 11621 19907
rect 11621 19873 11655 19907
rect 11655 19873 11664 19907
rect 11612 19864 11664 19873
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 13912 19932 13964 19984
rect 17316 20000 17368 20052
rect 17868 20000 17920 20052
rect 19340 20043 19392 20052
rect 19340 20009 19349 20043
rect 19349 20009 19383 20043
rect 19383 20009 19392 20043
rect 19340 20000 19392 20009
rect 20076 20000 20128 20052
rect 24124 20000 24176 20052
rect 17684 19932 17736 19984
rect 10140 19728 10192 19780
rect 12624 19796 12676 19848
rect 12716 19839 12768 19848
rect 12716 19805 12725 19839
rect 12725 19805 12759 19839
rect 12759 19805 12768 19839
rect 12716 19796 12768 19805
rect 17040 19864 17092 19916
rect 19156 19864 19208 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 21180 19907 21232 19916
rect 21180 19873 21189 19907
rect 21189 19873 21223 19907
rect 21223 19873 21232 19907
rect 21180 19864 21232 19873
rect 22928 19907 22980 19916
rect 22928 19873 22937 19907
rect 22937 19873 22971 19907
rect 22971 19873 22980 19907
rect 22928 19864 22980 19873
rect 27620 20000 27672 20052
rect 11612 19660 11664 19712
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 17500 19796 17552 19848
rect 18604 19839 18656 19848
rect 18604 19805 18613 19839
rect 18613 19805 18647 19839
rect 18647 19805 18656 19839
rect 18604 19796 18656 19805
rect 17224 19728 17276 19780
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 20076 19796 20128 19848
rect 20536 19796 20588 19848
rect 20720 19796 20772 19848
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 16028 19660 16080 19712
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 18880 19660 18932 19712
rect 23020 19728 23072 19780
rect 23388 19796 23440 19848
rect 25412 19932 25464 19984
rect 28172 20043 28224 20052
rect 28172 20009 28181 20043
rect 28181 20009 28215 20043
rect 28215 20009 28224 20043
rect 28172 20000 28224 20009
rect 28264 20000 28316 20052
rect 29460 20000 29512 20052
rect 30288 20000 30340 20052
rect 29092 19975 29144 19984
rect 29092 19941 29101 19975
rect 29101 19941 29135 19975
rect 29135 19941 29144 19975
rect 29092 19932 29144 19941
rect 25780 19864 25832 19916
rect 27988 19864 28040 19916
rect 28908 19907 28960 19916
rect 28908 19873 28917 19907
rect 28917 19873 28951 19907
rect 28951 19873 28960 19907
rect 28908 19864 28960 19873
rect 29276 19864 29328 19916
rect 24216 19728 24268 19780
rect 28632 19728 28684 19780
rect 29276 19728 29328 19780
rect 23480 19660 23532 19712
rect 24492 19703 24544 19712
rect 24492 19669 24501 19703
rect 24501 19669 24535 19703
rect 24535 19669 24544 19703
rect 24492 19660 24544 19669
rect 25228 19703 25280 19712
rect 25228 19669 25237 19703
rect 25237 19669 25271 19703
rect 25271 19669 25280 19703
rect 25228 19660 25280 19669
rect 29092 19660 29144 19712
rect 29644 19660 29696 19712
rect 5324 19558 5376 19610
rect 5388 19558 5440 19610
rect 5452 19558 5504 19610
rect 5516 19558 5568 19610
rect 5580 19558 5632 19610
rect 12752 19558 12804 19610
rect 12816 19558 12868 19610
rect 12880 19558 12932 19610
rect 12944 19558 12996 19610
rect 13008 19558 13060 19610
rect 20180 19558 20232 19610
rect 20244 19558 20296 19610
rect 20308 19558 20360 19610
rect 20372 19558 20424 19610
rect 20436 19558 20488 19610
rect 27608 19558 27660 19610
rect 27672 19558 27724 19610
rect 27736 19558 27788 19610
rect 27800 19558 27852 19610
rect 27864 19558 27916 19610
rect 4712 19456 4764 19508
rect 6460 19456 6512 19508
rect 6828 19456 6880 19508
rect 8484 19456 8536 19508
rect 9496 19456 9548 19508
rect 10232 19456 10284 19508
rect 10416 19456 10468 19508
rect 7932 19388 7984 19440
rect 8576 19388 8628 19440
rect 9128 19388 9180 19440
rect 7564 19363 7616 19372
rect 7564 19329 7573 19363
rect 7573 19329 7607 19363
rect 7607 19329 7616 19363
rect 7564 19320 7616 19329
rect 4988 19295 5040 19304
rect 4988 19261 4997 19295
rect 4997 19261 5031 19295
rect 5031 19261 5040 19295
rect 4988 19252 5040 19261
rect 4528 19184 4580 19236
rect 5080 19184 5132 19236
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 9772 19252 9824 19304
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 5540 19159 5592 19168
rect 5540 19125 5549 19159
rect 5549 19125 5583 19159
rect 5583 19125 5592 19159
rect 5540 19116 5592 19125
rect 12624 19184 12676 19236
rect 13636 19184 13688 19236
rect 13912 19320 13964 19372
rect 14096 19184 14148 19236
rect 16028 19456 16080 19508
rect 14464 19431 14516 19440
rect 14464 19397 14473 19431
rect 14473 19397 14507 19431
rect 14507 19397 14516 19431
rect 14464 19388 14516 19397
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 16764 19456 16816 19508
rect 17408 19499 17460 19508
rect 17408 19465 17417 19499
rect 17417 19465 17451 19499
rect 17451 19465 17460 19499
rect 17408 19456 17460 19465
rect 18420 19456 18472 19508
rect 18696 19456 18748 19508
rect 18788 19456 18840 19508
rect 19432 19499 19484 19508
rect 19432 19465 19441 19499
rect 19441 19465 19475 19499
rect 19475 19465 19484 19499
rect 19432 19456 19484 19465
rect 20076 19456 20128 19508
rect 21916 19456 21968 19508
rect 16948 19363 17000 19372
rect 16948 19329 16965 19363
rect 16965 19329 17000 19363
rect 16948 19320 17000 19329
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 17684 19320 17736 19372
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 20536 19388 20588 19440
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18144 19320 18196 19329
rect 18604 19320 18656 19372
rect 18880 19320 18932 19372
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 19156 19320 19208 19372
rect 19340 19320 19392 19372
rect 17592 19252 17644 19304
rect 17776 19252 17828 19304
rect 14832 19184 14884 19236
rect 17224 19184 17276 19236
rect 13360 19159 13412 19168
rect 13360 19125 13369 19159
rect 13369 19125 13403 19159
rect 13403 19125 13412 19159
rect 13360 19116 13412 19125
rect 13820 19116 13872 19168
rect 20812 19320 20864 19372
rect 23388 19388 23440 19440
rect 20720 19252 20772 19304
rect 18144 19116 18196 19168
rect 18880 19116 18932 19168
rect 21180 19295 21232 19304
rect 21180 19261 21189 19295
rect 21189 19261 21223 19295
rect 21223 19261 21232 19295
rect 21180 19252 21232 19261
rect 21916 19320 21968 19372
rect 23020 19363 23072 19372
rect 23020 19329 23029 19363
rect 23029 19329 23063 19363
rect 23063 19329 23072 19363
rect 23020 19320 23072 19329
rect 23480 19363 23532 19372
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 22928 19252 22980 19304
rect 24216 19388 24268 19440
rect 24492 19456 24544 19508
rect 25228 19456 25280 19508
rect 24952 19388 25004 19440
rect 25780 19388 25832 19440
rect 23940 19320 23992 19372
rect 26792 19456 26844 19508
rect 26516 19431 26568 19440
rect 26516 19397 26525 19431
rect 26525 19397 26559 19431
rect 26559 19397 26568 19431
rect 26516 19388 26568 19397
rect 30288 19456 30340 19508
rect 26332 19363 26384 19372
rect 26332 19329 26341 19363
rect 26341 19329 26375 19363
rect 26375 19329 26384 19363
rect 26332 19320 26384 19329
rect 26424 19363 26476 19372
rect 26424 19329 26433 19363
rect 26433 19329 26467 19363
rect 26467 19329 26476 19363
rect 26424 19320 26476 19329
rect 27988 19320 28040 19372
rect 26240 19252 26292 19304
rect 26884 19252 26936 19304
rect 29368 19363 29420 19372
rect 29368 19329 29377 19363
rect 29377 19329 29411 19363
rect 29411 19329 29420 19363
rect 29368 19320 29420 19329
rect 30104 19363 30156 19372
rect 30104 19329 30113 19363
rect 30113 19329 30147 19363
rect 30147 19329 30156 19363
rect 30104 19320 30156 19329
rect 20904 19116 20956 19168
rect 23296 19116 23348 19168
rect 27344 19116 27396 19168
rect 27896 19116 27948 19168
rect 28264 19116 28316 19168
rect 28816 19116 28868 19168
rect 28908 19159 28960 19168
rect 28908 19125 28917 19159
rect 28917 19125 28951 19159
rect 28951 19125 28960 19159
rect 28908 19116 28960 19125
rect 29276 19184 29328 19236
rect 29184 19116 29236 19168
rect 4664 19014 4716 19066
rect 4728 19014 4780 19066
rect 4792 19014 4844 19066
rect 4856 19014 4908 19066
rect 4920 19014 4972 19066
rect 12092 19014 12144 19066
rect 12156 19014 12208 19066
rect 12220 19014 12272 19066
rect 12284 19014 12336 19066
rect 12348 19014 12400 19066
rect 19520 19014 19572 19066
rect 19584 19014 19636 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 26948 19014 27000 19066
rect 27012 19014 27064 19066
rect 27076 19014 27128 19066
rect 27140 19014 27192 19066
rect 27204 19014 27256 19066
rect 7380 18912 7432 18964
rect 7472 18912 7524 18964
rect 8576 18912 8628 18964
rect 9864 18912 9916 18964
rect 13820 18912 13872 18964
rect 13912 18955 13964 18964
rect 13912 18921 13921 18955
rect 13921 18921 13955 18955
rect 13955 18921 13964 18955
rect 13912 18912 13964 18921
rect 16764 18912 16816 18964
rect 17316 18955 17368 18964
rect 17316 18921 17325 18955
rect 17325 18921 17359 18955
rect 17359 18921 17368 18955
rect 17316 18912 17368 18921
rect 17592 18955 17644 18964
rect 17592 18921 17601 18955
rect 17601 18921 17635 18955
rect 17635 18921 17644 18955
rect 17592 18912 17644 18921
rect 18328 18912 18380 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 19156 18912 19208 18964
rect 26332 18912 26384 18964
rect 4528 18819 4580 18828
rect 4528 18785 4537 18819
rect 4537 18785 4571 18819
rect 4571 18785 4580 18819
rect 4528 18776 4580 18785
rect 3700 18708 3752 18760
rect 3792 18708 3844 18760
rect 7564 18776 7616 18828
rect 9496 18776 9548 18828
rect 7656 18708 7708 18760
rect 940 18572 992 18624
rect 3148 18615 3200 18624
rect 3148 18581 3157 18615
rect 3157 18581 3191 18615
rect 3191 18581 3200 18615
rect 3148 18572 3200 18581
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 4436 18640 4488 18692
rect 4344 18615 4396 18624
rect 4344 18581 4353 18615
rect 4353 18581 4387 18615
rect 4387 18581 4396 18615
rect 4344 18572 4396 18581
rect 4896 18572 4948 18624
rect 6092 18640 6144 18692
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 5540 18572 5592 18624
rect 11704 18572 11756 18624
rect 15108 18708 15160 18760
rect 15384 18708 15436 18760
rect 18144 18844 18196 18896
rect 18972 18887 19024 18896
rect 18972 18853 18981 18887
rect 18981 18853 19015 18887
rect 19015 18853 19024 18887
rect 18972 18844 19024 18853
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 16212 18708 16264 18760
rect 17040 18708 17092 18760
rect 17316 18708 17368 18760
rect 17500 18708 17552 18760
rect 17592 18708 17644 18760
rect 19248 18776 19300 18828
rect 23848 18844 23900 18896
rect 28080 18912 28132 18964
rect 29276 18887 29328 18896
rect 22928 18776 22980 18828
rect 26516 18776 26568 18828
rect 16856 18572 16908 18624
rect 18972 18708 19024 18760
rect 19892 18708 19944 18760
rect 23020 18751 23072 18760
rect 23020 18717 23029 18751
rect 23029 18717 23063 18751
rect 23063 18717 23072 18751
rect 23020 18708 23072 18717
rect 20904 18640 20956 18692
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 24584 18751 24636 18760
rect 24584 18717 24593 18751
rect 24593 18717 24627 18751
rect 24627 18717 24636 18751
rect 24584 18708 24636 18717
rect 27436 18751 27488 18760
rect 27436 18717 27445 18751
rect 27445 18717 27479 18751
rect 27479 18717 27488 18751
rect 27436 18708 27488 18717
rect 29276 18853 29285 18887
rect 29285 18853 29319 18887
rect 29319 18853 29328 18887
rect 29276 18844 29328 18853
rect 23388 18640 23440 18692
rect 28172 18751 28224 18760
rect 28172 18717 28181 18751
rect 28181 18717 28215 18751
rect 28215 18717 28224 18751
rect 28172 18708 28224 18717
rect 28448 18708 28500 18760
rect 28816 18640 28868 18692
rect 29184 18640 29236 18692
rect 24400 18615 24452 18624
rect 24400 18581 24409 18615
rect 24409 18581 24443 18615
rect 24443 18581 24452 18615
rect 24400 18572 24452 18581
rect 25964 18572 26016 18624
rect 26240 18572 26292 18624
rect 28264 18572 28316 18624
rect 28356 18572 28408 18624
rect 5324 18470 5376 18522
rect 5388 18470 5440 18522
rect 5452 18470 5504 18522
rect 5516 18470 5568 18522
rect 5580 18470 5632 18522
rect 12752 18470 12804 18522
rect 12816 18470 12868 18522
rect 12880 18470 12932 18522
rect 12944 18470 12996 18522
rect 13008 18470 13060 18522
rect 20180 18470 20232 18522
rect 20244 18470 20296 18522
rect 20308 18470 20360 18522
rect 20372 18470 20424 18522
rect 20436 18470 20488 18522
rect 27608 18470 27660 18522
rect 27672 18470 27724 18522
rect 27736 18470 27788 18522
rect 27800 18470 27852 18522
rect 27864 18470 27916 18522
rect 3148 18368 3200 18420
rect 3700 18368 3752 18420
rect 3516 18300 3568 18352
rect 4988 18368 5040 18420
rect 6092 18411 6144 18420
rect 6092 18377 6101 18411
rect 6101 18377 6135 18411
rect 6135 18377 6144 18411
rect 6092 18368 6144 18377
rect 7656 18368 7708 18420
rect 2504 18232 2556 18284
rect 7196 18232 7248 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 11428 18368 11480 18420
rect 11888 18368 11940 18420
rect 13360 18368 13412 18420
rect 14280 18368 14332 18420
rect 6736 18207 6788 18216
rect 6736 18173 6745 18207
rect 6745 18173 6779 18207
rect 6779 18173 6788 18207
rect 6736 18164 6788 18173
rect 7012 18096 7064 18148
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 9772 18096 9824 18148
rect 9864 18096 9916 18148
rect 3700 18028 3752 18080
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 9588 18028 9640 18080
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 11428 18232 11480 18284
rect 12072 18300 12124 18352
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 18880 18368 18932 18420
rect 24400 18368 24452 18420
rect 24584 18368 24636 18420
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 10140 18096 10192 18148
rect 10600 18096 10652 18148
rect 12624 18164 12676 18216
rect 13452 18164 13504 18216
rect 14464 18207 14516 18216
rect 14464 18173 14473 18207
rect 14473 18173 14507 18207
rect 14507 18173 14516 18207
rect 14464 18164 14516 18173
rect 14832 18232 14884 18284
rect 15016 18096 15068 18148
rect 17224 18232 17276 18284
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 17592 18164 17644 18216
rect 17776 18096 17828 18148
rect 20536 18232 20588 18284
rect 20076 18164 20128 18216
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 20996 18232 21048 18284
rect 24860 18300 24912 18352
rect 22928 18232 22980 18284
rect 23020 18232 23072 18284
rect 23388 18232 23440 18284
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 26148 18275 26200 18284
rect 25412 18164 25464 18216
rect 26148 18241 26157 18275
rect 26157 18241 26191 18275
rect 26191 18241 26200 18275
rect 26148 18232 26200 18241
rect 26792 18232 26844 18284
rect 27344 18300 27396 18352
rect 27988 18300 28040 18352
rect 28172 18300 28224 18352
rect 28448 18411 28500 18420
rect 28448 18377 28457 18411
rect 28457 18377 28491 18411
rect 28491 18377 28500 18411
rect 28448 18368 28500 18377
rect 29184 18411 29236 18420
rect 29184 18377 29193 18411
rect 29193 18377 29227 18411
rect 29227 18377 29236 18411
rect 29184 18368 29236 18377
rect 28632 18300 28684 18352
rect 30104 18300 30156 18352
rect 29184 18275 29236 18284
rect 29184 18241 29193 18275
rect 29193 18241 29227 18275
rect 29227 18241 29236 18275
rect 29184 18232 29236 18241
rect 30012 18232 30064 18284
rect 26056 18164 26108 18216
rect 11060 18028 11112 18080
rect 11888 18028 11940 18080
rect 14096 18028 14148 18080
rect 16580 18028 16632 18080
rect 17960 18028 18012 18080
rect 19248 18028 19300 18080
rect 19432 18028 19484 18080
rect 20628 18028 20680 18080
rect 23480 18028 23532 18080
rect 27528 18028 27580 18080
rect 28080 18028 28132 18080
rect 4664 17926 4716 17978
rect 4728 17926 4780 17978
rect 4792 17926 4844 17978
rect 4856 17926 4908 17978
rect 4920 17926 4972 17978
rect 12092 17926 12144 17978
rect 12156 17926 12208 17978
rect 12220 17926 12272 17978
rect 12284 17926 12336 17978
rect 12348 17926 12400 17978
rect 19520 17926 19572 17978
rect 19584 17926 19636 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 26948 17926 27000 17978
rect 27012 17926 27064 17978
rect 27076 17926 27128 17978
rect 27140 17926 27192 17978
rect 27204 17926 27256 17978
rect 6460 17824 6512 17876
rect 3792 17663 3844 17672
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 5724 17620 5776 17672
rect 6736 17824 6788 17876
rect 8300 17824 8352 17876
rect 9864 17824 9916 17876
rect 10508 17867 10560 17876
rect 10508 17833 10517 17867
rect 10517 17833 10551 17867
rect 10551 17833 10560 17867
rect 10508 17824 10560 17833
rect 11060 17867 11112 17876
rect 11060 17833 11069 17867
rect 11069 17833 11103 17867
rect 11103 17833 11112 17867
rect 11060 17824 11112 17833
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 6920 17756 6972 17808
rect 7288 17756 7340 17808
rect 12348 17756 12400 17808
rect 4068 17595 4120 17604
rect 4068 17561 4077 17595
rect 4077 17561 4111 17595
rect 4111 17561 4120 17595
rect 4068 17552 4120 17561
rect 4528 17552 4580 17604
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 7196 17552 7248 17604
rect 6460 17484 6512 17536
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 8208 17663 8260 17672
rect 8208 17629 8217 17663
rect 8217 17629 8251 17663
rect 8251 17629 8260 17663
rect 8208 17620 8260 17629
rect 8852 17688 8904 17740
rect 10048 17688 10100 17740
rect 8668 17620 8720 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9772 17620 9824 17672
rect 10140 17620 10192 17672
rect 8484 17552 8536 17604
rect 8668 17484 8720 17536
rect 11060 17552 11112 17604
rect 12072 17620 12124 17672
rect 14740 17620 14792 17672
rect 17960 17799 18012 17808
rect 17960 17765 17969 17799
rect 17969 17765 18003 17799
rect 18003 17765 18012 17799
rect 17960 17756 18012 17765
rect 18972 17824 19024 17876
rect 19156 17824 19208 17876
rect 19892 17824 19944 17876
rect 20168 17756 20220 17808
rect 15660 17688 15712 17740
rect 16580 17688 16632 17740
rect 12624 17595 12676 17604
rect 12624 17561 12633 17595
rect 12633 17561 12667 17595
rect 12667 17561 12676 17595
rect 12624 17552 12676 17561
rect 17040 17552 17092 17604
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 27436 17824 27488 17876
rect 27620 17824 27672 17876
rect 28172 17824 28224 17876
rect 29184 17867 29236 17876
rect 29184 17833 29193 17867
rect 29193 17833 29227 17867
rect 29227 17833 29236 17867
rect 29184 17824 29236 17833
rect 22928 17688 22980 17740
rect 27344 17731 27396 17740
rect 27344 17697 27353 17731
rect 27353 17697 27387 17731
rect 27387 17697 27396 17731
rect 27344 17688 27396 17697
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 23020 17663 23072 17672
rect 23020 17629 23029 17663
rect 23029 17629 23063 17663
rect 23063 17629 23072 17663
rect 23020 17620 23072 17629
rect 23572 17663 23624 17672
rect 23572 17629 23581 17663
rect 23581 17629 23615 17663
rect 23615 17629 23624 17663
rect 23572 17620 23624 17629
rect 25044 17620 25096 17672
rect 27988 17663 28040 17672
rect 23388 17552 23440 17604
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28080 17552 28132 17604
rect 30012 17867 30064 17876
rect 30012 17833 30021 17867
rect 30021 17833 30055 17867
rect 30055 17833 30064 17867
rect 30012 17824 30064 17833
rect 11888 17484 11940 17536
rect 19340 17484 19392 17536
rect 19892 17484 19944 17536
rect 20168 17484 20220 17536
rect 24032 17484 24084 17536
rect 26148 17484 26200 17536
rect 5324 17382 5376 17434
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 12752 17382 12804 17434
rect 12816 17382 12868 17434
rect 12880 17382 12932 17434
rect 12944 17382 12996 17434
rect 13008 17382 13060 17434
rect 20180 17382 20232 17434
rect 20244 17382 20296 17434
rect 20308 17382 20360 17434
rect 20372 17382 20424 17434
rect 20436 17382 20488 17434
rect 27608 17382 27660 17434
rect 27672 17382 27724 17434
rect 27736 17382 27788 17434
rect 27800 17382 27852 17434
rect 27864 17382 27916 17434
rect 4068 17280 4120 17332
rect 4528 17323 4580 17332
rect 4528 17289 4537 17323
rect 4537 17289 4571 17323
rect 4571 17289 4580 17323
rect 4528 17280 4580 17289
rect 5724 17280 5776 17332
rect 6828 17323 6880 17332
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7840 17280 7892 17332
rect 9588 17280 9640 17332
rect 12624 17280 12676 17332
rect 14832 17280 14884 17332
rect 7932 17212 7984 17264
rect 13728 17212 13780 17264
rect 14556 17212 14608 17264
rect 4068 17076 4120 17128
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 6920 17144 6972 17196
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 9680 17144 9732 17196
rect 11060 17144 11112 17196
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 6276 17076 6328 17128
rect 4344 17008 4396 17060
rect 8116 17076 8168 17128
rect 12072 17144 12124 17196
rect 11980 17076 12032 17128
rect 12348 17187 12400 17196
rect 12348 17153 12357 17187
rect 12357 17153 12391 17187
rect 12391 17153 12400 17187
rect 12348 17144 12400 17153
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 13452 17187 13504 17196
rect 13452 17153 13461 17187
rect 13461 17153 13495 17187
rect 13495 17153 13504 17187
rect 13452 17144 13504 17153
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 13820 17119 13872 17128
rect 13820 17085 13829 17119
rect 13829 17085 13863 17119
rect 13863 17085 13872 17119
rect 13820 17076 13872 17085
rect 15568 17144 15620 17196
rect 15844 17144 15896 17196
rect 16856 17280 16908 17332
rect 17040 17323 17092 17332
rect 17040 17289 17049 17323
rect 17049 17289 17083 17323
rect 17083 17289 17092 17323
rect 17040 17280 17092 17289
rect 17224 17323 17276 17332
rect 17224 17289 17233 17323
rect 17233 17289 17267 17323
rect 17267 17289 17276 17323
rect 17224 17280 17276 17289
rect 17868 17280 17920 17332
rect 17960 17280 18012 17332
rect 19340 17280 19392 17332
rect 21088 17280 21140 17332
rect 19892 17212 19944 17264
rect 23480 17255 23532 17264
rect 23480 17221 23489 17255
rect 23489 17221 23523 17255
rect 23523 17221 23532 17255
rect 23480 17212 23532 17221
rect 24952 17280 25004 17332
rect 26424 17280 26476 17332
rect 18328 17144 18380 17196
rect 20076 17187 20128 17196
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 20904 17144 20956 17196
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 23664 17187 23716 17196
rect 23664 17153 23673 17187
rect 23673 17153 23707 17187
rect 23707 17153 23716 17187
rect 23664 17144 23716 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 25136 17144 25188 17196
rect 27528 17187 27580 17196
rect 27528 17153 27537 17187
rect 27537 17153 27571 17187
rect 27571 17153 27580 17187
rect 27528 17144 27580 17153
rect 28172 17144 28224 17196
rect 6460 16983 6512 16992
rect 6460 16949 6469 16983
rect 6469 16949 6503 16983
rect 6503 16949 6512 16983
rect 6460 16940 6512 16949
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 7380 16940 7432 16992
rect 9036 16940 9088 16992
rect 11244 16940 11296 16992
rect 12256 16940 12308 16992
rect 18328 17008 18380 17060
rect 23204 17008 23256 17060
rect 28264 17076 28316 17128
rect 13268 16940 13320 16992
rect 14004 16940 14056 16992
rect 17040 16940 17092 16992
rect 19892 16940 19944 16992
rect 23020 16940 23072 16992
rect 23112 16940 23164 16992
rect 27804 17008 27856 17060
rect 28080 16940 28132 16992
rect 4664 16838 4716 16890
rect 4728 16838 4780 16890
rect 4792 16838 4844 16890
rect 4856 16838 4908 16890
rect 4920 16838 4972 16890
rect 12092 16838 12144 16890
rect 12156 16838 12208 16890
rect 12220 16838 12272 16890
rect 12284 16838 12336 16890
rect 12348 16838 12400 16890
rect 19520 16838 19572 16890
rect 19584 16838 19636 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 26948 16838 27000 16890
rect 27012 16838 27064 16890
rect 27076 16838 27128 16890
rect 27140 16838 27192 16890
rect 27204 16838 27256 16890
rect 5264 16736 5316 16788
rect 8116 16736 8168 16788
rect 5724 16668 5776 16720
rect 6184 16668 6236 16720
rect 6276 16668 6328 16720
rect 9588 16736 9640 16788
rect 9680 16736 9732 16788
rect 10508 16736 10560 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 13820 16736 13872 16788
rect 14556 16736 14608 16788
rect 15200 16736 15252 16788
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 18420 16736 18472 16788
rect 18880 16736 18932 16788
rect 19892 16736 19944 16788
rect 20536 16736 20588 16788
rect 21088 16736 21140 16788
rect 11796 16668 11848 16720
rect 4528 16600 4580 16652
rect 5264 16600 5316 16652
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 9496 16600 9548 16652
rect 9588 16600 9640 16652
rect 8576 16532 8628 16584
rect 9036 16532 9088 16584
rect 9128 16532 9180 16584
rect 11152 16600 11204 16652
rect 5172 16464 5224 16516
rect 2688 16396 2740 16448
rect 4160 16439 4212 16448
rect 4160 16405 4169 16439
rect 4169 16405 4203 16439
rect 4203 16405 4212 16439
rect 4160 16396 4212 16405
rect 6552 16396 6604 16448
rect 8392 16464 8444 16516
rect 8116 16396 8168 16448
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 13268 16600 13320 16652
rect 17960 16668 18012 16720
rect 19156 16668 19208 16720
rect 20076 16668 20128 16720
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 15568 16600 15620 16652
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15844 16532 15896 16584
rect 18788 16532 18840 16584
rect 19984 16600 20036 16652
rect 20996 16600 21048 16652
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 26792 16736 26844 16788
rect 27988 16736 28040 16788
rect 23020 16668 23072 16720
rect 23756 16668 23808 16720
rect 11980 16464 12032 16516
rect 18144 16507 18196 16516
rect 18144 16473 18153 16507
rect 18153 16473 18187 16507
rect 18187 16473 18196 16507
rect 18144 16464 18196 16473
rect 18512 16464 18564 16516
rect 11888 16396 11940 16448
rect 13452 16396 13504 16448
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 18880 16464 18932 16516
rect 23112 16532 23164 16584
rect 23664 16532 23716 16584
rect 20628 16507 20680 16516
rect 20628 16473 20637 16507
rect 20637 16473 20671 16507
rect 20671 16473 20680 16507
rect 20628 16464 20680 16473
rect 21088 16464 21140 16516
rect 22008 16464 22060 16516
rect 24860 16600 24912 16652
rect 27436 16600 27488 16652
rect 21824 16396 21876 16448
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 23480 16439 23532 16448
rect 23480 16405 23489 16439
rect 23489 16405 23523 16439
rect 23523 16405 23532 16439
rect 23480 16396 23532 16405
rect 23940 16439 23992 16448
rect 23940 16405 23949 16439
rect 23949 16405 23983 16439
rect 23983 16405 23992 16439
rect 23940 16396 23992 16405
rect 25412 16464 25464 16516
rect 26148 16464 26200 16516
rect 26516 16507 26568 16516
rect 26516 16473 26525 16507
rect 26525 16473 26559 16507
rect 26559 16473 26568 16507
rect 26516 16464 26568 16473
rect 27528 16464 27580 16516
rect 28264 16507 28316 16516
rect 28264 16473 28273 16507
rect 28273 16473 28307 16507
rect 28307 16473 28316 16507
rect 28264 16464 28316 16473
rect 26240 16439 26292 16448
rect 26240 16405 26249 16439
rect 26249 16405 26283 16439
rect 26283 16405 26292 16439
rect 26240 16396 26292 16405
rect 30380 16464 30432 16516
rect 5324 16294 5376 16346
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 12752 16294 12804 16346
rect 12816 16294 12868 16346
rect 12880 16294 12932 16346
rect 12944 16294 12996 16346
rect 13008 16294 13060 16346
rect 20180 16294 20232 16346
rect 20244 16294 20296 16346
rect 20308 16294 20360 16346
rect 20372 16294 20424 16346
rect 20436 16294 20488 16346
rect 27608 16294 27660 16346
rect 27672 16294 27724 16346
rect 27736 16294 27788 16346
rect 27800 16294 27852 16346
rect 27864 16294 27916 16346
rect 4160 16192 4212 16244
rect 6920 16192 6972 16244
rect 3976 16124 4028 16176
rect 8300 16167 8352 16176
rect 8300 16133 8309 16167
rect 8309 16133 8343 16167
rect 8343 16133 8352 16167
rect 8300 16124 8352 16133
rect 8668 16192 8720 16244
rect 9404 16192 9456 16244
rect 18236 16192 18288 16244
rect 13544 16124 13596 16176
rect 1860 15988 1912 16040
rect 2320 16031 2372 16040
rect 2320 15997 2329 16031
rect 2329 15997 2363 16031
rect 2363 15997 2372 16031
rect 2320 15988 2372 15997
rect 3608 16056 3660 16108
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 4344 16056 4396 16108
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 5172 16056 5224 16108
rect 5724 16056 5776 16108
rect 6000 16099 6052 16108
rect 6000 16065 6009 16099
rect 6009 16065 6043 16099
rect 6043 16065 6052 16099
rect 6000 16056 6052 16065
rect 1676 15852 1728 15904
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 6736 16099 6788 16108
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 8116 16099 8168 16108
rect 8116 16065 8125 16099
rect 8125 16065 8159 16099
rect 8159 16065 8168 16099
rect 8116 16056 8168 16065
rect 6368 15988 6420 16040
rect 8392 16099 8444 16108
rect 8392 16065 8427 16099
rect 8427 16065 8444 16099
rect 8392 16056 8444 16065
rect 8576 16099 8628 16108
rect 8576 16065 8585 16099
rect 8585 16065 8619 16099
rect 8619 16065 8628 16099
rect 8576 16056 8628 16065
rect 8852 16056 8904 16108
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 11060 16056 11112 16108
rect 13268 16056 13320 16108
rect 13912 16056 13964 16108
rect 14372 16124 14424 16176
rect 16856 16124 16908 16176
rect 17040 16124 17092 16176
rect 18144 16124 18196 16176
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 19340 16192 19392 16244
rect 23204 16235 23256 16244
rect 23204 16201 23213 16235
rect 23213 16201 23247 16235
rect 23247 16201 23256 16235
rect 23204 16192 23256 16201
rect 24860 16192 24912 16244
rect 25136 16192 25188 16244
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 18696 16124 18748 16176
rect 15844 16056 15896 16108
rect 4988 15852 5040 15904
rect 6184 15852 6236 15904
rect 7472 15852 7524 15904
rect 9404 15988 9456 16040
rect 11704 15988 11756 16040
rect 13544 15988 13596 16040
rect 13728 15988 13780 16040
rect 14832 15988 14884 16040
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 20536 16056 20588 16108
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 18604 15988 18656 16040
rect 18788 15988 18840 16040
rect 23480 16056 23532 16108
rect 23572 16056 23624 16108
rect 25044 16056 25096 16108
rect 25320 16099 25372 16108
rect 25320 16065 25329 16099
rect 25329 16065 25363 16099
rect 25363 16065 25372 16099
rect 25320 16056 25372 16065
rect 22100 15988 22152 16040
rect 27436 16124 27488 16176
rect 26240 16056 26292 16108
rect 26700 16056 26752 16108
rect 26792 16056 26844 16108
rect 27620 16056 27672 16108
rect 27988 16056 28040 16108
rect 26056 16031 26108 16040
rect 26056 15997 26065 16031
rect 26065 15997 26099 16031
rect 26099 15997 26108 16031
rect 26056 15988 26108 15997
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 19432 15920 19484 15972
rect 21916 15920 21968 15972
rect 13084 15852 13136 15904
rect 14188 15852 14240 15904
rect 15660 15852 15712 15904
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 17040 15852 17092 15861
rect 18604 15895 18656 15904
rect 18604 15861 18621 15895
rect 18621 15861 18655 15895
rect 18655 15861 18656 15895
rect 18604 15852 18656 15861
rect 20168 15895 20220 15904
rect 20168 15861 20177 15895
rect 20177 15861 20211 15895
rect 20211 15861 20220 15895
rect 20168 15852 20220 15861
rect 21640 15895 21692 15904
rect 21640 15861 21649 15895
rect 21649 15861 21683 15895
rect 21683 15861 21692 15895
rect 21640 15852 21692 15861
rect 23296 15852 23348 15904
rect 26332 15852 26384 15904
rect 27620 15920 27672 15972
rect 28172 15895 28224 15904
rect 28172 15861 28181 15895
rect 28181 15861 28215 15895
rect 28215 15861 28224 15895
rect 28172 15852 28224 15861
rect 4664 15750 4716 15802
rect 4728 15750 4780 15802
rect 4792 15750 4844 15802
rect 4856 15750 4908 15802
rect 4920 15750 4972 15802
rect 12092 15750 12144 15802
rect 12156 15750 12208 15802
rect 12220 15750 12272 15802
rect 12284 15750 12336 15802
rect 12348 15750 12400 15802
rect 19520 15750 19572 15802
rect 19584 15750 19636 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 26948 15750 27000 15802
rect 27012 15750 27064 15802
rect 27076 15750 27128 15802
rect 27140 15750 27192 15802
rect 27204 15750 27256 15802
rect 2320 15648 2372 15700
rect 6000 15648 6052 15700
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 8484 15648 8536 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 11244 15648 11296 15700
rect 11980 15648 12032 15700
rect 13636 15648 13688 15700
rect 13728 15648 13780 15700
rect 13360 15580 13412 15632
rect 4344 15512 4396 15564
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 5172 15512 5224 15564
rect 6092 15512 6144 15564
rect 6184 15512 6236 15564
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 6828 15512 6880 15564
rect 7012 15555 7064 15564
rect 7012 15521 7021 15555
rect 7021 15521 7055 15555
rect 7055 15521 7064 15555
rect 7012 15512 7064 15521
rect 7196 15512 7248 15564
rect 6552 15487 6604 15496
rect 6552 15453 6561 15487
rect 6561 15453 6595 15487
rect 6595 15453 6604 15487
rect 6552 15444 6604 15453
rect 9036 15444 9088 15496
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 10876 15555 10928 15564
rect 10876 15521 10885 15555
rect 10885 15521 10919 15555
rect 10919 15521 10928 15555
rect 10876 15512 10928 15521
rect 11152 15512 11204 15564
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 5724 15308 5776 15360
rect 6644 15308 6696 15360
rect 6828 15376 6880 15428
rect 11336 15444 11388 15496
rect 13544 15512 13596 15564
rect 11612 15376 11664 15428
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 13452 15444 13504 15496
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 13820 15444 13872 15496
rect 14372 15512 14424 15564
rect 15016 15648 15068 15700
rect 18144 15648 18196 15700
rect 18420 15691 18472 15700
rect 18420 15657 18429 15691
rect 18429 15657 18463 15691
rect 18463 15657 18472 15691
rect 18420 15648 18472 15657
rect 18880 15648 18932 15700
rect 17868 15580 17920 15632
rect 18604 15580 18656 15632
rect 20996 15691 21048 15700
rect 20996 15657 21005 15691
rect 21005 15657 21039 15691
rect 21039 15657 21048 15691
rect 20996 15648 21048 15657
rect 21640 15648 21692 15700
rect 22468 15648 22520 15700
rect 23296 15691 23348 15700
rect 23296 15657 23305 15691
rect 23305 15657 23339 15691
rect 23339 15657 23348 15691
rect 23296 15648 23348 15657
rect 23480 15648 23532 15700
rect 15844 15512 15896 15564
rect 19984 15512 20036 15564
rect 23756 15580 23808 15632
rect 23940 15648 23992 15700
rect 26056 15648 26108 15700
rect 17960 15444 18012 15496
rect 18696 15444 18748 15496
rect 9956 15308 10008 15360
rect 11244 15308 11296 15360
rect 14096 15308 14148 15360
rect 14648 15308 14700 15360
rect 15660 15308 15712 15360
rect 15936 15351 15988 15360
rect 15936 15317 15945 15351
rect 15945 15317 15979 15351
rect 15979 15317 15988 15351
rect 15936 15308 15988 15317
rect 16304 15419 16356 15428
rect 16304 15385 16313 15419
rect 16313 15385 16347 15419
rect 16347 15385 16356 15419
rect 16304 15376 16356 15385
rect 17040 15376 17092 15428
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 21640 15512 21692 15564
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 23296 15512 23348 15564
rect 24308 15512 24360 15564
rect 22836 15487 22888 15496
rect 22836 15453 22845 15487
rect 22845 15453 22879 15487
rect 22879 15453 22888 15487
rect 22836 15444 22888 15453
rect 20168 15376 20220 15428
rect 19708 15308 19760 15360
rect 20996 15308 21048 15360
rect 21180 15308 21232 15360
rect 21916 15376 21968 15428
rect 22100 15308 22152 15360
rect 23204 15308 23256 15360
rect 23940 15487 23992 15496
rect 23940 15453 23949 15487
rect 23949 15453 23983 15487
rect 23983 15453 23992 15487
rect 23940 15444 23992 15453
rect 24952 15444 25004 15496
rect 25964 15444 26016 15496
rect 26240 15487 26292 15496
rect 26240 15453 26249 15487
rect 26249 15453 26283 15487
rect 26283 15453 26292 15487
rect 26240 15444 26292 15453
rect 26332 15444 26384 15496
rect 28172 15512 28224 15564
rect 27528 15487 27580 15496
rect 27528 15453 27537 15487
rect 27537 15453 27571 15487
rect 27571 15453 27580 15487
rect 27528 15444 27580 15453
rect 23848 15376 23900 15428
rect 28264 15444 28316 15496
rect 25044 15351 25096 15360
rect 25044 15317 25053 15351
rect 25053 15317 25087 15351
rect 25087 15317 25096 15351
rect 25044 15308 25096 15317
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 5324 15206 5376 15258
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 12752 15206 12804 15258
rect 12816 15206 12868 15258
rect 12880 15206 12932 15258
rect 12944 15206 12996 15258
rect 13008 15206 13060 15258
rect 20180 15206 20232 15258
rect 20244 15206 20296 15258
rect 20308 15206 20360 15258
rect 20372 15206 20424 15258
rect 20436 15206 20488 15258
rect 27608 15206 27660 15258
rect 27672 15206 27724 15258
rect 27736 15206 27788 15258
rect 27800 15206 27852 15258
rect 27864 15206 27916 15258
rect 6736 15104 6788 15156
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 6552 15036 6604 15088
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 4528 14900 4580 14952
rect 6736 14900 6788 14952
rect 7012 15036 7064 15088
rect 7104 15036 7156 15088
rect 8208 15036 8260 15088
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 10232 15104 10284 15156
rect 11060 15104 11112 15156
rect 9680 15036 9732 15088
rect 13820 15104 13872 15156
rect 12072 15079 12124 15088
rect 12072 15045 12081 15079
rect 12081 15045 12115 15079
rect 12115 15045 12124 15079
rect 12072 15036 12124 15045
rect 13636 15036 13688 15088
rect 16304 15104 16356 15156
rect 18052 15104 18104 15156
rect 18420 15104 18472 15156
rect 19708 15147 19760 15156
rect 19708 15113 19717 15147
rect 19717 15113 19751 15147
rect 19751 15113 19760 15147
rect 19708 15104 19760 15113
rect 20996 15104 21048 15156
rect 21088 15104 21140 15156
rect 11152 14968 11204 15020
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 7196 14900 7248 14952
rect 9772 14900 9824 14952
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 10876 14900 10928 14952
rect 2964 14764 3016 14816
rect 3884 14764 3936 14816
rect 4068 14764 4120 14816
rect 11796 14832 11848 14884
rect 11980 14832 12032 14884
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 14004 14968 14056 15020
rect 13360 14943 13412 14952
rect 13360 14909 13369 14943
rect 13369 14909 13403 14943
rect 13403 14909 13412 14943
rect 13360 14900 13412 14909
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 14740 15011 14792 15020
rect 14740 14977 14749 15011
rect 14749 14977 14783 15011
rect 14783 14977 14792 15011
rect 14740 14968 14792 14977
rect 15936 14968 15988 15020
rect 19340 15036 19392 15088
rect 21824 15104 21876 15156
rect 22652 15104 22704 15156
rect 25596 15104 25648 15156
rect 18788 15011 18840 15020
rect 18788 14977 18797 15011
rect 18797 14977 18831 15011
rect 18831 14977 18840 15011
rect 18788 14968 18840 14977
rect 19248 14968 19300 15020
rect 14280 14832 14332 14884
rect 18512 14900 18564 14952
rect 20812 14900 20864 14952
rect 13636 14764 13688 14816
rect 13820 14764 13872 14816
rect 15384 14764 15436 14816
rect 15660 14764 15712 14816
rect 17224 14764 17276 14816
rect 18696 14764 18748 14816
rect 19064 14832 19116 14884
rect 21180 14832 21232 14884
rect 21088 14764 21140 14816
rect 21732 14968 21784 15020
rect 21916 14968 21968 15020
rect 22008 15011 22060 15020
rect 22008 14977 22015 15011
rect 22015 14977 22049 15011
rect 22049 14977 22060 15011
rect 22008 14968 22060 14977
rect 22468 15079 22520 15088
rect 22468 15045 22477 15079
rect 22477 15045 22511 15079
rect 22511 15045 22520 15079
rect 22468 15036 22520 15045
rect 26240 15104 26292 15156
rect 21364 14900 21416 14952
rect 23756 14968 23808 15020
rect 24308 14968 24360 15020
rect 22284 14764 22336 14816
rect 25872 15011 25924 15020
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 26056 15011 26108 15020
rect 26056 14977 26065 15011
rect 26065 14977 26099 15011
rect 26099 14977 26108 15011
rect 26056 14968 26108 14977
rect 26148 15011 26200 15020
rect 26148 14977 26157 15011
rect 26157 14977 26191 15011
rect 26191 14977 26200 15011
rect 26148 14968 26200 14977
rect 26700 14968 26752 15020
rect 25964 14832 26016 14884
rect 27528 14900 27580 14952
rect 27712 14807 27764 14816
rect 27712 14773 27721 14807
rect 27721 14773 27755 14807
rect 27755 14773 27764 14807
rect 27712 14764 27764 14773
rect 28264 14807 28316 14816
rect 28264 14773 28273 14807
rect 28273 14773 28307 14807
rect 28307 14773 28316 14807
rect 28264 14764 28316 14773
rect 4664 14662 4716 14714
rect 4728 14662 4780 14714
rect 4792 14662 4844 14714
rect 4856 14662 4908 14714
rect 4920 14662 4972 14714
rect 12092 14662 12144 14714
rect 12156 14662 12208 14714
rect 12220 14662 12272 14714
rect 12284 14662 12336 14714
rect 12348 14662 12400 14714
rect 19520 14662 19572 14714
rect 19584 14662 19636 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 26948 14662 27000 14714
rect 27012 14662 27064 14714
rect 27076 14662 27128 14714
rect 27140 14662 27192 14714
rect 27204 14662 27256 14714
rect 3516 14560 3568 14612
rect 5724 14560 5776 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 6828 14560 6880 14612
rect 9680 14560 9732 14612
rect 9772 14603 9824 14612
rect 9772 14569 9781 14603
rect 9781 14569 9815 14603
rect 9815 14569 9824 14603
rect 9772 14560 9824 14569
rect 11152 14560 11204 14612
rect 11888 14560 11940 14612
rect 4988 14492 5040 14544
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 3976 14356 4028 14408
rect 4344 14356 4396 14408
rect 7380 14467 7432 14476
rect 7380 14433 7389 14467
rect 7389 14433 7423 14467
rect 7423 14433 7432 14467
rect 7380 14424 7432 14433
rect 2136 14331 2188 14340
rect 2136 14297 2145 14331
rect 2145 14297 2179 14331
rect 2179 14297 2188 14331
rect 2136 14288 2188 14297
rect 3148 14288 3200 14340
rect 4528 14288 4580 14340
rect 1676 14220 1728 14272
rect 3884 14220 3936 14272
rect 4068 14220 4120 14272
rect 4160 14220 4212 14272
rect 6828 14356 6880 14408
rect 7104 14356 7156 14408
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 7748 14331 7800 14340
rect 7748 14297 7757 14331
rect 7757 14297 7791 14331
rect 7791 14297 7800 14331
rect 7748 14288 7800 14297
rect 8024 14331 8076 14340
rect 8024 14297 8033 14331
rect 8033 14297 8067 14331
rect 8067 14297 8076 14331
rect 8024 14288 8076 14297
rect 8116 14331 8168 14340
rect 8116 14297 8125 14331
rect 8125 14297 8159 14331
rect 8159 14297 8168 14331
rect 8116 14288 8168 14297
rect 8208 14288 8260 14340
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 11796 14492 11848 14544
rect 16948 14560 17000 14612
rect 17224 14560 17276 14612
rect 20536 14560 20588 14612
rect 21364 14560 21416 14612
rect 9956 14399 10008 14408
rect 9956 14365 9965 14399
rect 9965 14365 9999 14399
rect 9999 14365 10008 14399
rect 9956 14356 10008 14365
rect 11520 14424 11572 14476
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 12072 14424 12124 14476
rect 18788 14492 18840 14544
rect 13176 14356 13228 14408
rect 13544 14356 13596 14408
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 16120 14356 16172 14408
rect 6736 14220 6788 14272
rect 7932 14220 7984 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 11244 14288 11296 14340
rect 16580 14288 16632 14340
rect 17776 14356 17828 14408
rect 17868 14356 17920 14408
rect 17684 14331 17736 14340
rect 17684 14297 17693 14331
rect 17693 14297 17727 14331
rect 17727 14297 17736 14331
rect 17684 14288 17736 14297
rect 18972 14356 19024 14408
rect 19248 14424 19300 14476
rect 19524 14356 19576 14408
rect 20076 14356 20128 14408
rect 18880 14288 18932 14340
rect 19156 14288 19208 14340
rect 22100 14424 22152 14476
rect 22468 14492 22520 14544
rect 23112 14560 23164 14612
rect 23664 14603 23716 14612
rect 23664 14569 23673 14603
rect 23673 14569 23707 14603
rect 23707 14569 23716 14603
rect 23664 14560 23716 14569
rect 23940 14560 23992 14612
rect 24308 14560 24360 14612
rect 24952 14560 25004 14612
rect 25044 14560 25096 14612
rect 21916 14399 21968 14408
rect 21916 14365 21925 14399
rect 21925 14365 21959 14399
rect 21959 14365 21968 14399
rect 21916 14356 21968 14365
rect 25872 14492 25924 14544
rect 27712 14603 27764 14612
rect 27712 14569 27721 14603
rect 27721 14569 27755 14603
rect 27755 14569 27764 14603
rect 27712 14560 27764 14569
rect 28264 14560 28316 14612
rect 24032 14356 24084 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 22008 14288 22060 14340
rect 22284 14288 22336 14340
rect 23848 14288 23900 14340
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 25228 14399 25280 14408
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 25320 14356 25372 14408
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 26148 14356 26200 14408
rect 25504 14331 25556 14340
rect 25504 14297 25513 14331
rect 25513 14297 25547 14331
rect 25547 14297 25556 14331
rect 25504 14288 25556 14297
rect 13268 14220 13320 14272
rect 14648 14220 14700 14272
rect 16212 14263 16264 14272
rect 16212 14229 16221 14263
rect 16221 14229 16255 14263
rect 16255 14229 16264 14263
rect 16212 14220 16264 14229
rect 16856 14220 16908 14272
rect 18144 14220 18196 14272
rect 19248 14220 19300 14272
rect 22192 14220 22244 14272
rect 22744 14263 22796 14272
rect 22744 14229 22753 14263
rect 22753 14229 22787 14263
rect 22787 14229 22796 14263
rect 22744 14220 22796 14229
rect 23204 14220 23256 14272
rect 24860 14220 24912 14272
rect 24952 14220 25004 14272
rect 26148 14220 26200 14272
rect 26332 14220 26384 14272
rect 5324 14118 5376 14170
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 12752 14118 12804 14170
rect 12816 14118 12868 14170
rect 12880 14118 12932 14170
rect 12944 14118 12996 14170
rect 13008 14118 13060 14170
rect 20180 14118 20232 14170
rect 20244 14118 20296 14170
rect 20308 14118 20360 14170
rect 20372 14118 20424 14170
rect 20436 14118 20488 14170
rect 27608 14118 27660 14170
rect 27672 14118 27724 14170
rect 27736 14118 27788 14170
rect 27800 14118 27852 14170
rect 27864 14118 27916 14170
rect 2136 14016 2188 14068
rect 940 13880 992 13932
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2964 14016 3016 14068
rect 3148 14016 3200 14068
rect 3516 14016 3568 14068
rect 4344 14016 4396 14068
rect 7288 14016 7340 14068
rect 4068 13880 4120 13932
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 7472 13948 7524 14000
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 3608 13744 3660 13796
rect 6644 13855 6696 13864
rect 6644 13821 6653 13855
rect 6653 13821 6687 13855
rect 6687 13821 6696 13855
rect 6644 13812 6696 13821
rect 8116 14016 8168 14068
rect 7932 13948 7984 14000
rect 8484 14016 8536 14068
rect 9128 14016 9180 14068
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 9680 14016 9732 14068
rect 8024 13923 8076 13932
rect 8024 13889 8033 13923
rect 8033 13889 8067 13923
rect 8067 13889 8076 13923
rect 8024 13880 8076 13889
rect 7932 13855 7984 13864
rect 7932 13821 7941 13855
rect 7941 13821 7975 13855
rect 7975 13821 7984 13855
rect 7932 13812 7984 13821
rect 3976 13676 4028 13728
rect 4068 13676 4120 13728
rect 5540 13744 5592 13796
rect 8116 13812 8168 13864
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 10140 13948 10192 14000
rect 10876 13948 10928 14000
rect 11152 14016 11204 14068
rect 11796 14016 11848 14068
rect 11612 13948 11664 14000
rect 11704 13948 11756 14000
rect 9680 13880 9732 13932
rect 9220 13812 9272 13864
rect 9588 13812 9640 13864
rect 13084 13880 13136 13932
rect 13912 13880 13964 13932
rect 14556 14016 14608 14068
rect 16120 13880 16172 13932
rect 17684 14016 17736 14068
rect 17776 14016 17828 14068
rect 19064 14016 19116 14068
rect 22744 14016 22796 14068
rect 23664 14016 23716 14068
rect 24860 14016 24912 14068
rect 25504 14016 25556 14068
rect 25872 14016 25924 14068
rect 18880 13880 18932 13932
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19248 13923 19300 13932
rect 19248 13889 19257 13923
rect 19257 13889 19291 13923
rect 19291 13889 19300 13923
rect 19248 13880 19300 13889
rect 19616 13880 19668 13932
rect 21456 13948 21508 14000
rect 20996 13880 21048 13932
rect 21088 13880 21140 13932
rect 22100 13880 22152 13932
rect 11980 13855 12032 13864
rect 11980 13821 11989 13855
rect 11989 13821 12023 13855
rect 12023 13821 12032 13855
rect 11980 13812 12032 13821
rect 13544 13812 13596 13864
rect 9956 13744 10008 13796
rect 9496 13676 9548 13728
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14648 13812 14700 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 16856 13812 16908 13864
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 22008 13744 22060 13796
rect 22836 13744 22888 13796
rect 15292 13676 15344 13728
rect 22744 13676 22796 13728
rect 23204 13880 23256 13932
rect 25044 13948 25096 14000
rect 23480 13880 23532 13932
rect 24768 13880 24820 13932
rect 23848 13744 23900 13796
rect 24032 13744 24084 13796
rect 25320 13880 25372 13932
rect 26240 13855 26292 13864
rect 26240 13821 26249 13855
rect 26249 13821 26283 13855
rect 26283 13821 26292 13855
rect 26240 13812 26292 13821
rect 25136 13719 25188 13728
rect 25136 13685 25145 13719
rect 25145 13685 25179 13719
rect 25179 13685 25188 13719
rect 25136 13676 25188 13685
rect 26148 13719 26200 13728
rect 26148 13685 26157 13719
rect 26157 13685 26191 13719
rect 26191 13685 26200 13719
rect 26148 13676 26200 13685
rect 26516 13719 26568 13728
rect 26516 13685 26525 13719
rect 26525 13685 26559 13719
rect 26559 13685 26568 13719
rect 26516 13676 26568 13685
rect 4664 13574 4716 13626
rect 4728 13574 4780 13626
rect 4792 13574 4844 13626
rect 4856 13574 4908 13626
rect 4920 13574 4972 13626
rect 12092 13574 12144 13626
rect 12156 13574 12208 13626
rect 12220 13574 12272 13626
rect 12284 13574 12336 13626
rect 12348 13574 12400 13626
rect 19520 13574 19572 13626
rect 19584 13574 19636 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 26948 13574 27000 13626
rect 27012 13574 27064 13626
rect 27076 13574 27128 13626
rect 27140 13574 27192 13626
rect 27204 13574 27256 13626
rect 6644 13515 6696 13524
rect 4252 13268 4304 13320
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 8300 13472 8352 13524
rect 8852 13472 8904 13524
rect 16580 13472 16632 13524
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 23756 13472 23808 13524
rect 26240 13472 26292 13524
rect 28356 13472 28408 13524
rect 9404 13404 9456 13456
rect 9588 13404 9640 13456
rect 19432 13404 19484 13456
rect 7196 13336 7248 13388
rect 11888 13336 11940 13388
rect 5540 13268 5592 13320
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 8024 13311 8076 13320
rect 8024 13277 8033 13311
rect 8033 13277 8067 13311
rect 8067 13277 8076 13311
rect 8024 13268 8076 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10232 13268 10284 13320
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 16212 13336 16264 13388
rect 14556 13268 14608 13320
rect 15292 13268 15344 13320
rect 11428 13243 11480 13252
rect 11428 13209 11437 13243
rect 11437 13209 11471 13243
rect 11471 13209 11480 13243
rect 11428 13200 11480 13209
rect 12164 13200 12216 13252
rect 16672 13268 16724 13320
rect 17776 13336 17828 13388
rect 18512 13336 18564 13388
rect 20812 13336 20864 13388
rect 21088 13336 21140 13388
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 18144 13311 18196 13320
rect 18144 13277 18153 13311
rect 18153 13277 18187 13311
rect 18187 13277 18196 13311
rect 18144 13268 18196 13277
rect 18880 13268 18932 13320
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 8668 13132 8720 13184
rect 11244 13132 11296 13184
rect 13084 13132 13136 13184
rect 16948 13200 17000 13252
rect 18328 13200 18380 13252
rect 20996 13268 21048 13320
rect 22192 13379 22244 13388
rect 22192 13345 22201 13379
rect 22201 13345 22235 13379
rect 22235 13345 22244 13379
rect 22192 13336 22244 13345
rect 22284 13379 22336 13388
rect 22284 13345 22293 13379
rect 22293 13345 22327 13379
rect 22327 13345 22336 13379
rect 22284 13336 22336 13345
rect 22744 13336 22796 13388
rect 22836 13336 22888 13388
rect 23480 13336 23532 13388
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 21364 13200 21416 13252
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 24768 13336 24820 13388
rect 26516 13447 26568 13456
rect 26516 13413 26525 13447
rect 26525 13413 26559 13447
rect 26559 13413 26568 13447
rect 26516 13404 26568 13413
rect 27344 13336 27396 13388
rect 25136 13268 25188 13320
rect 16856 13175 16908 13184
rect 16856 13141 16865 13175
rect 16865 13141 16899 13175
rect 16899 13141 16908 13175
rect 16856 13132 16908 13141
rect 20628 13132 20680 13184
rect 24676 13132 24728 13184
rect 25504 13132 25556 13184
rect 26332 13311 26384 13320
rect 26332 13277 26341 13311
rect 26341 13277 26375 13311
rect 26375 13277 26384 13311
rect 26332 13268 26384 13277
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26148 13200 26200 13252
rect 5324 13030 5376 13082
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 12752 13030 12804 13082
rect 12816 13030 12868 13082
rect 12880 13030 12932 13082
rect 12944 13030 12996 13082
rect 13008 13030 13060 13082
rect 20180 13030 20232 13082
rect 20244 13030 20296 13082
rect 20308 13030 20360 13082
rect 20372 13030 20424 13082
rect 20436 13030 20488 13082
rect 27608 13030 27660 13082
rect 27672 13030 27724 13082
rect 27736 13030 27788 13082
rect 27800 13030 27852 13082
rect 27864 13030 27916 13082
rect 7104 12928 7156 12980
rect 3976 12860 4028 12912
rect 2780 12835 2832 12844
rect 2780 12801 2789 12835
rect 2789 12801 2823 12835
rect 2823 12801 2832 12835
rect 2780 12792 2832 12801
rect 4160 12792 4212 12844
rect 4528 12792 4580 12844
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 6460 12860 6512 12912
rect 8760 12928 8812 12980
rect 8852 12903 8904 12912
rect 8852 12869 8861 12903
rect 8861 12869 8895 12903
rect 8895 12869 8904 12903
rect 8852 12860 8904 12869
rect 9772 12928 9824 12980
rect 9588 12860 9640 12912
rect 11336 12928 11388 12980
rect 11428 12928 11480 12980
rect 8300 12792 8352 12844
rect 9312 12792 9364 12844
rect 9404 12792 9456 12844
rect 9680 12792 9732 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 10600 12792 10652 12844
rect 13084 12928 13136 12980
rect 13912 12928 13964 12980
rect 11888 12860 11940 12912
rect 12164 12903 12216 12912
rect 12164 12869 12173 12903
rect 12173 12869 12207 12903
rect 12207 12869 12216 12903
rect 12164 12860 12216 12869
rect 14556 12903 14608 12912
rect 14556 12869 14565 12903
rect 14565 12869 14599 12903
rect 14599 12869 14608 12903
rect 14556 12860 14608 12869
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 16672 12971 16724 12980
rect 16672 12937 16681 12971
rect 16681 12937 16715 12971
rect 16715 12937 16724 12971
rect 16672 12928 16724 12937
rect 16856 12928 16908 12980
rect 16948 12928 17000 12980
rect 17040 12928 17092 12980
rect 17684 12928 17736 12980
rect 19984 12928 20036 12980
rect 22284 12928 22336 12980
rect 22468 12928 22520 12980
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 26424 12928 26476 12980
rect 1860 12724 1912 12776
rect 7012 12724 7064 12776
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 8944 12724 8996 12776
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 6092 12699 6144 12708
rect 6092 12665 6101 12699
rect 6101 12665 6135 12699
rect 6135 12665 6144 12699
rect 6092 12656 6144 12665
rect 10508 12724 10560 12776
rect 11244 12656 11296 12708
rect 17132 12724 17184 12776
rect 17224 12724 17276 12776
rect 18236 12860 18288 12912
rect 17408 12699 17460 12708
rect 17408 12665 17417 12699
rect 17417 12665 17451 12699
rect 17451 12665 17460 12699
rect 17408 12656 17460 12665
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 7472 12588 7524 12640
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 9404 12588 9456 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 11612 12588 11664 12640
rect 11980 12588 12032 12640
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 16212 12588 16264 12640
rect 18696 12792 18748 12844
rect 20536 12860 20588 12912
rect 23204 12835 23256 12844
rect 23204 12801 23213 12835
rect 23213 12801 23247 12835
rect 23247 12801 23256 12835
rect 23204 12792 23256 12801
rect 23020 12724 23072 12776
rect 23572 12792 23624 12844
rect 24032 12792 24084 12844
rect 24676 12835 24728 12844
rect 24676 12801 24685 12835
rect 24685 12801 24719 12835
rect 24719 12801 24728 12835
rect 24676 12792 24728 12801
rect 25504 12835 25556 12844
rect 25504 12801 25513 12835
rect 25513 12801 25547 12835
rect 25547 12801 25556 12835
rect 25504 12792 25556 12801
rect 21548 12631 21600 12640
rect 21548 12597 21557 12631
rect 21557 12597 21591 12631
rect 21591 12597 21600 12631
rect 21548 12588 21600 12597
rect 25136 12724 25188 12776
rect 25964 12860 26016 12912
rect 26148 12792 26200 12844
rect 4664 12486 4716 12538
rect 4728 12486 4780 12538
rect 4792 12486 4844 12538
rect 4856 12486 4908 12538
rect 4920 12486 4972 12538
rect 12092 12486 12144 12538
rect 12156 12486 12208 12538
rect 12220 12486 12272 12538
rect 12284 12486 12336 12538
rect 12348 12486 12400 12538
rect 19520 12486 19572 12538
rect 19584 12486 19636 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 26948 12486 27000 12538
rect 27012 12486 27064 12538
rect 27076 12486 27128 12538
rect 27140 12486 27192 12538
rect 27204 12486 27256 12538
rect 2780 12384 2832 12436
rect 1860 12291 1912 12300
rect 1860 12257 1869 12291
rect 1869 12257 1903 12291
rect 1903 12257 1912 12291
rect 1860 12248 1912 12257
rect 2596 12248 2648 12300
rect 3976 12248 4028 12300
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 5080 12248 5132 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 3240 12180 3292 12232
rect 3792 12180 3844 12232
rect 6460 12180 6512 12232
rect 7472 12316 7524 12368
rect 8300 12427 8352 12436
rect 8300 12393 8309 12427
rect 8309 12393 8343 12427
rect 8343 12393 8352 12427
rect 8300 12384 8352 12393
rect 9220 12384 9272 12436
rect 9312 12384 9364 12436
rect 9680 12384 9732 12436
rect 10048 12384 10100 12436
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 8484 12291 8536 12300
rect 8484 12257 8507 12291
rect 8507 12257 8536 12291
rect 8484 12248 8536 12257
rect 6920 12044 6972 12096
rect 7656 12112 7708 12164
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 14188 12384 14240 12436
rect 21364 12427 21416 12436
rect 21364 12393 21373 12427
rect 21373 12393 21407 12427
rect 21407 12393 21416 12427
rect 21364 12384 21416 12393
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 15568 12248 15620 12300
rect 17132 12248 17184 12300
rect 19340 12248 19392 12300
rect 19984 12248 20036 12300
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 16212 12180 16264 12232
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 19248 12180 19300 12232
rect 21548 12180 21600 12232
rect 21732 12223 21784 12232
rect 21732 12189 21741 12223
rect 21741 12189 21775 12223
rect 21775 12189 21784 12223
rect 21732 12180 21784 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 19984 12112 20036 12164
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 15200 12087 15252 12096
rect 15200 12053 15209 12087
rect 15209 12053 15243 12087
rect 15243 12053 15252 12087
rect 15200 12044 15252 12053
rect 15384 12087 15436 12096
rect 15384 12053 15393 12087
rect 15393 12053 15427 12087
rect 15427 12053 15436 12087
rect 15384 12044 15436 12053
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 17776 12044 17828 12096
rect 18696 12044 18748 12096
rect 21916 12087 21968 12096
rect 21916 12053 21925 12087
rect 21925 12053 21959 12087
rect 21959 12053 21968 12087
rect 21916 12044 21968 12053
rect 23020 12044 23072 12096
rect 5324 11942 5376 11994
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 12752 11942 12804 11994
rect 12816 11942 12868 11994
rect 12880 11942 12932 11994
rect 12944 11942 12996 11994
rect 13008 11942 13060 11994
rect 20180 11942 20232 11994
rect 20244 11942 20296 11994
rect 20308 11942 20360 11994
rect 20372 11942 20424 11994
rect 20436 11942 20488 11994
rect 27608 11942 27660 11994
rect 27672 11942 27724 11994
rect 27736 11942 27788 11994
rect 27800 11942 27852 11994
rect 27864 11942 27916 11994
rect 3240 11883 3292 11892
rect 3240 11849 3249 11883
rect 3249 11849 3283 11883
rect 3283 11849 3292 11883
rect 3240 11840 3292 11849
rect 3608 11840 3660 11892
rect 5172 11840 5224 11892
rect 6460 11840 6512 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 9680 11840 9732 11892
rect 10784 11840 10836 11892
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 10140 11772 10192 11824
rect 12440 11772 12492 11824
rect 3332 11704 3384 11713
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11244 11704 11296 11756
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 13452 11704 13504 11756
rect 14188 11772 14240 11824
rect 15200 11840 15252 11892
rect 16948 11815 17000 11824
rect 16948 11781 16957 11815
rect 16957 11781 16991 11815
rect 16991 11781 17000 11815
rect 16948 11772 17000 11781
rect 19984 11840 20036 11892
rect 21732 11840 21784 11892
rect 21916 11840 21968 11892
rect 6184 11611 6236 11620
rect 6184 11577 6193 11611
rect 6193 11577 6227 11611
rect 6227 11577 6236 11611
rect 6184 11568 6236 11577
rect 10048 11568 10100 11620
rect 17316 11704 17368 11756
rect 17408 11704 17460 11756
rect 17684 11704 17736 11756
rect 17224 11636 17276 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 20076 11704 20128 11756
rect 20628 11704 20680 11756
rect 23020 11772 23072 11824
rect 20996 11636 21048 11688
rect 21088 11679 21140 11688
rect 21088 11645 21097 11679
rect 21097 11645 21131 11679
rect 21131 11645 21140 11679
rect 21088 11636 21140 11645
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 23940 11704 23992 11756
rect 9404 11500 9456 11552
rect 9680 11500 9732 11552
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 14924 11500 14976 11552
rect 17776 11500 17828 11552
rect 18236 11500 18288 11552
rect 18328 11500 18380 11552
rect 18420 11500 18472 11552
rect 19432 11500 19484 11552
rect 19984 11500 20036 11552
rect 23848 11636 23900 11688
rect 24308 11543 24360 11552
rect 24308 11509 24317 11543
rect 24317 11509 24351 11543
rect 24351 11509 24360 11543
rect 24308 11500 24360 11509
rect 4664 11398 4716 11450
rect 4728 11398 4780 11450
rect 4792 11398 4844 11450
rect 4856 11398 4908 11450
rect 4920 11398 4972 11450
rect 12092 11398 12144 11450
rect 12156 11398 12208 11450
rect 12220 11398 12272 11450
rect 12284 11398 12336 11450
rect 12348 11398 12400 11450
rect 19520 11398 19572 11450
rect 19584 11398 19636 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 26948 11398 27000 11450
rect 27012 11398 27064 11450
rect 27076 11398 27128 11450
rect 27140 11398 27192 11450
rect 27204 11398 27256 11450
rect 1860 11296 1912 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 9588 11296 9640 11348
rect 10140 11296 10192 11348
rect 11152 11296 11204 11348
rect 12440 11296 12492 11348
rect 9128 11228 9180 11280
rect 3148 11092 3200 11144
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 5724 11024 5776 11076
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 10048 11092 10100 11144
rect 14924 11296 14976 11348
rect 15476 11339 15528 11348
rect 15476 11305 15485 11339
rect 15485 11305 15519 11339
rect 15519 11305 15528 11339
rect 15476 11296 15528 11305
rect 16948 11296 17000 11348
rect 13544 11228 13596 11280
rect 15844 11271 15896 11280
rect 15844 11237 15853 11271
rect 15853 11237 15887 11271
rect 15887 11237 15896 11271
rect 15844 11228 15896 11237
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 13452 11160 13504 11212
rect 15016 11160 15068 11212
rect 13636 11092 13688 11144
rect 17776 11160 17828 11212
rect 17132 11135 17184 11144
rect 6644 10956 6696 11008
rect 8576 10956 8628 11008
rect 11796 11024 11848 11076
rect 13452 11024 13504 11076
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 16488 11024 16540 11076
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 17408 11024 17460 11076
rect 18328 11024 18380 11076
rect 21088 11296 21140 11348
rect 21180 11296 21232 11348
rect 24308 11296 24360 11348
rect 25044 11296 25096 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 21824 11228 21876 11280
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 23940 11228 23992 11280
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 23480 11092 23532 11144
rect 23848 11135 23900 11144
rect 23848 11101 23857 11135
rect 23857 11101 23891 11135
rect 23891 11101 23900 11135
rect 23848 11092 23900 11101
rect 13820 10999 13872 11008
rect 13820 10965 13829 10999
rect 13829 10965 13863 10999
rect 13863 10965 13872 10999
rect 13820 10956 13872 10965
rect 14832 10956 14884 11008
rect 15568 10956 15620 11008
rect 19892 11024 19944 11076
rect 21824 11067 21876 11076
rect 21824 11033 21833 11067
rect 21833 11033 21867 11067
rect 21867 11033 21876 11067
rect 21824 11024 21876 11033
rect 24492 11135 24544 11144
rect 24492 11101 24501 11135
rect 24501 11101 24535 11135
rect 24535 11101 24544 11135
rect 24492 11092 24544 11101
rect 24676 11135 24728 11144
rect 24676 11101 24683 11135
rect 24683 11101 24728 11135
rect 24676 11092 24728 11101
rect 24860 11160 24912 11212
rect 25044 11160 25096 11212
rect 25504 11203 25556 11212
rect 25504 11169 25513 11203
rect 25513 11169 25547 11203
rect 25547 11169 25556 11203
rect 25504 11160 25556 11169
rect 20076 10956 20128 11008
rect 20628 10956 20680 11008
rect 23204 10956 23256 11008
rect 23848 10956 23900 11008
rect 25412 10956 25464 11008
rect 5324 10854 5376 10906
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 12752 10854 12804 10906
rect 12816 10854 12868 10906
rect 12880 10854 12932 10906
rect 12944 10854 12996 10906
rect 13008 10854 13060 10906
rect 20180 10854 20232 10906
rect 20244 10854 20296 10906
rect 20308 10854 20360 10906
rect 20372 10854 20424 10906
rect 20436 10854 20488 10906
rect 27608 10854 27660 10906
rect 27672 10854 27724 10906
rect 27736 10854 27788 10906
rect 27800 10854 27852 10906
rect 27864 10854 27916 10906
rect 2044 10752 2096 10804
rect 3148 10752 3200 10804
rect 3792 10752 3844 10804
rect 3976 10752 4028 10804
rect 4896 10684 4948 10736
rect 7380 10752 7432 10804
rect 7656 10752 7708 10804
rect 8392 10752 8444 10804
rect 13360 10752 13412 10804
rect 3332 10659 3384 10668
rect 3332 10625 3341 10659
rect 3341 10625 3375 10659
rect 3375 10625 3384 10659
rect 3332 10616 3384 10625
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4160 10616 4212 10668
rect 4528 10616 4580 10668
rect 4804 10616 4856 10668
rect 5724 10684 5776 10736
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 6828 10616 6880 10668
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 8300 10659 8352 10668
rect 8300 10625 8309 10659
rect 8309 10625 8343 10659
rect 8343 10625 8352 10659
rect 8300 10616 8352 10625
rect 8392 10616 8444 10668
rect 9220 10684 9272 10736
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 5080 10480 5132 10532
rect 9036 10591 9088 10600
rect 9036 10557 9045 10591
rect 9045 10557 9079 10591
rect 9079 10557 9088 10591
rect 9036 10548 9088 10557
rect 10048 10548 10100 10600
rect 12624 10616 12676 10668
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 13820 10616 13872 10668
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 15108 10752 15160 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 15384 10752 15436 10804
rect 17132 10752 17184 10804
rect 18512 10752 18564 10804
rect 8852 10412 8904 10464
rect 13912 10480 13964 10532
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 13176 10455 13228 10464
rect 13176 10421 13185 10455
rect 13185 10421 13219 10455
rect 13219 10421 13228 10455
rect 13176 10412 13228 10421
rect 15476 10616 15528 10668
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 16948 10616 17000 10668
rect 17316 10659 17368 10668
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 16488 10548 16540 10600
rect 17960 10616 18012 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 19984 10752 20036 10804
rect 19892 10684 19944 10736
rect 21824 10684 21876 10736
rect 22192 10752 22244 10804
rect 23940 10752 23992 10804
rect 24492 10752 24544 10804
rect 24860 10752 24912 10804
rect 25412 10752 25464 10804
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 23020 10616 23072 10668
rect 23848 10616 23900 10668
rect 24308 10616 24360 10668
rect 24584 10616 24636 10668
rect 15568 10480 15620 10532
rect 17132 10480 17184 10532
rect 19248 10480 19300 10532
rect 21088 10548 21140 10600
rect 22744 10548 22796 10600
rect 25320 10548 25372 10600
rect 15936 10412 15988 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 19892 10412 19944 10464
rect 22284 10455 22336 10464
rect 22284 10421 22293 10455
rect 22293 10421 22327 10455
rect 22327 10421 22336 10455
rect 22284 10412 22336 10421
rect 22560 10455 22612 10464
rect 22560 10421 22569 10455
rect 22569 10421 22603 10455
rect 22603 10421 22612 10455
rect 22560 10412 22612 10421
rect 4664 10310 4716 10362
rect 4728 10310 4780 10362
rect 4792 10310 4844 10362
rect 4856 10310 4908 10362
rect 4920 10310 4972 10362
rect 12092 10310 12144 10362
rect 12156 10310 12208 10362
rect 12220 10310 12272 10362
rect 12284 10310 12336 10362
rect 12348 10310 12400 10362
rect 19520 10310 19572 10362
rect 19584 10310 19636 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 26948 10310 27000 10362
rect 27012 10310 27064 10362
rect 27076 10310 27128 10362
rect 27140 10310 27192 10362
rect 27204 10310 27256 10362
rect 7932 10208 7984 10260
rect 9864 10208 9916 10260
rect 9956 10208 10008 10260
rect 13176 10208 13228 10260
rect 5172 10004 5224 10056
rect 6276 10004 6328 10056
rect 13544 10208 13596 10260
rect 9220 10004 9272 10056
rect 9312 10004 9364 10056
rect 9036 9979 9088 9988
rect 9036 9945 9045 9979
rect 9045 9945 9079 9979
rect 9079 9945 9088 9979
rect 9036 9936 9088 9945
rect 6736 9868 6788 9920
rect 8576 9868 8628 9920
rect 10600 9911 10652 9920
rect 10600 9877 10609 9911
rect 10609 9877 10643 9911
rect 10643 9877 10652 9911
rect 10600 9868 10652 9877
rect 12532 9868 12584 9920
rect 13084 10004 13136 10056
rect 13360 10004 13412 10056
rect 15384 10208 15436 10260
rect 17316 10208 17368 10260
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 16856 10072 16908 10124
rect 17316 10115 17368 10124
rect 17316 10081 17325 10115
rect 17325 10081 17359 10115
rect 17359 10081 17368 10115
rect 17316 10072 17368 10081
rect 19340 10072 19392 10124
rect 19524 10004 19576 10056
rect 20812 10140 20864 10192
rect 20904 10183 20956 10192
rect 20904 10149 20913 10183
rect 20913 10149 20947 10183
rect 20947 10149 20956 10183
rect 20904 10140 20956 10149
rect 20536 10072 20588 10124
rect 16488 9936 16540 9988
rect 16580 9868 16632 9920
rect 16764 9911 16816 9920
rect 16764 9877 16773 9911
rect 16773 9877 16807 9911
rect 16807 9877 16816 9911
rect 16764 9868 16816 9877
rect 17500 9936 17552 9988
rect 21180 10004 21232 10056
rect 22008 10072 22060 10124
rect 22284 10208 22336 10260
rect 23020 10208 23072 10260
rect 25504 10208 25556 10260
rect 25964 10251 26016 10260
rect 25964 10217 25973 10251
rect 25973 10217 26007 10251
rect 26007 10217 26016 10251
rect 25964 10208 26016 10217
rect 24768 10183 24820 10192
rect 24768 10149 24777 10183
rect 24777 10149 24811 10183
rect 24811 10149 24820 10183
rect 24768 10140 24820 10149
rect 25780 10072 25832 10124
rect 18236 9868 18288 9920
rect 19156 9868 19208 9920
rect 20904 9936 20956 9988
rect 20628 9868 20680 9920
rect 22376 10004 22428 10056
rect 22560 10047 22612 10056
rect 22560 10013 22569 10047
rect 22569 10013 22603 10047
rect 22603 10013 22612 10047
rect 22560 10004 22612 10013
rect 24860 10004 24912 10056
rect 24584 9936 24636 9988
rect 25412 9936 25464 9988
rect 22652 9911 22704 9920
rect 22652 9877 22661 9911
rect 22661 9877 22695 9911
rect 22695 9877 22704 9911
rect 22652 9868 22704 9877
rect 23020 9868 23072 9920
rect 25964 9868 26016 9920
rect 5324 9766 5376 9818
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 12752 9766 12804 9818
rect 12816 9766 12868 9818
rect 12880 9766 12932 9818
rect 12944 9766 12996 9818
rect 13008 9766 13060 9818
rect 20180 9766 20232 9818
rect 20244 9766 20296 9818
rect 20308 9766 20360 9818
rect 20372 9766 20424 9818
rect 20436 9766 20488 9818
rect 27608 9766 27660 9818
rect 27672 9766 27724 9818
rect 27736 9766 27788 9818
rect 27800 9766 27852 9818
rect 27864 9766 27916 9818
rect 3608 9596 3660 9648
rect 4068 9596 4120 9648
rect 9312 9664 9364 9716
rect 12624 9707 12676 9716
rect 12624 9673 12633 9707
rect 12633 9673 12667 9707
rect 12667 9673 12676 9707
rect 12624 9664 12676 9673
rect 6736 9596 6788 9648
rect 12348 9596 12400 9648
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5356 9528 5408 9580
rect 5540 9528 5592 9580
rect 3332 9324 3384 9376
rect 4160 9367 4212 9376
rect 4160 9333 4169 9367
rect 4169 9333 4203 9367
rect 4203 9333 4212 9367
rect 4160 9324 4212 9333
rect 6184 9503 6236 9512
rect 6184 9469 6193 9503
rect 6193 9469 6227 9503
rect 6227 9469 6236 9503
rect 6184 9460 6236 9469
rect 8576 9528 8628 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9680 9571 9732 9580
rect 9680 9537 9682 9571
rect 9682 9537 9716 9571
rect 9716 9537 9732 9571
rect 9680 9528 9732 9537
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12440 9528 12492 9580
rect 13268 9664 13320 9716
rect 16764 9664 16816 9716
rect 16580 9596 16632 9648
rect 5172 9392 5224 9444
rect 8576 9435 8628 9444
rect 8576 9401 8585 9435
rect 8585 9401 8619 9435
rect 8619 9401 8628 9435
rect 8576 9392 8628 9401
rect 9220 9460 9272 9512
rect 9496 9392 9548 9444
rect 11244 9460 11296 9512
rect 12716 9392 12768 9444
rect 12624 9324 12676 9376
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 14188 9528 14240 9580
rect 15016 9528 15068 9580
rect 15844 9528 15896 9580
rect 16856 9528 16908 9580
rect 17132 9571 17184 9580
rect 17132 9537 17141 9571
rect 17141 9537 17175 9571
rect 17175 9537 17184 9571
rect 17132 9528 17184 9537
rect 16028 9460 16080 9512
rect 16948 9460 17000 9512
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 19156 9664 19208 9716
rect 22560 9664 22612 9716
rect 22652 9664 22704 9716
rect 17316 9528 17368 9537
rect 18144 9528 18196 9580
rect 22836 9639 22888 9648
rect 22836 9605 22845 9639
rect 22845 9605 22879 9639
rect 22879 9605 22888 9639
rect 22836 9596 22888 9605
rect 23480 9596 23532 9648
rect 24768 9596 24820 9648
rect 24952 9596 25004 9648
rect 17408 9460 17460 9512
rect 16396 9392 16448 9444
rect 13176 9367 13228 9376
rect 13176 9333 13185 9367
rect 13185 9333 13219 9367
rect 13219 9333 13228 9367
rect 13176 9324 13228 9333
rect 16764 9324 16816 9376
rect 18236 9324 18288 9376
rect 19524 9324 19576 9376
rect 20536 9324 20588 9376
rect 22744 9528 22796 9580
rect 22928 9460 22980 9512
rect 25044 9571 25096 9580
rect 25044 9537 25053 9571
rect 25053 9537 25087 9571
rect 25087 9537 25096 9571
rect 25044 9528 25096 9537
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 25688 9528 25740 9580
rect 25964 9528 26016 9580
rect 22468 9392 22520 9444
rect 22560 9392 22612 9444
rect 26148 9503 26200 9512
rect 26148 9469 26157 9503
rect 26157 9469 26191 9503
rect 26191 9469 26200 9503
rect 26148 9460 26200 9469
rect 24216 9367 24268 9376
rect 24216 9333 24225 9367
rect 24225 9333 24259 9367
rect 24259 9333 24268 9367
rect 24216 9324 24268 9333
rect 4664 9222 4716 9274
rect 4728 9222 4780 9274
rect 4792 9222 4844 9274
rect 4856 9222 4908 9274
rect 4920 9222 4972 9274
rect 12092 9222 12144 9274
rect 12156 9222 12208 9274
rect 12220 9222 12272 9274
rect 12284 9222 12336 9274
rect 12348 9222 12400 9274
rect 19520 9222 19572 9274
rect 19584 9222 19636 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 26948 9222 27000 9274
rect 27012 9222 27064 9274
rect 27076 9222 27128 9274
rect 27140 9222 27192 9274
rect 27204 9222 27256 9274
rect 2596 9120 2648 9172
rect 3608 9120 3660 9172
rect 4160 9120 4212 9172
rect 4344 9120 4396 9172
rect 4896 9120 4948 9172
rect 5172 9120 5224 9172
rect 9496 9120 9548 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 13176 9120 13228 9172
rect 14556 9163 14608 9172
rect 14556 9129 14565 9163
rect 14565 9129 14599 9163
rect 14599 9129 14608 9163
rect 14556 9120 14608 9129
rect 14924 9120 14976 9172
rect 22928 9163 22980 9172
rect 22928 9129 22937 9163
rect 22937 9129 22971 9163
rect 22971 9129 22980 9163
rect 22928 9120 22980 9129
rect 25044 9120 25096 9172
rect 3424 8916 3476 8968
rect 4528 8916 4580 8968
rect 5356 8984 5408 9036
rect 6184 8984 6236 9036
rect 12440 9052 12492 9104
rect 8300 8984 8352 9036
rect 11336 8984 11388 9036
rect 13084 9052 13136 9104
rect 3976 8848 4028 8900
rect 4988 8959 5040 8968
rect 4988 8925 4997 8959
rect 4997 8925 5031 8959
rect 5031 8925 5040 8959
rect 4988 8916 5040 8925
rect 5080 8916 5132 8968
rect 5172 8848 5224 8900
rect 5356 8848 5408 8900
rect 4988 8780 5040 8832
rect 5448 8780 5500 8832
rect 9312 8916 9364 8968
rect 9680 8916 9732 8968
rect 15476 9052 15528 9104
rect 25412 9095 25464 9104
rect 20812 8984 20864 9036
rect 25412 9061 25421 9095
rect 25421 9061 25455 9095
rect 25455 9061 25464 9095
rect 25412 9052 25464 9061
rect 22008 8984 22060 9036
rect 26148 9120 26200 9172
rect 12716 8916 12768 8968
rect 14188 8916 14240 8968
rect 14372 8916 14424 8968
rect 15200 8959 15252 8968
rect 15200 8925 15209 8959
rect 15209 8925 15243 8959
rect 15243 8925 15252 8959
rect 15200 8916 15252 8925
rect 7656 8891 7708 8900
rect 7656 8857 7665 8891
rect 7665 8857 7699 8891
rect 7699 8857 7708 8891
rect 7656 8848 7708 8857
rect 11888 8848 11940 8900
rect 16764 8848 16816 8900
rect 18420 8916 18472 8968
rect 21732 8959 21784 8968
rect 21732 8925 21741 8959
rect 21741 8925 21775 8959
rect 21775 8925 21784 8959
rect 21732 8916 21784 8925
rect 22376 8916 22428 8968
rect 25780 8959 25832 8968
rect 25780 8925 25789 8959
rect 25789 8925 25823 8959
rect 25823 8925 25832 8959
rect 25780 8916 25832 8925
rect 22928 8848 22980 8900
rect 25872 8848 25924 8900
rect 7564 8780 7616 8832
rect 10508 8780 10560 8832
rect 12532 8780 12584 8832
rect 12716 8780 12768 8832
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 16580 8780 16632 8832
rect 18144 8780 18196 8832
rect 25136 8780 25188 8832
rect 5324 8678 5376 8730
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 12752 8678 12804 8730
rect 12816 8678 12868 8730
rect 12880 8678 12932 8730
rect 12944 8678 12996 8730
rect 13008 8678 13060 8730
rect 20180 8678 20232 8730
rect 20244 8678 20296 8730
rect 20308 8678 20360 8730
rect 20372 8678 20424 8730
rect 20436 8678 20488 8730
rect 27608 8678 27660 8730
rect 27672 8678 27724 8730
rect 27736 8678 27788 8730
rect 27800 8678 27852 8730
rect 27864 8678 27916 8730
rect 8300 8576 8352 8628
rect 10784 8576 10836 8628
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 14188 8576 14240 8628
rect 15200 8576 15252 8628
rect 7196 8440 7248 8492
rect 7564 8440 7616 8492
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8760 8508 8812 8560
rect 9496 8508 9548 8560
rect 9680 8508 9732 8560
rect 6368 8304 6420 8356
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 7380 8236 7432 8288
rect 9220 8440 9272 8492
rect 8760 8347 8812 8356
rect 8760 8313 8769 8347
rect 8769 8313 8803 8347
rect 8803 8313 8812 8347
rect 8760 8304 8812 8313
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 10968 8440 11020 8492
rect 11336 8440 11388 8492
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 13636 8440 13688 8492
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 15476 8508 15528 8560
rect 16764 8508 16816 8560
rect 14372 8440 14424 8449
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 10876 8372 10928 8424
rect 14556 8372 14608 8424
rect 15844 8372 15896 8424
rect 16396 8483 16448 8492
rect 16396 8449 16405 8483
rect 16405 8449 16439 8483
rect 16439 8449 16448 8483
rect 16396 8440 16448 8449
rect 21732 8576 21784 8628
rect 17960 8508 18012 8560
rect 20536 8508 20588 8560
rect 22744 8576 22796 8628
rect 23388 8619 23440 8628
rect 23388 8585 23397 8619
rect 23397 8585 23431 8619
rect 23431 8585 23440 8619
rect 23388 8576 23440 8585
rect 24584 8619 24636 8628
rect 24584 8585 24593 8619
rect 24593 8585 24627 8619
rect 24627 8585 24636 8619
rect 24584 8576 24636 8585
rect 24768 8576 24820 8628
rect 25596 8576 25648 8628
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 10600 8304 10652 8356
rect 11244 8304 11296 8356
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 18144 8415 18196 8424
rect 18144 8381 18153 8415
rect 18153 8381 18187 8415
rect 18187 8381 18196 8415
rect 18144 8372 18196 8381
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 20812 8415 20864 8424
rect 20812 8381 20821 8415
rect 20821 8381 20855 8415
rect 20855 8381 20864 8415
rect 20812 8372 20864 8381
rect 22376 8415 22428 8424
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 23388 8372 23440 8424
rect 17316 8304 17368 8356
rect 18420 8304 18472 8356
rect 25136 8483 25188 8492
rect 25136 8449 25145 8483
rect 25145 8449 25179 8483
rect 25179 8449 25188 8483
rect 25136 8440 25188 8449
rect 25412 8440 25464 8492
rect 25872 8440 25924 8492
rect 8944 8279 8996 8288
rect 8944 8245 8953 8279
rect 8953 8245 8987 8279
rect 8987 8245 8996 8279
rect 8944 8236 8996 8245
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9220 8236 9272 8288
rect 9404 8236 9456 8288
rect 14556 8236 14608 8288
rect 16580 8236 16632 8288
rect 16764 8279 16816 8288
rect 16764 8245 16773 8279
rect 16773 8245 16807 8279
rect 16807 8245 16816 8279
rect 16764 8236 16816 8245
rect 19800 8236 19852 8288
rect 20260 8236 20312 8288
rect 22008 8279 22060 8288
rect 22008 8245 22017 8279
rect 22017 8245 22051 8279
rect 22051 8245 22060 8279
rect 22008 8236 22060 8245
rect 24676 8304 24728 8356
rect 25688 8347 25740 8356
rect 25688 8313 25697 8347
rect 25697 8313 25731 8347
rect 25731 8313 25740 8347
rect 25688 8304 25740 8313
rect 25320 8236 25372 8288
rect 4664 8134 4716 8186
rect 4728 8134 4780 8186
rect 4792 8134 4844 8186
rect 4856 8134 4908 8186
rect 4920 8134 4972 8186
rect 12092 8134 12144 8186
rect 12156 8134 12208 8186
rect 12220 8134 12272 8186
rect 12284 8134 12336 8186
rect 12348 8134 12400 8186
rect 19520 8134 19572 8186
rect 19584 8134 19636 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 26948 8134 27000 8186
rect 27012 8134 27064 8186
rect 27076 8134 27128 8186
rect 27140 8134 27192 8186
rect 27204 8134 27256 8186
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7564 8032 7616 8084
rect 8208 8032 8260 8084
rect 8852 8032 8904 8084
rect 9404 8032 9456 8084
rect 10692 8032 10744 8084
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 12440 8032 12492 8084
rect 15292 8032 15344 8084
rect 16028 8032 16080 8084
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17960 8075 18012 8084
rect 17960 8041 17969 8075
rect 17969 8041 18003 8075
rect 18003 8041 18012 8075
rect 17960 8032 18012 8041
rect 4068 7964 4120 8016
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 8116 7964 8168 8016
rect 8760 7964 8812 8016
rect 5724 7896 5776 7948
rect 6920 7896 6972 7948
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5172 7871 5224 7880
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 7380 7828 7432 7880
rect 9220 7896 9272 7948
rect 9312 7896 9364 7948
rect 9496 7828 9548 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 18788 8032 18840 8084
rect 19892 8032 19944 8084
rect 7196 7760 7248 7812
rect 9128 7803 9180 7812
rect 9128 7769 9137 7803
rect 9137 7769 9171 7803
rect 9171 7769 9180 7803
rect 9128 7760 9180 7769
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 10968 7828 11020 7837
rect 12624 7896 12676 7948
rect 16028 7896 16080 7948
rect 17224 7896 17276 7948
rect 18052 7896 18104 7948
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 16764 7828 16816 7880
rect 11980 7760 12032 7812
rect 15384 7760 15436 7812
rect 6368 7692 6420 7744
rect 9404 7735 9456 7744
rect 9404 7701 9413 7735
rect 9413 7701 9447 7735
rect 9447 7701 9456 7735
rect 9404 7692 9456 7701
rect 10048 7735 10100 7744
rect 10048 7701 10057 7735
rect 10057 7701 10091 7735
rect 10091 7701 10100 7735
rect 10048 7692 10100 7701
rect 10508 7692 10560 7744
rect 10784 7692 10836 7744
rect 13820 7692 13872 7744
rect 18328 7692 18380 7744
rect 18788 7896 18840 7948
rect 19800 7896 19852 7948
rect 20260 7896 20312 7948
rect 22008 8032 22060 8084
rect 25964 8032 26016 8084
rect 22376 7964 22428 8016
rect 22652 7964 22704 8016
rect 25596 7964 25648 8016
rect 19432 7828 19484 7880
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 20076 7828 20128 7880
rect 20812 7828 20864 7880
rect 24676 7828 24728 7880
rect 20720 7760 20772 7812
rect 25044 7760 25096 7812
rect 25412 7803 25464 7812
rect 25412 7769 25421 7803
rect 25421 7769 25455 7803
rect 25455 7769 25464 7803
rect 25412 7760 25464 7769
rect 19708 7692 19760 7744
rect 19984 7692 20036 7744
rect 5324 7590 5376 7642
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 12752 7590 12804 7642
rect 12816 7590 12868 7642
rect 12880 7590 12932 7642
rect 12944 7590 12996 7642
rect 13008 7590 13060 7642
rect 20180 7590 20232 7642
rect 20244 7590 20296 7642
rect 20308 7590 20360 7642
rect 20372 7590 20424 7642
rect 20436 7590 20488 7642
rect 27608 7590 27660 7642
rect 27672 7590 27724 7642
rect 27736 7590 27788 7642
rect 27800 7590 27852 7642
rect 27864 7590 27916 7642
rect 3792 7488 3844 7540
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 5724 7488 5776 7540
rect 7196 7488 7248 7540
rect 4160 7420 4212 7472
rect 9404 7488 9456 7540
rect 10048 7488 10100 7540
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 3332 7284 3384 7336
rect 6276 7284 6328 7336
rect 4068 7148 4120 7200
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 9036 7352 9088 7404
rect 10784 7352 10836 7404
rect 15936 7531 15988 7540
rect 15936 7497 15945 7531
rect 15945 7497 15979 7531
rect 15979 7497 15988 7531
rect 15936 7488 15988 7497
rect 16580 7488 16632 7540
rect 11152 7352 11204 7404
rect 11612 7352 11664 7404
rect 11980 7352 12032 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 13360 7395 13412 7404
rect 13360 7361 13395 7395
rect 13395 7361 13412 7395
rect 13360 7352 13412 7361
rect 13912 7352 13964 7404
rect 13728 7284 13780 7336
rect 14556 7352 14608 7404
rect 14096 7216 14148 7268
rect 8944 7148 8996 7200
rect 12716 7148 12768 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 12808 7148 12860 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13176 7148 13228 7200
rect 14464 7148 14516 7200
rect 15292 7284 15344 7336
rect 15476 7352 15528 7404
rect 15660 7352 15712 7404
rect 15568 7216 15620 7268
rect 15292 7148 15344 7200
rect 18052 7488 18104 7540
rect 20076 7488 20128 7540
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 20720 7488 20772 7540
rect 24216 7488 24268 7540
rect 24676 7488 24728 7540
rect 25044 7531 25096 7540
rect 25044 7497 25053 7531
rect 25053 7497 25087 7531
rect 25087 7497 25096 7531
rect 25044 7488 25096 7497
rect 25596 7531 25648 7540
rect 25596 7497 25605 7531
rect 25605 7497 25639 7531
rect 25639 7497 25648 7531
rect 25596 7488 25648 7497
rect 18328 7352 18380 7404
rect 18788 7352 18840 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 19800 7352 19852 7404
rect 22376 7420 22428 7472
rect 22008 7352 22060 7404
rect 24584 7395 24636 7404
rect 24584 7361 24593 7395
rect 24593 7361 24627 7395
rect 24627 7361 24636 7395
rect 24584 7352 24636 7361
rect 20168 7284 20220 7336
rect 23020 7327 23072 7336
rect 17960 7191 18012 7200
rect 17960 7157 17969 7191
rect 17969 7157 18003 7191
rect 18003 7157 18012 7191
rect 17960 7148 18012 7157
rect 19892 7148 19944 7200
rect 20260 7148 20312 7200
rect 23020 7293 23029 7327
rect 23029 7293 23063 7327
rect 23063 7293 23072 7327
rect 23020 7284 23072 7293
rect 22928 7216 22980 7268
rect 23664 7191 23716 7200
rect 23664 7157 23673 7191
rect 23673 7157 23707 7191
rect 23707 7157 23716 7191
rect 23664 7148 23716 7157
rect 4664 7046 4716 7098
rect 4728 7046 4780 7098
rect 4792 7046 4844 7098
rect 4856 7046 4908 7098
rect 4920 7046 4972 7098
rect 12092 7046 12144 7098
rect 12156 7046 12208 7098
rect 12220 7046 12272 7098
rect 12284 7046 12336 7098
rect 12348 7046 12400 7098
rect 19520 7046 19572 7098
rect 19584 7046 19636 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 26948 7046 27000 7098
rect 27012 7046 27064 7098
rect 27076 7046 27128 7098
rect 27140 7046 27192 7098
rect 27204 7046 27256 7098
rect 4988 6944 5040 6996
rect 3976 6876 4028 6928
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 12716 6944 12768 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 13268 6987 13320 6996
rect 13268 6953 13277 6987
rect 13277 6953 13311 6987
rect 13311 6953 13320 6987
rect 13268 6944 13320 6953
rect 13820 6944 13872 6996
rect 14924 6944 14976 6996
rect 16396 6944 16448 6996
rect 8300 6808 8352 6860
rect 11704 6808 11756 6860
rect 9312 6740 9364 6792
rect 6092 6604 6144 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 12900 6740 12952 6792
rect 13912 6876 13964 6928
rect 15200 6808 15252 6860
rect 15844 6851 15896 6860
rect 15844 6817 15853 6851
rect 15853 6817 15887 6851
rect 15887 6817 15896 6851
rect 20260 6944 20312 6996
rect 17960 6876 18012 6928
rect 15844 6808 15896 6817
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18788 6808 18840 6860
rect 21364 6851 21416 6860
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 21916 6808 21968 6860
rect 22836 6808 22888 6860
rect 23020 6808 23072 6860
rect 13728 6783 13780 6792
rect 13728 6749 13773 6783
rect 13773 6749 13780 6783
rect 13728 6740 13780 6749
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 7472 6604 7524 6656
rect 9496 6604 9548 6656
rect 11244 6672 11296 6724
rect 10692 6604 10744 6656
rect 11520 6647 11572 6656
rect 11520 6613 11529 6647
rect 11529 6613 11563 6647
rect 11563 6613 11572 6647
rect 11520 6604 11572 6613
rect 12808 6672 12860 6724
rect 13268 6672 13320 6724
rect 13452 6604 13504 6656
rect 13636 6715 13688 6724
rect 13636 6681 13645 6715
rect 13645 6681 13679 6715
rect 13679 6681 13688 6715
rect 13636 6672 13688 6681
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 15292 6783 15344 6792
rect 15292 6749 15301 6783
rect 15301 6749 15335 6783
rect 15335 6749 15344 6783
rect 15292 6740 15344 6749
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 15476 6672 15528 6724
rect 19432 6740 19484 6792
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20076 6672 20128 6724
rect 23664 6740 23716 6792
rect 16396 6647 16448 6656
rect 16396 6613 16405 6647
rect 16405 6613 16439 6647
rect 16439 6613 16448 6647
rect 16396 6604 16448 6613
rect 17776 6604 17828 6656
rect 21364 6604 21416 6656
rect 23572 6604 23624 6656
rect 23848 6604 23900 6656
rect 5324 6502 5376 6554
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 12752 6502 12804 6554
rect 12816 6502 12868 6554
rect 12880 6502 12932 6554
rect 12944 6502 12996 6554
rect 13008 6502 13060 6554
rect 20180 6502 20232 6554
rect 20244 6502 20296 6554
rect 20308 6502 20360 6554
rect 20372 6502 20424 6554
rect 20436 6502 20488 6554
rect 27608 6502 27660 6554
rect 27672 6502 27724 6554
rect 27736 6502 27788 6554
rect 27800 6502 27852 6554
rect 27864 6502 27916 6554
rect 9312 6400 9364 6452
rect 10600 6400 10652 6452
rect 11244 6400 11296 6452
rect 11520 6400 11572 6452
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 8392 6196 8444 6205
rect 11152 6264 11204 6316
rect 13728 6400 13780 6452
rect 15384 6400 15436 6452
rect 16028 6400 16080 6452
rect 15568 6264 15620 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16396 6264 16448 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 18420 6264 18472 6316
rect 20168 6332 20220 6384
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 22560 6332 22612 6384
rect 23848 6400 23900 6452
rect 24676 6400 24728 6452
rect 24400 6332 24452 6384
rect 9128 6128 9180 6180
rect 9496 6060 9548 6112
rect 14832 6196 14884 6248
rect 15292 6196 15344 6248
rect 11244 6171 11296 6180
rect 11244 6137 11253 6171
rect 11253 6137 11287 6171
rect 11287 6137 11296 6171
rect 11244 6128 11296 6137
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 20536 6128 20588 6180
rect 23572 6171 23624 6180
rect 23572 6137 23581 6171
rect 23581 6137 23615 6171
rect 23615 6137 23624 6171
rect 24584 6196 24636 6248
rect 23572 6128 23624 6137
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 16304 6060 16356 6112
rect 4664 5958 4716 6010
rect 4728 5958 4780 6010
rect 4792 5958 4844 6010
rect 4856 5958 4908 6010
rect 4920 5958 4972 6010
rect 12092 5958 12144 6010
rect 12156 5958 12208 6010
rect 12220 5958 12272 6010
rect 12284 5958 12336 6010
rect 12348 5958 12400 6010
rect 19520 5958 19572 6010
rect 19584 5958 19636 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 26948 5958 27000 6010
rect 27012 5958 27064 6010
rect 27076 5958 27128 6010
rect 27140 5958 27192 6010
rect 27204 5958 27256 6010
rect 6092 5856 6144 5908
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 11244 5856 11296 5908
rect 4068 5720 4120 5772
rect 7012 5720 7064 5772
rect 11520 5720 11572 5772
rect 13360 5856 13412 5908
rect 14280 5856 14332 5908
rect 17776 5899 17828 5908
rect 13452 5788 13504 5840
rect 9128 5652 9180 5704
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 17776 5865 17785 5899
rect 17785 5865 17819 5899
rect 17819 5865 17828 5899
rect 17776 5856 17828 5865
rect 19432 5899 19484 5908
rect 19432 5865 19441 5899
rect 19441 5865 19475 5899
rect 19475 5865 19484 5899
rect 19432 5856 19484 5865
rect 20168 5856 20220 5908
rect 22560 5856 22612 5908
rect 24400 5856 24452 5908
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 16028 5763 16080 5772
rect 16028 5729 16037 5763
rect 16037 5729 16071 5763
rect 16071 5729 16080 5763
rect 16028 5720 16080 5729
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 18236 5652 18288 5704
rect 19892 5652 19944 5704
rect 6736 5584 6788 5636
rect 11520 5584 11572 5636
rect 13268 5584 13320 5636
rect 12256 5559 12308 5568
rect 12256 5525 12265 5559
rect 12265 5525 12299 5559
rect 12299 5525 12308 5559
rect 12256 5516 12308 5525
rect 13452 5516 13504 5568
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 14832 5559 14884 5568
rect 14832 5525 14841 5559
rect 14841 5525 14875 5559
rect 14875 5525 14884 5559
rect 14832 5516 14884 5525
rect 5324 5414 5376 5466
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 12752 5414 12804 5466
rect 12816 5414 12868 5466
rect 12880 5414 12932 5466
rect 12944 5414 12996 5466
rect 13008 5414 13060 5466
rect 20180 5414 20232 5466
rect 20244 5414 20296 5466
rect 20308 5414 20360 5466
rect 20372 5414 20424 5466
rect 20436 5414 20488 5466
rect 27608 5414 27660 5466
rect 27672 5414 27724 5466
rect 27736 5414 27788 5466
rect 27800 5414 27852 5466
rect 27864 5414 27916 5466
rect 11520 5312 11572 5364
rect 12532 5312 12584 5364
rect 11888 5176 11940 5228
rect 12256 5219 12308 5228
rect 12256 5185 12265 5219
rect 12265 5185 12299 5219
rect 12299 5185 12308 5219
rect 12256 5176 12308 5185
rect 13636 5312 13688 5364
rect 14096 5312 14148 5364
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 13452 5244 13504 5296
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 13268 5108 13320 5160
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 4664 4870 4716 4922
rect 4728 4870 4780 4922
rect 4792 4870 4844 4922
rect 4856 4870 4908 4922
rect 4920 4870 4972 4922
rect 12092 4870 12144 4922
rect 12156 4870 12208 4922
rect 12220 4870 12272 4922
rect 12284 4870 12336 4922
rect 12348 4870 12400 4922
rect 19520 4870 19572 4922
rect 19584 4870 19636 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 26948 4870 27000 4922
rect 27012 4870 27064 4922
rect 27076 4870 27128 4922
rect 27140 4870 27192 4922
rect 27204 4870 27256 4922
rect 5324 4326 5376 4378
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 12752 4326 12804 4378
rect 12816 4326 12868 4378
rect 12880 4326 12932 4378
rect 12944 4326 12996 4378
rect 13008 4326 13060 4378
rect 20180 4326 20232 4378
rect 20244 4326 20296 4378
rect 20308 4326 20360 4378
rect 20372 4326 20424 4378
rect 20436 4326 20488 4378
rect 27608 4326 27660 4378
rect 27672 4326 27724 4378
rect 27736 4326 27788 4378
rect 27800 4326 27852 4378
rect 27864 4326 27916 4378
rect 14832 4088 14884 4140
rect 16120 4088 16172 4140
rect 17408 4088 17460 4140
rect 18144 4088 18196 4140
rect 4664 3782 4716 3834
rect 4728 3782 4780 3834
rect 4792 3782 4844 3834
rect 4856 3782 4908 3834
rect 4920 3782 4972 3834
rect 12092 3782 12144 3834
rect 12156 3782 12208 3834
rect 12220 3782 12272 3834
rect 12284 3782 12336 3834
rect 12348 3782 12400 3834
rect 19520 3782 19572 3834
rect 19584 3782 19636 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 26948 3782 27000 3834
rect 27012 3782 27064 3834
rect 27076 3782 27128 3834
rect 27140 3782 27192 3834
rect 27204 3782 27256 3834
rect 5324 3238 5376 3290
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 12752 3238 12804 3290
rect 12816 3238 12868 3290
rect 12880 3238 12932 3290
rect 12944 3238 12996 3290
rect 13008 3238 13060 3290
rect 20180 3238 20232 3290
rect 20244 3238 20296 3290
rect 20308 3238 20360 3290
rect 20372 3238 20424 3290
rect 20436 3238 20488 3290
rect 27608 3238 27660 3290
rect 27672 3238 27724 3290
rect 27736 3238 27788 3290
rect 27800 3238 27852 3290
rect 27864 3238 27916 3290
rect 4664 2694 4716 2746
rect 4728 2694 4780 2746
rect 4792 2694 4844 2746
rect 4856 2694 4908 2746
rect 4920 2694 4972 2746
rect 12092 2694 12144 2746
rect 12156 2694 12208 2746
rect 12220 2694 12272 2746
rect 12284 2694 12336 2746
rect 12348 2694 12400 2746
rect 19520 2694 19572 2746
rect 19584 2694 19636 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 26948 2694 27000 2746
rect 27012 2694 27064 2746
rect 27076 2694 27128 2746
rect 27140 2694 27192 2746
rect 27204 2694 27256 2746
rect 5324 2150 5376 2202
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 12752 2150 12804 2202
rect 12816 2150 12868 2202
rect 12880 2150 12932 2202
rect 12944 2150 12996 2202
rect 13008 2150 13060 2202
rect 20180 2150 20232 2202
rect 20244 2150 20296 2202
rect 20308 2150 20360 2202
rect 20372 2150 20424 2202
rect 20436 2150 20488 2202
rect 27608 2150 27660 2202
rect 27672 2150 27724 2202
rect 27736 2150 27788 2202
rect 27800 2150 27852 2202
rect 27864 2150 27916 2202
<< metal2 >>
rect 12898 31200 12954 32000
rect 14830 31200 14886 32000
rect 15474 31200 15530 32000
rect 18050 31362 18106 32000
rect 18050 31334 18184 31362
rect 18050 31200 18106 31334
rect 12912 30002 12940 31200
rect 12912 29974 13124 30002
rect 5324 29404 5632 29413
rect 5324 29402 5330 29404
rect 5386 29402 5410 29404
rect 5466 29402 5490 29404
rect 5546 29402 5570 29404
rect 5626 29402 5632 29404
rect 5386 29350 5388 29402
rect 5568 29350 5570 29402
rect 5324 29348 5330 29350
rect 5386 29348 5410 29350
rect 5466 29348 5490 29350
rect 5546 29348 5570 29350
rect 5626 29348 5632 29350
rect 5324 29339 5632 29348
rect 12752 29404 13060 29413
rect 12752 29402 12758 29404
rect 12814 29402 12838 29404
rect 12894 29402 12918 29404
rect 12974 29402 12998 29404
rect 13054 29402 13060 29404
rect 12814 29350 12816 29402
rect 12996 29350 12998 29402
rect 12752 29348 12758 29350
rect 12814 29348 12838 29350
rect 12894 29348 12918 29350
rect 12974 29348 12998 29350
rect 13054 29348 13060 29350
rect 12752 29339 13060 29348
rect 13096 29306 13124 29974
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 4664 28860 4972 28869
rect 4664 28858 4670 28860
rect 4726 28858 4750 28860
rect 4806 28858 4830 28860
rect 4886 28858 4910 28860
rect 4966 28858 4972 28860
rect 4726 28806 4728 28858
rect 4908 28806 4910 28858
rect 4664 28804 4670 28806
rect 4726 28804 4750 28806
rect 4806 28804 4830 28806
rect 4886 28804 4910 28806
rect 4966 28804 4972 28806
rect 4664 28795 4972 28804
rect 12092 28860 12400 28869
rect 12092 28858 12098 28860
rect 12154 28858 12178 28860
rect 12234 28858 12258 28860
rect 12314 28858 12338 28860
rect 12394 28858 12400 28860
rect 12154 28806 12156 28858
rect 12336 28806 12338 28858
rect 12092 28804 12098 28806
rect 12154 28804 12178 28806
rect 12234 28804 12258 28806
rect 12314 28804 12338 28806
rect 12394 28804 12400 28806
rect 12092 28795 12400 28804
rect 5324 28316 5632 28325
rect 5324 28314 5330 28316
rect 5386 28314 5410 28316
rect 5466 28314 5490 28316
rect 5546 28314 5570 28316
rect 5626 28314 5632 28316
rect 5386 28262 5388 28314
rect 5568 28262 5570 28314
rect 5324 28260 5330 28262
rect 5386 28260 5410 28262
rect 5466 28260 5490 28262
rect 5546 28260 5570 28262
rect 5626 28260 5632 28262
rect 5324 28251 5632 28260
rect 12752 28316 13060 28325
rect 12752 28314 12758 28316
rect 12814 28314 12838 28316
rect 12894 28314 12918 28316
rect 12974 28314 12998 28316
rect 13054 28314 13060 28316
rect 12814 28262 12816 28314
rect 12996 28262 12998 28314
rect 12752 28260 12758 28262
rect 12814 28260 12838 28262
rect 12894 28260 12918 28262
rect 12974 28260 12998 28262
rect 13054 28260 13060 28262
rect 12752 28251 13060 28260
rect 4664 27772 4972 27781
rect 4664 27770 4670 27772
rect 4726 27770 4750 27772
rect 4806 27770 4830 27772
rect 4886 27770 4910 27772
rect 4966 27770 4972 27772
rect 4726 27718 4728 27770
rect 4908 27718 4910 27770
rect 4664 27716 4670 27718
rect 4726 27716 4750 27718
rect 4806 27716 4830 27718
rect 4886 27716 4910 27718
rect 4966 27716 4972 27718
rect 4664 27707 4972 27716
rect 12092 27772 12400 27781
rect 12092 27770 12098 27772
rect 12154 27770 12178 27772
rect 12234 27770 12258 27772
rect 12314 27770 12338 27772
rect 12394 27770 12400 27772
rect 12154 27718 12156 27770
rect 12336 27718 12338 27770
rect 12092 27716 12098 27718
rect 12154 27716 12178 27718
rect 12234 27716 12258 27718
rect 12314 27716 12338 27718
rect 12394 27716 12400 27718
rect 12092 27707 12400 27716
rect 5324 27228 5632 27237
rect 5324 27226 5330 27228
rect 5386 27226 5410 27228
rect 5466 27226 5490 27228
rect 5546 27226 5570 27228
rect 5626 27226 5632 27228
rect 5386 27174 5388 27226
rect 5568 27174 5570 27226
rect 5324 27172 5330 27174
rect 5386 27172 5410 27174
rect 5466 27172 5490 27174
rect 5546 27172 5570 27174
rect 5626 27172 5632 27174
rect 5324 27163 5632 27172
rect 12752 27228 13060 27237
rect 12752 27226 12758 27228
rect 12814 27226 12838 27228
rect 12894 27226 12918 27228
rect 12974 27226 12998 27228
rect 13054 27226 13060 27228
rect 12814 27174 12816 27226
rect 12996 27174 12998 27226
rect 12752 27172 12758 27174
rect 12814 27172 12838 27174
rect 12894 27172 12918 27174
rect 12974 27172 12998 27174
rect 13054 27172 13060 27174
rect 12752 27163 13060 27172
rect 4664 26684 4972 26693
rect 4664 26682 4670 26684
rect 4726 26682 4750 26684
rect 4806 26682 4830 26684
rect 4886 26682 4910 26684
rect 4966 26682 4972 26684
rect 4726 26630 4728 26682
rect 4908 26630 4910 26682
rect 4664 26628 4670 26630
rect 4726 26628 4750 26630
rect 4806 26628 4830 26630
rect 4886 26628 4910 26630
rect 4966 26628 4972 26630
rect 4664 26619 4972 26628
rect 12092 26684 12400 26693
rect 12092 26682 12098 26684
rect 12154 26682 12178 26684
rect 12234 26682 12258 26684
rect 12314 26682 12338 26684
rect 12394 26682 12400 26684
rect 12154 26630 12156 26682
rect 12336 26630 12338 26682
rect 12092 26628 12098 26630
rect 12154 26628 12178 26630
rect 12234 26628 12258 26630
rect 12314 26628 12338 26630
rect 12394 26628 12400 26630
rect 12092 26619 12400 26628
rect 5324 26140 5632 26149
rect 5324 26138 5330 26140
rect 5386 26138 5410 26140
rect 5466 26138 5490 26140
rect 5546 26138 5570 26140
rect 5626 26138 5632 26140
rect 5386 26086 5388 26138
rect 5568 26086 5570 26138
rect 5324 26084 5330 26086
rect 5386 26084 5410 26086
rect 5466 26084 5490 26086
rect 5546 26084 5570 26086
rect 5626 26084 5632 26086
rect 5324 26075 5632 26084
rect 12752 26140 13060 26149
rect 12752 26138 12758 26140
rect 12814 26138 12838 26140
rect 12894 26138 12918 26140
rect 12974 26138 12998 26140
rect 13054 26138 13060 26140
rect 12814 26086 12816 26138
rect 12996 26086 12998 26138
rect 12752 26084 12758 26086
rect 12814 26084 12838 26086
rect 12894 26084 12918 26086
rect 12974 26084 12998 26086
rect 13054 26084 13060 26086
rect 12752 26075 13060 26084
rect 3974 25936 4030 25945
rect 3974 25871 4030 25880
rect 12808 25900 12860 25906
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 952 21185 980 21286
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20641 1532 20742
rect 1490 20632 1546 20641
rect 1490 20567 1546 20576
rect 938 19816 994 19825
rect 938 19751 994 19760
rect 952 19718 980 19751
rect 940 19712 992 19718
rect 940 19654 992 19660
rect 1492 19168 1544 19174
rect 1490 19136 1492 19145
rect 1544 19136 1546 19145
rect 1490 19071 1546 19080
rect 940 18624 992 18630
rect 940 18566 992 18572
rect 952 18465 980 18566
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1688 15910 1716 21490
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 2516 18290 2544 20334
rect 2792 20058 2820 20334
rect 3896 20058 3924 20402
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3712 18766 3740 19790
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3160 18426 3188 18566
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3528 18358 3556 18566
rect 3712 18426 3740 18702
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3516 18352 3568 18358
rect 3516 18294 3568 18300
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 3700 18080 3752 18086
rect 3804 18034 3832 18702
rect 3752 18028 3832 18034
rect 3700 18022 3832 18028
rect 3712 18006 3832 18022
rect 3804 17678 3832 18006
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1872 14414 1900 15982
rect 2332 15706 2360 15982
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2700 15502 2728 16390
rect 3988 16182 4016 25871
rect 12808 25842 12860 25848
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 4664 25596 4972 25605
rect 4664 25594 4670 25596
rect 4726 25594 4750 25596
rect 4806 25594 4830 25596
rect 4886 25594 4910 25596
rect 4966 25594 4972 25596
rect 4726 25542 4728 25594
rect 4908 25542 4910 25594
rect 4664 25540 4670 25542
rect 4726 25540 4750 25542
rect 4806 25540 4830 25542
rect 4886 25540 4910 25542
rect 4966 25540 4972 25542
rect 4664 25531 4972 25540
rect 10888 25362 10916 25774
rect 12092 25596 12400 25605
rect 12092 25594 12098 25596
rect 12154 25594 12178 25596
rect 12234 25594 12258 25596
rect 12314 25594 12338 25596
rect 12394 25594 12400 25596
rect 12154 25542 12156 25594
rect 12336 25542 12338 25594
rect 12092 25540 12098 25542
rect 12154 25540 12178 25542
rect 12234 25540 12258 25542
rect 12314 25540 12338 25542
rect 12394 25540 12400 25542
rect 12092 25531 12400 25540
rect 12820 25498 12848 25842
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 13004 25498 13032 25638
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 5324 25052 5632 25061
rect 5324 25050 5330 25052
rect 5386 25050 5410 25052
rect 5466 25050 5490 25052
rect 5546 25050 5570 25052
rect 5626 25050 5632 25052
rect 5386 24998 5388 25050
rect 5568 24998 5570 25050
rect 5324 24996 5330 24998
rect 5386 24996 5410 24998
rect 5466 24996 5490 24998
rect 5546 24996 5570 24998
rect 5626 24996 5632 24998
rect 5324 24987 5632 24996
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6460 24608 6512 24614
rect 6460 24550 6512 24556
rect 4664 24508 4972 24517
rect 4664 24506 4670 24508
rect 4726 24506 4750 24508
rect 4806 24506 4830 24508
rect 4886 24506 4910 24508
rect 4966 24506 4972 24508
rect 4726 24454 4728 24506
rect 4908 24454 4910 24506
rect 4664 24452 4670 24454
rect 4726 24452 4750 24454
rect 4806 24452 4830 24454
rect 4886 24452 4910 24454
rect 4966 24452 4972 24454
rect 4664 24443 4972 24452
rect 6472 24274 6500 24550
rect 6656 24410 6684 24686
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 7944 24206 7972 24550
rect 8404 24410 8432 24754
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8496 24342 8524 25094
rect 9416 24886 9444 25094
rect 10888 24954 10916 25298
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 10980 24954 11008 25162
rect 11900 24954 11928 25162
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 12360 24818 12388 25094
rect 12752 25052 13060 25061
rect 12752 25050 12758 25052
rect 12814 25050 12838 25052
rect 12894 25050 12918 25052
rect 12974 25050 12998 25052
rect 13054 25050 13060 25052
rect 12814 24998 12816 25050
rect 12996 24998 12998 25050
rect 12752 24996 12758 24998
rect 12814 24996 12838 24998
rect 12894 24996 12918 24998
rect 12974 24996 12998 24998
rect 13054 24996 13060 24998
rect 12752 24987 13060 24996
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 9312 24744 9364 24750
rect 9232 24704 9312 24732
rect 8484 24336 8536 24342
rect 8404 24284 8484 24290
rect 8404 24278 8536 24284
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8404 24262 8524 24278
rect 7104 24200 7156 24206
rect 7104 24142 7156 24148
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6920 24132 6972 24138
rect 6920 24074 6972 24080
rect 4448 23066 4476 24074
rect 5324 23964 5632 23973
rect 5324 23962 5330 23964
rect 5386 23962 5410 23964
rect 5466 23962 5490 23964
rect 5546 23962 5570 23964
rect 5626 23962 5632 23964
rect 5386 23910 5388 23962
rect 5568 23910 5570 23962
rect 5324 23908 5330 23910
rect 5386 23908 5410 23910
rect 5466 23908 5490 23910
rect 5546 23908 5570 23910
rect 5626 23908 5632 23910
rect 5324 23899 5632 23908
rect 5736 23866 5764 24074
rect 6196 23866 6224 24074
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 4664 23420 4972 23429
rect 4664 23418 4670 23420
rect 4726 23418 4750 23420
rect 4806 23418 4830 23420
rect 4886 23418 4910 23420
rect 4966 23418 4972 23420
rect 4726 23366 4728 23418
rect 4908 23366 4910 23418
rect 4664 23364 4670 23366
rect 4726 23364 4750 23366
rect 4806 23364 4830 23366
rect 4886 23364 4910 23366
rect 4966 23364 4972 23366
rect 4664 23355 4972 23364
rect 6564 23322 6592 23666
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 4448 23038 4568 23066
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4172 22234 4200 22510
rect 4160 22228 4212 22234
rect 4160 22170 4212 22176
rect 4448 22098 4476 22714
rect 4436 22092 4488 22098
rect 4436 22034 4488 22040
rect 4344 22024 4396 22030
rect 4344 21966 4396 21972
rect 4356 21690 4384 21966
rect 4540 21894 4568 23038
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 5324 22876 5632 22885
rect 5324 22874 5330 22876
rect 5386 22874 5410 22876
rect 5466 22874 5490 22876
rect 5546 22874 5570 22876
rect 5626 22874 5632 22876
rect 5386 22822 5388 22874
rect 5568 22822 5570 22874
rect 5324 22820 5330 22822
rect 5386 22820 5410 22822
rect 5466 22820 5490 22822
rect 5546 22820 5570 22822
rect 5626 22820 5632 22822
rect 5324 22811 5632 22820
rect 5172 22704 5224 22710
rect 5172 22646 5224 22652
rect 6092 22704 6144 22710
rect 6092 22646 6144 22652
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4664 22332 4972 22341
rect 4664 22330 4670 22332
rect 4726 22330 4750 22332
rect 4806 22330 4830 22332
rect 4886 22330 4910 22332
rect 4966 22330 4972 22332
rect 4726 22278 4728 22330
rect 4908 22278 4910 22330
rect 4664 22276 4670 22278
rect 4726 22276 4750 22278
rect 4806 22276 4830 22278
rect 4886 22276 4910 22278
rect 4966 22276 4972 22278
rect 4664 22267 4972 22276
rect 5000 22234 5028 22374
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 5092 22094 5120 22374
rect 5184 22098 5212 22646
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 5920 22234 5948 22578
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5000 22066 5120 22094
rect 5172 22092 5224 22098
rect 5000 22030 5028 22066
rect 5172 22034 5224 22040
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4528 21888 4580 21894
rect 4528 21830 4580 21836
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4448 21350 4476 21830
rect 4540 21622 4568 21830
rect 4528 21616 4580 21622
rect 4528 21558 4580 21564
rect 4632 21434 4660 21830
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 4540 21406 4660 21434
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4172 20398 4200 20878
rect 4264 20602 4292 20878
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 17338 4108 17546
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 4080 16114 4108 17070
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16250 4200 16390
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 2964 14816 3016 14822
rect 2964 14758 3016 14764
rect 1860 14408 1912 14414
rect 938 14376 994 14385
rect 1860 14350 1912 14356
rect 938 14311 994 14320
rect 952 13938 980 14311
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 13938 1716 14214
rect 940 13932 992 13938
rect 940 13874 992 13880
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1872 12782 1900 14350
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 14074 2176 14282
rect 2976 14074 3004 14758
rect 3528 14618 3556 14962
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14074 3188 14282
rect 3528 14074 3556 14554
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3620 13802 3648 16050
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3608 13796 3660 13802
rect 3608 13738 3660 13744
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 12306 1900 12718
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12306 2636 12582
rect 2792 12442 2820 12786
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 1872 11354 1900 12242
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11898 3280 12174
rect 3620 11898 3648 13738
rect 3804 12238 3832 14894
rect 4080 14822 4108 14991
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3896 14278 3924 14758
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3988 13734 4016 14350
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4080 13938 4108 14214
rect 4172 13938 4200 14214
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3976 13728 4028 13734
rect 4068 13728 4120 13734
rect 3976 13670 4028 13676
rect 4066 13696 4068 13705
rect 4120 13696 4122 13705
rect 3988 12918 4016 13670
rect 4066 13631 4122 13640
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3988 12434 4016 12854
rect 4172 12850 4200 13874
rect 4264 13326 4292 20402
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4356 20058 4384 20198
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4448 19938 4476 21286
rect 4540 20890 4568 21406
rect 4664 21244 4972 21253
rect 4664 21242 4670 21244
rect 4726 21242 4750 21244
rect 4806 21242 4830 21244
rect 4886 21242 4910 21244
rect 4966 21242 4972 21244
rect 4726 21190 4728 21242
rect 4908 21190 4910 21242
rect 4664 21188 4670 21190
rect 4726 21188 4750 21190
rect 4806 21188 4830 21190
rect 4886 21188 4910 21190
rect 4966 21188 4972 21190
rect 4664 21179 4972 21188
rect 4540 20862 4660 20890
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20602 4568 20742
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4632 20534 4660 20862
rect 4620 20528 4672 20534
rect 4620 20470 4672 20476
rect 4664 20156 4972 20165
rect 4664 20154 4670 20156
rect 4726 20154 4750 20156
rect 4806 20154 4830 20156
rect 4886 20154 4910 20156
rect 4966 20154 4972 20156
rect 4726 20102 4728 20154
rect 4908 20102 4910 20154
rect 4664 20100 4670 20102
rect 4726 20100 4750 20102
rect 4806 20100 4830 20102
rect 4886 20100 4910 20102
rect 4966 20100 4972 20102
rect 4664 20091 4972 20100
rect 5000 20040 5028 21558
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5092 21146 5120 21286
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5092 20602 5120 20878
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 5184 20534 5212 22034
rect 5324 21788 5632 21797
rect 5324 21786 5330 21788
rect 5386 21786 5410 21788
rect 5466 21786 5490 21788
rect 5546 21786 5570 21788
rect 5626 21786 5632 21788
rect 5386 21734 5388 21786
rect 5568 21734 5570 21786
rect 5324 21732 5330 21734
rect 5386 21732 5410 21734
rect 5466 21732 5490 21734
rect 5546 21732 5570 21734
rect 5626 21732 5632 21734
rect 5324 21723 5632 21732
rect 6104 21554 6132 22646
rect 6564 22574 6592 22918
rect 6656 22778 6684 23122
rect 6932 22778 6960 24074
rect 7116 23798 7144 24142
rect 7104 23792 7156 23798
rect 7104 23734 7156 23740
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 7024 22982 7052 23666
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6920 22636 6972 22642
rect 7024 22624 7052 22918
rect 6972 22596 7052 22624
rect 6920 22578 6972 22584
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6748 21554 6776 22170
rect 6932 22094 6960 22578
rect 6840 22066 6960 22094
rect 6840 21690 6868 22066
rect 7116 21690 7144 23122
rect 7208 22642 7236 24142
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7852 23254 7880 23462
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7208 22098 7236 22578
rect 7484 22438 7512 22918
rect 7668 22778 7696 23054
rect 7852 22982 7880 23190
rect 7944 23118 7972 24142
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8128 23730 8156 24006
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7656 22772 7708 22778
rect 7656 22714 7708 22720
rect 7760 22642 7788 22918
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 8036 22574 8064 23190
rect 8220 23118 8248 23462
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 5552 20942 5580 21490
rect 6104 21078 6132 21490
rect 6564 21146 6592 21490
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6840 21078 6868 21286
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 6828 21072 6880 21078
rect 6828 21014 6880 21020
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 6460 20936 6512 20942
rect 6736 20936 6788 20942
rect 6460 20878 6512 20884
rect 6656 20896 6736 20924
rect 5324 20700 5632 20709
rect 5324 20698 5330 20700
rect 5386 20698 5410 20700
rect 5466 20698 5490 20700
rect 5546 20698 5570 20700
rect 5626 20698 5632 20700
rect 5386 20646 5388 20698
rect 5568 20646 5570 20698
rect 5324 20644 5330 20646
rect 5386 20644 5410 20646
rect 5466 20644 5490 20646
rect 5546 20644 5570 20646
rect 5626 20644 5632 20646
rect 5324 20635 5632 20644
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 6472 20466 6500 20878
rect 6656 20806 6684 20896
rect 6736 20878 6788 20884
rect 6840 20856 6868 21014
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 6920 20868 6972 20874
rect 6840 20828 6920 20856
rect 6920 20810 6972 20816
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 7024 20602 7052 20946
rect 7576 20602 7604 20946
rect 7668 20806 7696 21626
rect 8220 21622 8248 23054
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 8220 20806 8248 21558
rect 8312 21434 8340 24210
rect 8404 24138 8432 24262
rect 9232 24206 9260 24704
rect 9312 24686 9364 24692
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9220 24200 9272 24206
rect 9220 24142 9272 24148
rect 8392 24132 8444 24138
rect 8392 24074 8444 24080
rect 9036 24132 9088 24138
rect 9036 24074 9088 24080
rect 9128 24132 9180 24138
rect 9128 24074 9180 24080
rect 8404 23798 8432 24074
rect 8392 23792 8444 23798
rect 8392 23734 8444 23740
rect 9048 23730 9076 24074
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8496 22642 8524 22918
rect 9140 22778 9168 24074
rect 9232 23118 9260 24142
rect 9692 23338 9720 24550
rect 10060 24410 10088 24686
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 10336 24274 10364 24686
rect 10416 24676 10468 24682
rect 10416 24618 10468 24624
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10428 23594 10456 24618
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10416 23588 10468 23594
rect 10416 23530 10468 23536
rect 9600 23322 9720 23338
rect 9588 23316 9720 23322
rect 9640 23310 9720 23316
rect 9588 23258 9640 23264
rect 9220 23112 9272 23118
rect 9220 23054 9272 23060
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8404 22094 8432 22578
rect 8588 22234 8616 22578
rect 8680 22234 8708 22578
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8404 22066 8616 22094
rect 8312 21406 8524 21434
rect 8496 21350 8524 21406
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7668 20466 7696 20742
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 4356 19910 4476 19938
rect 4908 20012 5028 20040
rect 4356 18630 4384 19910
rect 4908 19718 4936 20012
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4724 19514 4752 19654
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 5000 19310 5028 19858
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 4448 18698 4476 19110
rect 4540 18834 4568 19178
rect 4664 19068 4972 19077
rect 4664 19066 4670 19068
rect 4726 19066 4750 19068
rect 4806 19066 4830 19068
rect 4886 19066 4910 19068
rect 4966 19066 4972 19068
rect 4726 19014 4728 19066
rect 4908 19014 4910 19066
rect 4664 19012 4670 19014
rect 4726 19012 4750 19014
rect 4806 19012 4830 19014
rect 4886 19012 4910 19014
rect 4966 19012 4972 19014
rect 4664 19003 4972 19012
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4908 18306 4936 18566
rect 5000 18426 5028 19246
rect 5092 19242 5120 20334
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19922 5396 20198
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5552 19854 5580 20402
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5324 19612 5632 19621
rect 5324 19610 5330 19612
rect 5386 19610 5410 19612
rect 5466 19610 5490 19612
rect 5546 19610 5570 19612
rect 5626 19610 5632 19612
rect 5386 19558 5388 19610
rect 5568 19558 5570 19610
rect 5324 19556 5330 19558
rect 5386 19556 5410 19558
rect 5466 19556 5490 19558
rect 5546 19556 5570 19558
rect 5626 19556 5632 19558
rect 5324 19547 5632 19556
rect 6472 19514 6500 20402
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19514 6868 19654
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18630 5580 19110
rect 6092 18692 6144 18698
rect 6092 18634 6144 18640
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5324 18524 5632 18533
rect 5324 18522 5330 18524
rect 5386 18522 5410 18524
rect 5466 18522 5490 18524
rect 5546 18522 5570 18524
rect 5626 18522 5632 18524
rect 5386 18470 5388 18522
rect 5568 18470 5570 18522
rect 5324 18468 5330 18470
rect 5386 18468 5410 18470
rect 5466 18468 5490 18470
rect 5546 18468 5570 18470
rect 5626 18468 5632 18470
rect 5324 18459 5632 18468
rect 6104 18426 6132 18634
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 4908 18278 5028 18306
rect 4664 17980 4972 17989
rect 4664 17978 4670 17980
rect 4726 17978 4750 17980
rect 4806 17978 4830 17980
rect 4886 17978 4910 17980
rect 4966 17978 4972 17980
rect 4726 17926 4728 17978
rect 4908 17926 4910 17978
rect 4664 17924 4670 17926
rect 4726 17924 4750 17926
rect 4806 17924 4830 17926
rect 4886 17924 4910 17926
rect 4966 17924 4972 17926
rect 4664 17915 4972 17924
rect 4528 17604 4580 17610
rect 4528 17546 4580 17552
rect 4540 17338 4568 17546
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4356 16114 4384 17002
rect 4664 16892 4972 16901
rect 4664 16890 4670 16892
rect 4726 16890 4750 16892
rect 4806 16890 4830 16892
rect 4886 16890 4910 16892
rect 4966 16890 4972 16892
rect 4726 16838 4728 16890
rect 4908 16838 4910 16890
rect 4664 16836 4670 16838
rect 4726 16836 4750 16838
rect 4806 16836 4830 16838
rect 4886 16836 4910 16838
rect 4966 16836 4972 16838
rect 4664 16827 4972 16836
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4434 16416 4490 16425
rect 4434 16351 4490 16360
rect 4448 16114 4476 16351
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4342 15736 4398 15745
rect 4342 15671 4398 15680
rect 4356 15570 4384 15671
rect 4448 15570 4476 16050
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4540 14958 4568 16594
rect 5000 15910 5028 18278
rect 6472 17882 6500 19450
rect 7392 18970 7420 19858
rect 7668 19768 7696 20402
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7840 19780 7892 19786
rect 7668 19740 7840 19768
rect 7840 19722 7892 19728
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7484 18970 7512 19654
rect 7944 19446 7972 19994
rect 8036 19854 8064 20198
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8496 19514 8524 21286
rect 8588 21146 8616 22066
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8772 20534 8800 22578
rect 9232 22030 9260 23054
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9324 22098 9352 22918
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 22024 9272 22030
rect 9600 21978 9628 23258
rect 10520 22982 10548 23598
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10520 22778 10548 22918
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9220 21966 9272 21972
rect 9232 21690 9260 21966
rect 9416 21950 9628 21978
rect 9312 21888 9364 21894
rect 9416 21876 9444 21950
rect 9364 21848 9444 21876
rect 9496 21888 9548 21894
rect 9312 21830 9364 21836
rect 9496 21830 9548 21836
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9324 20874 9352 21830
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9312 20868 9364 20874
rect 9312 20810 9364 20816
rect 8760 20528 8812 20534
rect 8760 20470 8812 20476
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7576 18834 7604 19314
rect 8588 18970 8616 19382
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7668 18426 7696 18702
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6748 17882 6776 18158
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6472 17762 6500 17818
rect 6932 17814 6960 18022
rect 6380 17734 6500 17762
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5324 17436 5632 17445
rect 5324 17434 5330 17436
rect 5386 17434 5410 17436
rect 5466 17434 5490 17436
rect 5546 17434 5570 17436
rect 5626 17434 5632 17436
rect 5386 17382 5388 17434
rect 5568 17382 5570 17434
rect 5324 17380 5330 17382
rect 5386 17380 5410 17382
rect 5466 17380 5490 17382
rect 5546 17380 5570 17382
rect 5626 17380 5632 17382
rect 5324 17371 5632 17380
rect 5736 17338 5764 17614
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 6380 17202 6408 17734
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 5276 16794 5304 17070
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5276 16658 5304 16730
rect 6288 16726 6316 17070
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5184 16114 5212 16458
rect 5324 16348 5632 16357
rect 5324 16346 5330 16348
rect 5386 16346 5410 16348
rect 5466 16346 5490 16348
rect 5546 16346 5570 16348
rect 5626 16346 5632 16348
rect 5386 16294 5388 16346
rect 5568 16294 5570 16346
rect 5324 16292 5330 16294
rect 5386 16292 5410 16294
rect 5466 16292 5490 16294
rect 5546 16292 5570 16294
rect 5626 16292 5632 16294
rect 5324 16283 5632 16292
rect 5736 16114 5764 16662
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4664 15804 4972 15813
rect 4664 15802 4670 15804
rect 4726 15802 4750 15804
rect 4806 15802 4830 15804
rect 4886 15802 4910 15804
rect 4966 15802 4972 15804
rect 4726 15750 4728 15802
rect 4908 15750 4910 15802
rect 4664 15748 4670 15750
rect 4726 15748 4750 15750
rect 4806 15748 4830 15750
rect 4886 15748 4910 15750
rect 4966 15748 4972 15750
rect 4664 15739 4972 15748
rect 5184 15570 5212 16050
rect 6012 15706 6040 16050
rect 6196 15910 6224 16662
rect 6380 16046 6408 17138
rect 6472 16998 6500 17478
rect 6840 17338 6868 17614
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6104 15570 6132 15642
rect 6196 15570 6224 15846
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6472 15484 6500 16934
rect 6932 16658 6960 17138
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6564 16114 6592 16390
rect 6932 16250 6960 16594
rect 7024 16590 7052 18090
rect 7208 17610 7236 18226
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 7288 17808 7340 17814
rect 8312 17762 8340 17818
rect 8772 17762 8800 20470
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9048 19530 9076 19790
rect 9048 19502 9168 19530
rect 9140 19446 9168 19502
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 9324 19310 9352 19858
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 7288 17750 7340 17756
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 17202 7236 17546
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7300 16998 7328 17750
rect 8220 17734 8340 17762
rect 8220 17678 8248 17734
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 17338 7880 17478
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7944 17105 7972 17206
rect 8116 17128 8168 17134
rect 7930 17096 7986 17105
rect 8116 17070 8168 17076
rect 7930 17031 7986 17040
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6552 15496 6604 15502
rect 6472 15456 6552 15484
rect 6552 15438 6604 15444
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5324 15260 5632 15269
rect 5324 15258 5330 15260
rect 5386 15258 5410 15260
rect 5466 15258 5490 15260
rect 5546 15258 5570 15260
rect 5626 15258 5632 15260
rect 5386 15206 5388 15258
rect 5568 15206 5570 15258
rect 5324 15204 5330 15206
rect 5386 15204 5410 15206
rect 5466 15204 5490 15206
rect 5546 15204 5570 15206
rect 5626 15204 5632 15206
rect 5324 15195 5632 15204
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4664 14716 4972 14725
rect 4664 14714 4670 14716
rect 4726 14714 4750 14716
rect 4806 14714 4830 14716
rect 4886 14714 4910 14716
rect 4966 14714 4972 14716
rect 4726 14662 4728 14714
rect 4908 14662 4910 14714
rect 4664 14660 4670 14662
rect 4726 14660 4750 14662
rect 4806 14660 4830 14662
rect 4886 14660 4910 14662
rect 4966 14660 4972 14662
rect 4664 14651 4972 14660
rect 5736 14618 5764 15302
rect 6564 15094 6592 15438
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6656 14618 6684 15302
rect 6748 15162 6776 16050
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 6840 15434 6868 15506
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 7024 15094 7052 15506
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 4988 14544 5040 14550
rect 4988 14486 5040 14492
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4356 14074 4384 14350
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4540 12850 4568 14282
rect 4664 13628 4972 13637
rect 4664 13626 4670 13628
rect 4726 13626 4750 13628
rect 4806 13626 4830 13628
rect 4886 13626 4910 13628
rect 4966 13626 4972 13628
rect 4726 13574 4728 13626
rect 4908 13574 4910 13626
rect 4664 13572 4670 13574
rect 4726 13572 4750 13574
rect 4806 13572 4830 13574
rect 4886 13572 4910 13574
rect 4966 13572 4972 13574
rect 4664 13563 4972 13572
rect 5000 12850 5028 14486
rect 6748 14278 6776 14894
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 14414 6868 14554
rect 7116 14414 7144 15030
rect 7208 14958 7236 15506
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 5324 14172 5632 14181
rect 5324 14170 5330 14172
rect 5386 14170 5410 14172
rect 5466 14170 5490 14172
rect 5546 14170 5570 14172
rect 5626 14170 5632 14172
rect 5386 14118 5388 14170
rect 5568 14118 5570 14170
rect 5324 14116 5330 14118
rect 5386 14116 5410 14118
rect 5466 14116 5490 14118
rect 5546 14116 5570 14118
rect 5626 14116 5632 14118
rect 5324 14107 5632 14116
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13326 5580 13738
rect 6564 13326 6592 13874
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6656 13530 6684 13806
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 5324 13084 5632 13093
rect 5324 13082 5330 13084
rect 5386 13082 5410 13084
rect 5466 13082 5490 13084
rect 5546 13082 5570 13084
rect 5626 13082 5632 13084
rect 5386 13030 5388 13082
rect 5568 13030 5570 13082
rect 5324 13028 5330 13030
rect 5386 13028 5410 13030
rect 5466 13028 5490 13030
rect 5546 13028 5570 13030
rect 5626 13028 5632 13030
rect 5324 13019 5632 13028
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 3988 12406 4108 12434
rect 3974 12336 4030 12345
rect 3974 12271 3976 12280
rect 4028 12271 4030 12280
rect 3976 12242 4028 12248
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 2056 10810 2084 11018
rect 3160 10810 3188 11086
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3344 10674 3372 11698
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3974 10976 4030 10985
rect 3804 10810 3832 10950
rect 3974 10911 4030 10920
rect 3988 10810 4016 10911
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4080 10674 4108 12406
rect 4172 10674 4200 12786
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4356 11218 4384 12242
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3344 9674 3372 10610
rect 3344 9646 3464 9674
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 9178 2636 9454
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 3344 7342 3372 9318
rect 3436 8974 3464 9646
rect 3608 9648 3660 9654
rect 4068 9648 4120 9654
rect 3608 9590 3660 9596
rect 4066 9616 4068 9625
rect 4120 9616 4122 9625
rect 3620 9178 3648 9590
rect 4066 9551 4122 9560
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 9178 4200 9318
rect 4356 9178 4384 11154
rect 4540 10674 4568 12786
rect 4664 12540 4972 12549
rect 4664 12538 4670 12540
rect 4726 12538 4750 12540
rect 4806 12538 4830 12540
rect 4886 12538 4910 12540
rect 4966 12538 4972 12540
rect 4726 12486 4728 12538
rect 4908 12486 4910 12538
rect 4664 12484 4670 12486
rect 4726 12484 4750 12486
rect 4806 12484 4830 12486
rect 4886 12484 4910 12486
rect 4966 12484 4972 12486
rect 4664 12475 4972 12484
rect 4664 11452 4972 11461
rect 4664 11450 4670 11452
rect 4726 11450 4750 11452
rect 4806 11450 4830 11452
rect 4886 11450 4910 11452
rect 4966 11450 4972 11452
rect 4726 11398 4728 11450
rect 4908 11398 4910 11450
rect 4664 11396 4670 11398
rect 4726 11396 4750 11398
rect 4806 11396 4830 11398
rect 4886 11396 4910 11398
rect 4966 11396 4972 11398
rect 4664 11387 4972 11396
rect 5000 11200 5028 12786
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 12306 5120 12582
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5184 11898 5212 12242
rect 5324 11996 5632 12005
rect 5324 11994 5330 11996
rect 5386 11994 5410 11996
rect 5466 11994 5490 11996
rect 5546 11994 5570 11996
rect 5626 11994 5632 11996
rect 5386 11942 5388 11994
rect 5568 11942 5570 11994
rect 5324 11940 5330 11942
rect 5386 11940 5410 11942
rect 5466 11940 5490 11942
rect 5546 11940 5570 11942
rect 5626 11940 5632 11942
rect 5324 11931 5632 11940
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5736 11778 5764 13262
rect 7116 12986 7144 14350
rect 7208 13394 7236 14894
rect 7392 14498 7420 16934
rect 8128 16794 8156 17070
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 16114 8156 16390
rect 8312 16182 8340 17734
rect 8680 17734 8800 17762
rect 8852 17740 8904 17746
rect 8680 17678 8708 17734
rect 8852 17682 8904 17688
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8484 17604 8536 17610
rect 8536 17564 8616 17592
rect 8484 17546 8536 17552
rect 8588 16590 8616 17564
rect 8680 17542 8708 17614
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7300 14482 7420 14498
rect 7300 14476 7432 14482
rect 7300 14470 7380 14476
rect 7300 14074 7328 14470
rect 7380 14418 7432 14424
rect 7484 14414 7512 15846
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7484 14006 7512 14350
rect 8220 14346 8248 15030
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7760 13410 7788 14282
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 14006 7972 14214
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 8036 13938 8064 14282
rect 8128 14074 8156 14282
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7932 13864 7984 13870
rect 8116 13864 8168 13870
rect 7984 13812 8116 13818
rect 7932 13806 8168 13812
rect 7944 13790 8156 13806
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7392 13382 7788 13410
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6104 12434 6132 12650
rect 6104 12406 6224 12434
rect 5184 11750 5764 11778
rect 5184 11694 5212 11750
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 4816 11172 5028 11200
rect 4816 10674 4844 11172
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10742 4936 11018
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4540 8974 4568 10610
rect 4664 10364 4972 10373
rect 4664 10362 4670 10364
rect 4726 10362 4750 10364
rect 4806 10362 4830 10364
rect 4886 10362 4910 10364
rect 4966 10362 4972 10364
rect 4726 10310 4728 10362
rect 4908 10310 4910 10362
rect 4664 10308 4670 10310
rect 4726 10308 4750 10310
rect 4806 10308 4830 10310
rect 4886 10308 4910 10310
rect 4966 10308 4972 10310
rect 4664 10299 4972 10308
rect 4664 9276 4972 9285
rect 4664 9274 4670 9276
rect 4726 9274 4750 9276
rect 4806 9274 4830 9276
rect 4886 9274 4910 9276
rect 4966 9274 4972 9276
rect 4726 9222 4728 9274
rect 4908 9222 4910 9274
rect 4664 9220 4670 9222
rect 4726 9220 4750 9222
rect 4806 9220 4830 9222
rect 4886 9220 4910 9222
rect 4966 9220 4972 9222
rect 4664 9211 4972 9220
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3988 7834 4016 8842
rect 4908 8650 4936 9114
rect 5000 8974 5028 11172
rect 5184 10606 5212 11630
rect 6196 11626 6224 12406
rect 6472 12238 6500 12854
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11898 6500 12174
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11898 6960 12038
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5324 10908 5632 10917
rect 5324 10906 5330 10908
rect 5386 10906 5410 10908
rect 5466 10906 5490 10908
rect 5546 10906 5570 10908
rect 5626 10906 5632 10908
rect 5386 10854 5388 10906
rect 5568 10854 5570 10906
rect 5324 10852 5330 10854
rect 5386 10852 5410 10854
rect 5466 10852 5490 10854
rect 5546 10852 5570 10854
rect 5626 10852 5632 10854
rect 5324 10843 5632 10852
rect 5736 10742 5764 11018
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 6656 10674 6684 10950
rect 6840 10674 6868 11290
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 9568 5120 10474
rect 5184 10062 5212 10542
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 5324 9820 5632 9829
rect 5324 9818 5330 9820
rect 5386 9818 5410 9820
rect 5466 9818 5490 9820
rect 5546 9818 5570 9820
rect 5626 9818 5632 9820
rect 5386 9766 5388 9818
rect 5568 9766 5570 9818
rect 5324 9764 5330 9766
rect 5386 9764 5410 9766
rect 5466 9764 5490 9766
rect 5546 9764 5570 9766
rect 5626 9764 5632 9766
rect 5324 9755 5632 9764
rect 5172 9580 5224 9586
rect 5092 9540 5172 9568
rect 5092 8974 5120 9540
rect 5172 9522 5224 9528
rect 5356 9580 5408 9586
rect 5540 9580 5592 9586
rect 5356 9522 5408 9528
rect 5460 9540 5540 9568
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5184 9178 5212 9386
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5368 9042 5396 9522
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5000 8838 5028 8910
rect 5368 8906 5396 8978
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4908 8622 5028 8650
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4080 8022 4108 8191
rect 4664 8188 4972 8197
rect 4664 8186 4670 8188
rect 4726 8186 4750 8188
rect 4806 8186 4830 8188
rect 4886 8186 4910 8188
rect 4966 8186 4972 8188
rect 4726 8134 4728 8186
rect 4908 8134 4910 8186
rect 4664 8132 4670 8134
rect 4726 8132 4750 8134
rect 4806 8132 4830 8134
rect 4886 8132 4910 8134
rect 4966 8132 4972 8134
rect 4664 8123 4972 8132
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 5000 7954 5028 8622
rect 5184 8344 5212 8842
rect 5460 8838 5488 9540
rect 5540 9522 5592 9528
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 9042 6224 9454
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5324 8732 5632 8741
rect 5324 8730 5330 8732
rect 5386 8730 5410 8732
rect 5466 8730 5490 8732
rect 5546 8730 5570 8732
rect 5626 8730 5632 8732
rect 5386 8678 5388 8730
rect 5568 8678 5570 8730
rect 5324 8676 5330 8678
rect 5386 8676 5410 8678
rect 5466 8676 5490 8678
rect 5546 8676 5570 8678
rect 5626 8676 5632 8678
rect 5324 8667 5632 8676
rect 5184 8316 5396 8344
rect 5368 7954 5396 8316
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 4068 7880 4120 7886
rect 3988 7828 4068 7834
rect 3988 7822 4120 7828
rect 3988 7806 4108 7822
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3804 7546 3832 7686
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3988 6934 4016 7806
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7478 4200 7686
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4080 5778 4108 7142
rect 4664 7100 4972 7109
rect 4664 7098 4670 7100
rect 4726 7098 4750 7100
rect 4806 7098 4830 7100
rect 4886 7098 4910 7100
rect 4966 7098 4972 7100
rect 4726 7046 4728 7098
rect 4908 7046 4910 7098
rect 4664 7044 4670 7046
rect 4726 7044 4750 7046
rect 4806 7044 4830 7046
rect 4886 7044 4910 7046
rect 4966 7044 4972 7046
rect 4664 7035 4972 7044
rect 5000 7002 5028 7890
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5184 7546 5212 7822
rect 5324 7644 5632 7653
rect 5324 7642 5330 7644
rect 5386 7642 5410 7644
rect 5466 7642 5490 7644
rect 5546 7642 5570 7644
rect 5626 7642 5632 7644
rect 5386 7590 5388 7642
rect 5568 7590 5570 7642
rect 5324 7588 5330 7590
rect 5386 7588 5410 7590
rect 5466 7588 5490 7590
rect 5546 7588 5570 7590
rect 5626 7588 5632 7590
rect 5324 7579 5632 7588
rect 5736 7546 5764 7890
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 6288 7342 6316 9998
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9654 6776 9862
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6380 7750 6408 8298
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7954 6960 8230
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 5324 6556 5632 6565
rect 5324 6554 5330 6556
rect 5386 6554 5410 6556
rect 5466 6554 5490 6556
rect 5546 6554 5570 6556
rect 5626 6554 5632 6556
rect 5386 6502 5388 6554
rect 5568 6502 5570 6554
rect 5324 6500 5330 6502
rect 5386 6500 5410 6502
rect 5466 6500 5490 6502
rect 5546 6500 5570 6502
rect 5626 6500 5632 6502
rect 5324 6491 5632 6500
rect 4664 6012 4972 6021
rect 4664 6010 4670 6012
rect 4726 6010 4750 6012
rect 4806 6010 4830 6012
rect 4886 6010 4910 6012
rect 4966 6010 4972 6012
rect 4726 5958 4728 6010
rect 4908 5958 4910 6010
rect 4664 5956 4670 5958
rect 4726 5956 4750 5958
rect 4806 5956 4830 5958
rect 4886 5956 4910 5958
rect 4966 5956 4972 5958
rect 4664 5947 4972 5956
rect 6104 5914 6132 6598
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 6748 5642 6776 6598
rect 7024 5778 7052 12718
rect 7392 11150 7420 13382
rect 8036 13326 8064 13790
rect 8312 13530 8340 16118
rect 8404 16114 8432 16458
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8496 15162 8524 15642
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 14074 8524 14214
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 12374 7512 12582
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7852 12306 7880 13126
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12442 8340 12786
rect 8588 12782 8616 16050
rect 8680 15722 8708 16186
rect 8864 16114 8892 17682
rect 8956 16436 8984 18226
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9324 17678 9352 18158
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9048 16590 9076 16934
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 8956 16408 9076 16436
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8680 15694 8800 15722
rect 8956 15706 8984 16050
rect 8668 13864 8720 13870
rect 8666 13832 8668 13841
rect 8720 13832 8722 13841
rect 8666 13767 8722 13776
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11150 7696 12106
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 7392 10810 7420 11086
rect 7668 10810 7696 11086
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 8312 10674 8340 11086
rect 8404 10810 8432 11086
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8392 10668 8444 10674
rect 8496 10656 8524 12242
rect 8680 12238 8708 13126
rect 8772 12986 8800 15694
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9048 15502 9076 16408
rect 9036 15496 9088 15502
rect 9140 15484 9168 16526
rect 9416 16250 9444 21490
rect 9508 21146 9536 21830
rect 9692 21672 9720 22578
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 22166 9904 22442
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9772 21684 9824 21690
rect 9692 21644 9772 21672
rect 9772 21626 9824 21632
rect 9876 21486 9904 21830
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9692 21146 9720 21286
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9876 21078 9904 21422
rect 9968 21146 9996 22578
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21350 10088 21966
rect 10612 21690 10640 24754
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10704 23866 10732 24074
rect 11072 24070 11100 24754
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12092 24508 12400 24517
rect 12092 24506 12098 24508
rect 12154 24506 12178 24508
rect 12234 24506 12258 24508
rect 12314 24506 12338 24508
rect 12394 24506 12400 24508
rect 12154 24454 12156 24506
rect 12336 24454 12338 24506
rect 12092 24452 12098 24454
rect 12154 24452 12178 24454
rect 12234 24452 12258 24454
rect 12314 24452 12338 24454
rect 12394 24452 12400 24454
rect 12092 24443 12400 24452
rect 12452 24342 12480 24550
rect 12440 24336 12492 24342
rect 12440 24278 12492 24284
rect 13096 24070 13124 24686
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10796 22778 10824 23734
rect 11072 23730 11100 24006
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11072 23322 11100 23666
rect 11152 23588 11204 23594
rect 11152 23530 11204 23536
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11164 23254 11192 23530
rect 11152 23248 11204 23254
rect 11152 23190 11204 23196
rect 11992 23118 12020 24006
rect 12752 23964 13060 23973
rect 12752 23962 12758 23964
rect 12814 23962 12838 23964
rect 12894 23962 12918 23964
rect 12974 23962 12998 23964
rect 13054 23962 13060 23964
rect 12814 23910 12816 23962
rect 12996 23910 12998 23962
rect 12752 23908 12758 23910
rect 12814 23908 12838 23910
rect 12894 23908 12918 23910
rect 12974 23908 12998 23910
rect 13054 23908 13060 23910
rect 12752 23899 13060 23908
rect 12092 23420 12400 23429
rect 12092 23418 12098 23420
rect 12154 23418 12178 23420
rect 12234 23418 12258 23420
rect 12314 23418 12338 23420
rect 12394 23418 12400 23420
rect 12154 23366 12156 23418
rect 12336 23366 12338 23418
rect 12092 23364 12098 23366
rect 12154 23364 12178 23366
rect 12234 23364 12258 23366
rect 12314 23364 12338 23366
rect 12394 23364 12400 23366
rect 12092 23355 12400 23364
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 11428 22704 11480 22710
rect 11428 22646 11480 22652
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10704 21554 10732 22374
rect 10980 22166 11008 22374
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9692 20806 9720 20946
rect 10060 20942 10088 21286
rect 10428 21162 10456 21490
rect 10336 21134 10456 21162
rect 10520 21146 10548 21490
rect 10796 21146 10824 21490
rect 10508 21140 10560 21146
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9600 20618 9628 20742
rect 9600 20590 9812 20618
rect 9876 20602 9904 20810
rect 9784 19922 9812 20590
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9508 18834 9536 19450
rect 9784 19310 9812 19858
rect 10152 19786 10180 20810
rect 10336 19922 10364 21134
rect 10508 21082 10560 21088
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10244 19514 10272 19790
rect 10428 19514 10456 21014
rect 10980 21010 11008 22102
rect 11072 22098 11100 22578
rect 11440 22386 11468 22646
rect 11256 22358 11468 22386
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 11256 21434 11284 22358
rect 11428 21956 11480 21962
rect 11624 21944 11652 22918
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11716 22234 11744 22578
rect 11808 22506 11836 22578
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11704 21956 11756 21962
rect 11624 21916 11704 21944
rect 11428 21898 11480 21904
rect 11704 21898 11756 21904
rect 11072 21418 11284 21434
rect 11060 21412 11284 21418
rect 11112 21406 11284 21412
rect 11060 21354 11112 21360
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11072 20874 11100 21354
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10980 20602 11008 20810
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 19990 11100 20266
rect 11164 20058 11192 20810
rect 11256 20398 11284 21406
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9508 16658 9536 18770
rect 9784 18154 9812 19246
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9876 18154 9904 18906
rect 11440 18426 11468 21898
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11532 20602 11560 20878
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11520 20596 11572 20602
rect 11520 20538 11572 20544
rect 11624 20466 11652 20810
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11612 19916 11664 19922
rect 11716 19904 11744 21898
rect 11808 20942 11836 22442
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11808 20602 11836 20878
rect 11900 20602 11928 22986
rect 11992 22778 12020 23054
rect 12268 22982 12296 23258
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12268 22778 12296 22918
rect 11980 22772 12032 22778
rect 11980 22714 12032 22720
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11992 21622 12020 22578
rect 12256 22500 12308 22506
rect 12360 22488 12388 22646
rect 12308 22460 12388 22488
rect 12256 22442 12308 22448
rect 12092 22332 12400 22341
rect 12092 22330 12098 22332
rect 12154 22330 12178 22332
rect 12234 22330 12258 22332
rect 12314 22330 12338 22332
rect 12394 22330 12400 22332
rect 12154 22278 12156 22330
rect 12336 22278 12338 22330
rect 12092 22276 12098 22278
rect 12154 22276 12178 22278
rect 12234 22276 12258 22278
rect 12314 22276 12338 22278
rect 12394 22276 12400 22278
rect 12092 22267 12400 22276
rect 11980 21616 12032 21622
rect 11980 21558 12032 21564
rect 11992 21146 12020 21558
rect 12092 21244 12400 21253
rect 12092 21242 12098 21244
rect 12154 21242 12178 21244
rect 12234 21242 12258 21244
rect 12314 21242 12338 21244
rect 12394 21242 12400 21244
rect 12154 21190 12156 21242
rect 12336 21190 12338 21242
rect 12092 21188 12098 21190
rect 12154 21188 12178 21190
rect 12234 21188 12258 21190
rect 12314 21188 12338 21190
rect 12394 21188 12400 21190
rect 12092 21179 12400 21188
rect 12452 21146 12480 23122
rect 12752 22876 13060 22885
rect 12752 22874 12758 22876
rect 12814 22874 12838 22876
rect 12894 22874 12918 22876
rect 12974 22874 12998 22876
rect 13054 22874 13060 22876
rect 12814 22822 12816 22874
rect 12996 22822 12998 22874
rect 12752 22820 12758 22822
rect 12814 22820 12838 22822
rect 12894 22820 12918 22822
rect 12974 22820 12998 22822
rect 13054 22820 13060 22822
rect 12752 22811 13060 22820
rect 12532 22500 12584 22506
rect 12532 22442 12584 22448
rect 12544 22030 12572 22442
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 13096 21962 13124 24006
rect 13268 23248 13320 23254
rect 13268 23190 13320 23196
rect 13176 22976 13228 22982
rect 13176 22918 13228 22924
rect 13188 22030 13216 22918
rect 13280 22642 13308 23190
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 13188 21894 13216 21966
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 11980 21140 12032 21146
rect 12440 21140 12492 21146
rect 11980 21082 12032 21088
rect 12360 21100 12440 21128
rect 12072 20800 12124 20806
rect 12072 20742 12124 20748
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 12084 20466 12112 20742
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12360 20262 12388 21100
rect 12440 21082 12492 21088
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 20602 12480 20810
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12092 20156 12400 20165
rect 12092 20154 12098 20156
rect 12154 20154 12178 20156
rect 12234 20154 12258 20156
rect 12314 20154 12338 20156
rect 12394 20154 12400 20156
rect 12154 20102 12156 20154
rect 12336 20102 12338 20154
rect 12092 20100 12098 20102
rect 12154 20100 12178 20102
rect 12234 20100 12258 20102
rect 12314 20100 12338 20102
rect 12394 20100 12400 20102
rect 12092 20091 12400 20100
rect 12452 19938 12480 20402
rect 12544 20058 12572 21830
rect 12752 21788 13060 21797
rect 12752 21786 12758 21788
rect 12814 21786 12838 21788
rect 12894 21786 12918 21788
rect 12974 21786 12998 21788
rect 13054 21786 13060 21788
rect 12814 21734 12816 21786
rect 12996 21734 12998 21786
rect 12752 21732 12758 21734
rect 12814 21732 12838 21734
rect 12894 21732 12918 21734
rect 12974 21732 12998 21734
rect 13054 21732 13060 21734
rect 12752 21723 13060 21732
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 21078 12664 21490
rect 13188 21350 13216 21830
rect 13280 21690 13308 22374
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 12624 21072 12676 21078
rect 12624 21014 12676 21020
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12752 20700 13060 20709
rect 12752 20698 12758 20700
rect 12814 20698 12838 20700
rect 12894 20698 12918 20700
rect 12974 20698 12998 20700
rect 13054 20698 13060 20700
rect 12814 20646 12816 20698
rect 12996 20646 12998 20698
rect 12752 20644 12758 20646
rect 12814 20644 12838 20646
rect 12894 20644 12918 20646
rect 12974 20644 12998 20646
rect 13054 20644 13060 20646
rect 12752 20635 13060 20644
rect 13096 20602 13124 20878
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12532 20052 12584 20058
rect 12584 20012 12664 20040
rect 12532 19994 12584 20000
rect 12452 19910 12572 19938
rect 11664 19876 11744 19904
rect 11612 19858 11664 19864
rect 11624 19718 11652 19858
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 12544 19378 12572 19910
rect 12636 19854 12664 20012
rect 12728 19854 12756 20198
rect 13372 20058 13400 29106
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14108 26042 14136 26318
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14384 25906 14412 26318
rect 14568 26042 14596 26930
rect 14648 26784 14700 26790
rect 14648 26726 14700 26732
rect 14844 26738 14872 31200
rect 15488 29306 15516 31200
rect 18156 29306 18184 31334
rect 20626 31200 20682 32000
rect 20180 29404 20488 29413
rect 20180 29402 20186 29404
rect 20242 29402 20266 29404
rect 20322 29402 20346 29404
rect 20402 29402 20426 29404
rect 20482 29402 20488 29404
rect 20242 29350 20244 29402
rect 20424 29350 20426 29402
rect 20180 29348 20186 29350
rect 20242 29348 20266 29350
rect 20322 29348 20346 29350
rect 20402 29348 20426 29350
rect 20482 29348 20488 29350
rect 20180 29339 20488 29348
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 16396 29164 16448 29170
rect 16396 29106 16448 29112
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 14556 26036 14608 26042
rect 14556 25978 14608 25984
rect 14660 25974 14688 26726
rect 14844 26710 15148 26738
rect 14740 26308 14792 26314
rect 14740 26250 14792 26256
rect 14752 26042 14780 26250
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14384 25498 14412 25842
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 14200 24206 14228 24618
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 14384 24274 14412 24550
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14200 23866 14228 24142
rect 14292 23866 14320 24142
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13556 23322 13584 23666
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13648 23254 13676 23666
rect 14384 23662 14412 24210
rect 14556 23724 14608 23730
rect 14740 23724 14792 23730
rect 14608 23684 14740 23712
rect 14556 23666 14608 23672
rect 14740 23666 14792 23672
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13636 23248 13688 23254
rect 13636 23190 13688 23196
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 21894 13584 22578
rect 13648 22234 13676 23190
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13740 21554 13768 23462
rect 14384 22642 14412 23598
rect 14832 23520 14884 23526
rect 14832 23462 14884 23468
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14844 22030 14872 23462
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 14936 22778 14964 22918
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 20602 13768 20742
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13832 20466 13860 21830
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14016 20262 14044 21966
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14464 21344 14516 21350
rect 14568 21321 14596 21830
rect 14844 21554 14872 21966
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14464 21286 14516 21292
rect 14554 21312 14610 21321
rect 14292 20874 14320 21286
rect 14280 20868 14332 20874
rect 14280 20810 14332 20816
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12752 19612 13060 19621
rect 12752 19610 12758 19612
rect 12814 19610 12838 19612
rect 12894 19610 12918 19612
rect 12974 19610 12998 19612
rect 13054 19610 13060 19612
rect 12814 19558 12816 19610
rect 12996 19558 12998 19610
rect 12752 19556 12758 19558
rect 12814 19556 12838 19558
rect 12894 19556 12918 19558
rect 12974 19556 12998 19558
rect 13054 19556 13060 19558
rect 12752 19547 13060 19556
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 13648 19242 13676 20198
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13924 19378 13952 19926
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 12092 19068 12400 19077
rect 12092 19066 12098 19068
rect 12154 19066 12178 19068
rect 12234 19066 12258 19068
rect 12314 19066 12338 19068
rect 12394 19066 12400 19068
rect 12154 19014 12156 19066
rect 12336 19014 12338 19066
rect 12092 19012 12098 19014
rect 12154 19012 12178 19014
rect 12234 19012 12258 19014
rect 12314 19012 12338 19014
rect 12394 19012 12400 19014
rect 12092 19003 12400 19012
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 11716 18306 11744 18566
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 12072 18352 12124 18358
rect 11716 18300 12072 18306
rect 11716 18294 12124 18300
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11716 18278 12112 18294
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17338 9628 18022
rect 9784 17678 9812 18090
rect 9876 17882 9904 18090
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 10060 17746 10088 18158
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10152 17678 10180 18090
rect 10612 18034 10640 18090
rect 10520 18006 10640 18034
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10520 17882 10548 18006
rect 11072 17882 11100 18022
rect 11440 17882 11468 18226
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16794 9720 17138
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9600 16658 9628 16730
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15706 9444 15982
rect 9404 15700 9456 15706
rect 9456 15660 9628 15688
rect 9404 15642 9456 15648
rect 9220 15496 9272 15502
rect 9140 15456 9220 15484
rect 9036 15438 9088 15444
rect 9220 15438 9272 15444
rect 9128 14068 9180 14074
rect 9404 14068 9456 14074
rect 9180 14028 9404 14056
rect 9128 14010 9180 14016
rect 9404 14010 9456 14016
rect 9600 13954 9628 15660
rect 9692 15094 9720 16730
rect 9784 15502 9812 17614
rect 10520 16794 10548 17818
rect 11072 17610 11100 17818
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 11072 16114 11100 17138
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9968 14958 9996 15302
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9784 14618 9812 14894
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9692 14414 9720 14554
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9416 13938 9720 13954
rect 9416 13932 9732 13938
rect 9416 13926 9680 13932
rect 9220 13864 9272 13870
rect 9416 13852 9444 13926
rect 9680 13874 9732 13880
rect 9272 13824 9444 13852
rect 9588 13864 9640 13870
rect 9220 13806 9272 13812
rect 9588 13806 9640 13812
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8864 12918 8892 13466
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8864 12434 8892 12854
rect 9416 12850 9444 13398
rect 9508 12866 9536 13670
rect 9600 13462 9628 13806
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9588 12912 9640 12918
rect 9508 12860 9588 12866
rect 9508 12854 9640 12860
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9508 12838 9628 12854
rect 9692 12850 9720 13874
rect 9968 13802 9996 14350
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 10152 13326 10180 13942
rect 10244 13326 10272 15098
rect 10888 15042 10916 15506
rect 11072 15162 11100 16050
rect 11164 15570 11192 16594
rect 11256 15706 11284 16934
rect 11716 16046 11744 18278
rect 12636 18222 12664 19178
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 12752 18524 13060 18533
rect 12752 18522 12758 18524
rect 12814 18522 12838 18524
rect 12894 18522 12918 18524
rect 12974 18522 12998 18524
rect 13054 18522 13060 18524
rect 12814 18470 12816 18522
rect 12996 18470 12998 18522
rect 12752 18468 12758 18470
rect 12814 18468 12838 18470
rect 12894 18468 12918 18470
rect 12974 18468 12998 18470
rect 13054 18468 13060 18470
rect 12752 18459 13060 18468
rect 13372 18426 13400 19110
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17542 11928 18022
rect 12092 17980 12400 17989
rect 12092 17978 12098 17980
rect 12154 17978 12178 17980
rect 12234 17978 12258 17980
rect 12314 17978 12338 17980
rect 12394 17978 12400 17980
rect 12154 17926 12156 17978
rect 12336 17926 12338 17978
rect 12092 17924 12098 17926
rect 12154 17924 12178 17926
rect 12234 17924 12258 17926
rect 12314 17924 12338 17926
rect 12394 17924 12400 17926
rect 12092 17915 12400 17924
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 16794 11928 17478
rect 12084 17202 12112 17614
rect 12360 17202 12388 17750
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12636 17338 12664 17546
rect 12752 17436 13060 17445
rect 12752 17434 12758 17436
rect 12814 17434 12838 17436
rect 12894 17434 12918 17436
rect 12974 17434 12998 17436
rect 13054 17434 13060 17436
rect 12814 17382 12816 17434
rect 12996 17382 12998 17434
rect 12752 17380 12758 17382
rect 12814 17380 12838 17382
rect 12894 17380 12918 17382
rect 12974 17380 12998 17382
rect 13054 17380 13060 17382
rect 12752 17371 13060 17380
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 13464 17202 13492 18158
rect 12072 17196 12124 17202
rect 12348 17196 12400 17202
rect 12072 17138 12124 17144
rect 12268 17156 12348 17184
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10888 15014 11008 15042
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9680 12844 9732 12850
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8772 12406 8892 12434
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8444 10628 8524 10656
rect 8392 10610 8444 10616
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10266 7972 10406
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8588 10010 8616 10950
rect 8312 9982 8616 10010
rect 8312 9042 8340 9982
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 9586 8616 9862
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8588 9450 8616 9522
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8498 7604 8774
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7208 8090 7236 8434
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7208 7818 7236 8026
rect 7392 7886 7420 8230
rect 7576 8090 7604 8434
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7546 7236 7754
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6254 7512 6598
rect 7668 6254 7696 8842
rect 8312 8634 8340 8978
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8772 8566 8800 12406
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 10470 8892 10610
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 8560 8812 8566
rect 8680 8508 8760 8514
rect 8680 8502 8812 8508
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8680 8486 8800 8502
rect 8128 8022 8156 8434
rect 8220 8090 8248 8434
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8680 7478 8708 8486
rect 8956 8378 8984 12718
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 12442 9260 12582
rect 9324 12442 9352 12786
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9416 11558 9444 12582
rect 9508 12238 9536 12838
rect 9680 12786 9732 12792
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9784 12730 9812 12922
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9600 12238 9628 12718
rect 9784 12702 9904 12730
rect 9772 12640 9824 12646
rect 9692 12600 9772 12628
rect 9692 12442 9720 12600
rect 9772 12582 9824 12588
rect 9680 12436 9732 12442
rect 9876 12434 9904 12702
rect 10060 12442 10088 12786
rect 9680 12378 9732 12384
rect 9784 12406 9904 12434
rect 10048 12436 10100 12442
rect 9784 12238 9812 12406
rect 10048 12378 10100 12384
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9600 11354 9628 12174
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11898 9720 12038
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 10060 11626 10088 12378
rect 10152 11830 10180 13262
rect 10520 12782 10548 14350
rect 10888 14006 10916 14894
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10782 13832 10838 13841
rect 10782 13767 10838 13776
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10612 12850 10640 13262
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10796 11898 10824 13767
rect 10980 13682 11008 15014
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11164 14618 11192 14962
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11256 14346 11284 15302
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10980 13654 11100 13682
rect 11072 12481 11100 13654
rect 11058 12472 11114 12481
rect 11058 12407 11114 12416
rect 11164 11914 11192 14010
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11256 12714 11284 13126
rect 11348 12986 11376 15438
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11440 12986 11468 13194
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 11072 11886 11192 11914
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9140 10674 9168 11222
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9048 9994 9076 10542
rect 9232 10062 9260 10678
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10062 9352 10610
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 9232 9518 9260 9998
rect 9324 9722 9352 9998
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9692 9586 9720 11494
rect 10152 11354 10180 11494
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9876 10266 9904 11154
rect 10796 11150 10824 11834
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10060 10606 10088 11086
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9968 10266 9996 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9876 10146 9904 10202
rect 10060 10146 10088 10406
rect 9876 10118 10088 10146
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10612 9586 10640 9862
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9324 8974 9352 9522
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9178 9536 9386
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9312 8968 9364 8974
rect 9232 8928 9312 8956
rect 9232 8498 9260 8928
rect 9312 8910 9364 8916
rect 9508 8566 9536 9114
rect 9692 8974 9720 9522
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8566 9720 8910
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9312 8424 9364 8430
rect 8760 8356 8812 8362
rect 8956 8350 9076 8378
rect 9312 8366 9364 8372
rect 8760 8298 8812 8304
rect 8772 8022 8800 8298
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8760 8016 8812 8022
rect 8864 7993 8892 8026
rect 8760 7958 8812 7964
rect 8850 7984 8906 7993
rect 8850 7919 8906 7928
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8956 7206 8984 8230
rect 9048 7410 9076 8350
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9140 7818 9168 8230
rect 9232 7954 9260 8230
rect 9324 7954 9352 8366
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 8090 9444 8230
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8312 6866 8340 7142
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 7484 5914 7512 6190
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 5324 5468 5632 5477
rect 5324 5466 5330 5468
rect 5386 5466 5410 5468
rect 5466 5466 5490 5468
rect 5546 5466 5570 5468
rect 5626 5466 5632 5468
rect 5386 5414 5388 5466
rect 5568 5414 5570 5466
rect 5324 5412 5330 5414
rect 5386 5412 5410 5414
rect 5466 5412 5490 5414
rect 5546 5412 5570 5414
rect 5626 5412 5632 5414
rect 5324 5403 5632 5412
rect 4664 4924 4972 4933
rect 4664 4922 4670 4924
rect 4726 4922 4750 4924
rect 4806 4922 4830 4924
rect 4886 4922 4910 4924
rect 4966 4922 4972 4924
rect 4726 4870 4728 4922
rect 4908 4870 4910 4922
rect 4664 4868 4670 4870
rect 4726 4868 4750 4870
rect 4806 4868 4830 4870
rect 4886 4868 4910 4870
rect 4966 4868 4972 4870
rect 4664 4859 4972 4868
rect 5324 4380 5632 4389
rect 5324 4378 5330 4380
rect 5386 4378 5410 4380
rect 5466 4378 5490 4380
rect 5546 4378 5570 4380
rect 5626 4378 5632 4380
rect 5386 4326 5388 4378
rect 5568 4326 5570 4378
rect 5324 4324 5330 4326
rect 5386 4324 5410 4326
rect 5466 4324 5490 4326
rect 5546 4324 5570 4326
rect 5626 4324 5632 4326
rect 5324 4315 5632 4324
rect 4664 3836 4972 3845
rect 4664 3834 4670 3836
rect 4726 3834 4750 3836
rect 4806 3834 4830 3836
rect 4886 3834 4910 3836
rect 4966 3834 4972 3836
rect 4726 3782 4728 3834
rect 4908 3782 4910 3834
rect 4664 3780 4670 3782
rect 4726 3780 4750 3782
rect 4806 3780 4830 3782
rect 4886 3780 4910 3782
rect 4966 3780 4972 3782
rect 4664 3771 4972 3780
rect 5324 3292 5632 3301
rect 5324 3290 5330 3292
rect 5386 3290 5410 3292
rect 5466 3290 5490 3292
rect 5546 3290 5570 3292
rect 5626 3290 5632 3292
rect 5386 3238 5388 3290
rect 5568 3238 5570 3290
rect 5324 3236 5330 3238
rect 5386 3236 5410 3238
rect 5466 3236 5490 3238
rect 5546 3236 5570 3238
rect 5626 3236 5632 3238
rect 5324 3227 5632 3236
rect 4664 2748 4972 2757
rect 4664 2746 4670 2748
rect 4726 2746 4750 2748
rect 4806 2746 4830 2748
rect 4886 2746 4910 2748
rect 4966 2746 4972 2748
rect 4726 2694 4728 2746
rect 4908 2694 4910 2746
rect 4664 2692 4670 2694
rect 4726 2692 4750 2694
rect 4806 2692 4830 2694
rect 4886 2692 4910 2694
rect 4966 2692 4972 2694
rect 4664 2683 4972 2692
rect 5324 2204 5632 2213
rect 5324 2202 5330 2204
rect 5386 2202 5410 2204
rect 5466 2202 5490 2204
rect 5546 2202 5570 2204
rect 5626 2202 5632 2204
rect 5386 2150 5388 2202
rect 5568 2150 5570 2202
rect 5324 2148 5330 2150
rect 5386 2148 5410 2150
rect 5466 2148 5490 2150
rect 5546 2148 5570 2150
rect 5626 2148 5632 2150
rect 5324 2139 5632 2148
rect 8404 800 8432 6190
rect 9140 6186 9168 6938
rect 9324 6798 9352 7890
rect 9508 7886 9536 8502
rect 10520 8498 10548 8774
rect 10796 8634 10824 9522
rect 11072 9500 11100 11886
rect 11256 11762 11284 12650
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11164 11354 11192 11698
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11532 9586 11560 14418
rect 11624 14006 11652 15370
rect 11808 14890 11836 16662
rect 11992 16522 12020 17070
rect 12268 16998 12296 17156
rect 12348 17138 12400 17144
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12092 16892 12400 16901
rect 12092 16890 12098 16892
rect 12154 16890 12178 16892
rect 12234 16890 12258 16892
rect 12314 16890 12338 16892
rect 12394 16890 12400 16892
rect 12154 16838 12156 16890
rect 12336 16838 12338 16890
rect 12092 16836 12098 16838
rect 12154 16836 12178 16838
rect 12234 16836 12258 16838
rect 12314 16836 12338 16838
rect 12394 16836 12400 16838
rect 12092 16827 12400 16836
rect 12636 16658 12664 17138
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16658 13308 16934
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15586 11928 16390
rect 11992 15706 12020 16458
rect 13464 16454 13492 17138
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 12752 16348 13060 16357
rect 12752 16346 12758 16348
rect 12814 16346 12838 16348
rect 12894 16346 12918 16348
rect 12974 16346 12998 16348
rect 13054 16346 13060 16348
rect 12814 16294 12816 16346
rect 12996 16294 12998 16346
rect 12752 16292 12758 16294
rect 12814 16292 12838 16294
rect 12894 16292 12918 16294
rect 12974 16292 12998 16294
rect 13054 16292 13060 16294
rect 12752 16283 13060 16292
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12092 15804 12400 15813
rect 12092 15802 12098 15804
rect 12154 15802 12178 15804
rect 12234 15802 12258 15804
rect 12314 15802 12338 15804
rect 12394 15802 12400 15804
rect 12154 15750 12156 15802
rect 12336 15750 12338 15802
rect 12092 15748 12098 15750
rect 12154 15748 12178 15750
rect 12234 15748 12258 15750
rect 12314 15748 12338 15750
rect 12394 15748 12400 15750
rect 12092 15739 12400 15748
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11900 15558 12112 15586
rect 12084 15094 12112 15558
rect 13096 15502 13124 15846
rect 13280 15502 13308 16050
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13084 15496 13136 15502
rect 12530 15464 12586 15473
rect 13268 15496 13320 15502
rect 13084 15438 13136 15444
rect 13188 15456 13268 15484
rect 12530 15399 12586 15408
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11900 14618 11928 14962
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11992 14498 12020 14826
rect 12092 14716 12400 14725
rect 12092 14714 12098 14716
rect 12154 14714 12178 14716
rect 12234 14714 12258 14716
rect 12314 14714 12338 14716
rect 12394 14714 12400 14716
rect 12154 14662 12156 14714
rect 12336 14662 12338 14714
rect 12092 14660 12098 14662
rect 12154 14660 12178 14662
rect 12234 14660 12258 14662
rect 12314 14660 12338 14662
rect 12394 14660 12400 14662
rect 12092 14651 12400 14660
rect 11808 14074 11836 14486
rect 11992 14482 12112 14498
rect 11992 14476 12124 14482
rect 11992 14470 12072 14476
rect 12072 14418 12124 14424
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11624 12646 11652 13942
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11610 12472 11666 12481
rect 11610 12407 11666 12416
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11244 9512 11296 9518
rect 11072 9472 11244 9500
rect 11244 9454 11296 9460
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 9586 7984 9642 7993
rect 9586 7919 9642 7928
rect 9600 7886 9628 7919
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 9416 7546 9444 7686
rect 10060 7546 10088 7686
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10520 7002 10548 7686
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10612 6882 10640 8298
rect 10888 8090 10916 8366
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10704 7954 10732 8026
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10520 6854 10640 6882
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9324 6458 9352 6734
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9140 5710 9168 6122
rect 9324 5914 9352 6394
rect 9508 6118 9536 6598
rect 10520 6322 10548 6854
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6458 10640 6734
rect 10704 6662 10732 7890
rect 10980 7886 11008 8434
rect 11256 8362 11284 9454
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11348 8498 11376 8978
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 7410 10824 7686
rect 11624 7410 11652 12407
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 11164 6322 11192 7346
rect 11716 6866 11744 13942
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12918 11928 13330
rect 11888 12912 11940 12918
rect 11808 12860 11888 12866
rect 11808 12854 11940 12860
rect 11808 12838 11928 12854
rect 11808 11082 11836 12838
rect 11992 12764 12020 13806
rect 12092 13628 12400 13637
rect 12092 13626 12098 13628
rect 12154 13626 12178 13628
rect 12234 13626 12258 13628
rect 12314 13626 12338 13628
rect 12394 13626 12400 13628
rect 12154 13574 12156 13626
rect 12336 13574 12338 13626
rect 12092 13572 12098 13574
rect 12154 13572 12178 13574
rect 12234 13572 12258 13574
rect 12314 13572 12338 13574
rect 12394 13572 12400 13574
rect 12092 13563 12400 13572
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 12176 12918 12204 13194
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11900 12736 12020 12764
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 9466 11836 11018
rect 11900 9586 11928 12736
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 9586 12020 12582
rect 12092 12540 12400 12549
rect 12092 12538 12098 12540
rect 12154 12538 12178 12540
rect 12234 12538 12258 12540
rect 12314 12538 12338 12540
rect 12394 12538 12400 12540
rect 12154 12486 12156 12538
rect 12336 12486 12338 12538
rect 12092 12484 12098 12486
rect 12154 12484 12178 12486
rect 12234 12484 12258 12486
rect 12314 12484 12338 12486
rect 12394 12484 12400 12486
rect 12092 12475 12400 12484
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12092 11452 12400 11461
rect 12092 11450 12098 11452
rect 12154 11450 12178 11452
rect 12234 11450 12258 11452
rect 12314 11450 12338 11452
rect 12394 11450 12400 11452
rect 12154 11398 12156 11450
rect 12336 11398 12338 11450
rect 12092 11396 12098 11398
rect 12154 11396 12178 11398
rect 12234 11396 12258 11398
rect 12314 11396 12338 11398
rect 12394 11396 12400 11398
rect 12092 11387 12400 11396
rect 12452 11354 12480 11766
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12092 10364 12400 10373
rect 12092 10362 12098 10364
rect 12154 10362 12178 10364
rect 12234 10362 12258 10364
rect 12314 10362 12338 10364
rect 12394 10362 12400 10364
rect 12154 10310 12156 10362
rect 12336 10310 12338 10362
rect 12092 10308 12098 10310
rect 12154 10308 12178 10310
rect 12234 10308 12258 10310
rect 12314 10308 12338 10310
rect 12394 10308 12400 10310
rect 12092 10299 12400 10308
rect 12544 10010 12572 15399
rect 12752 15260 13060 15269
rect 12752 15258 12758 15260
rect 12814 15258 12838 15260
rect 12894 15258 12918 15260
rect 12974 15258 12998 15260
rect 13054 15258 13060 15260
rect 12814 15206 12816 15258
rect 12996 15206 12998 15258
rect 12752 15204 12758 15206
rect 12814 15204 12838 15206
rect 12894 15204 12918 15206
rect 12974 15204 12998 15206
rect 13054 15204 13060 15206
rect 12752 15195 13060 15204
rect 12752 14172 13060 14181
rect 12752 14170 12758 14172
rect 12814 14170 12838 14172
rect 12894 14170 12918 14172
rect 12974 14170 12998 14172
rect 13054 14170 13060 14172
rect 12814 14118 12816 14170
rect 12996 14118 12998 14170
rect 12752 14116 12758 14118
rect 12814 14116 12838 14118
rect 12894 14116 12918 14118
rect 12974 14116 12998 14118
rect 13054 14116 13060 14118
rect 12752 14107 13060 14116
rect 13096 13938 13124 15438
rect 13188 14414 13216 15456
rect 13268 15438 13320 15444
rect 13372 14958 13400 15574
rect 13464 15502 13492 16390
rect 13556 16182 13584 17070
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13556 15570 13584 15982
rect 13648 15706 13676 19178
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18970 13860 19110
rect 13924 18970 13952 19314
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 14016 18290 14044 20198
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14004 18284 14056 18290
rect 13924 18244 14004 18272
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13740 16046 13768 17206
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16794 13860 17070
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13924 16114 13952 18244
rect 14004 18226 14056 18232
rect 14108 18086 14136 19178
rect 14200 18290 14228 20742
rect 14292 20398 14320 20810
rect 14476 20534 14504 21286
rect 14554 21247 14610 21256
rect 14568 20942 14596 21247
rect 15028 21146 15056 21422
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14464 20528 14516 20534
rect 14464 20470 14516 20476
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18426 14320 18702
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14004 16992 14056 16998
rect 14108 16980 14136 18022
rect 14056 16952 14136 16980
rect 14004 16934 14056 16940
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13740 15586 13768 15642
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13648 15558 13768 15586
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13556 15026 13584 15506
rect 13648 15094 13676 15558
rect 13728 15496 13780 15502
rect 13726 15464 13728 15473
rect 13820 15496 13872 15502
rect 13780 15464 13782 15473
rect 13820 15438 13872 15444
rect 13726 15399 13782 15408
rect 13832 15162 13860 15438
rect 14108 15366 14136 16952
rect 14200 15910 14228 18226
rect 14476 18222 14504 19382
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14844 18290 14872 19178
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14568 16794 14596 17206
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12752 13084 13060 13093
rect 12752 13082 12758 13084
rect 12814 13082 12838 13084
rect 12894 13082 12918 13084
rect 12974 13082 12998 13084
rect 13054 13082 13060 13084
rect 12814 13030 12816 13082
rect 12996 13030 12998 13082
rect 12752 13028 12758 13030
rect 12814 13028 12838 13030
rect 12894 13028 12918 13030
rect 12974 13028 12998 13030
rect 13054 13028 13060 13030
rect 12752 13019 13060 13028
rect 13096 12986 13124 13126
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12752 11996 13060 12005
rect 12752 11994 12758 11996
rect 12814 11994 12838 11996
rect 12894 11994 12918 11996
rect 12974 11994 12998 11996
rect 13054 11994 13060 11996
rect 12814 11942 12816 11994
rect 12996 11942 12998 11994
rect 12752 11940 12758 11942
rect 12814 11940 12838 11942
rect 12894 11940 12918 11942
rect 12974 11940 12998 11942
rect 13054 11940 13060 11942
rect 12752 11931 13060 11940
rect 12752 10908 13060 10917
rect 12752 10906 12758 10908
rect 12814 10906 12838 10908
rect 12894 10906 12918 10908
rect 12974 10906 12998 10908
rect 13054 10906 13060 10908
rect 12814 10854 12816 10906
rect 12996 10854 12998 10906
rect 12752 10852 12758 10854
rect 12814 10852 12838 10854
rect 12894 10852 12918 10854
rect 12974 10852 12998 10854
rect 13054 10852 13060 10854
rect 12752 10843 13060 10852
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12360 9982 12572 10010
rect 12360 9654 12388 9982
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 11808 9438 11928 9466
rect 11900 8906 11928 9438
rect 12092 9276 12400 9285
rect 12092 9274 12098 9276
rect 12154 9274 12178 9276
rect 12234 9274 12258 9276
rect 12314 9274 12338 9276
rect 12394 9274 12400 9276
rect 12154 9222 12156 9274
rect 12336 9222 12338 9274
rect 12092 9220 12098 9222
rect 12154 9220 12178 9222
rect 12234 9220 12258 9222
rect 12314 9220 12338 9222
rect 12394 9220 12400 9222
rect 12092 9211 12400 9220
rect 12452 9110 12480 9522
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 6458 11284 6666
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6458 11560 6598
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5914 9536 6054
rect 11256 5914 11284 6122
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11532 5778 11560 6054
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11532 5370 11560 5578
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11900 5234 11928 8842
rect 12544 8838 12572 9862
rect 12636 9722 12664 10610
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 10266 13216 10406
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12752 9820 13060 9829
rect 12752 9818 12758 9820
rect 12814 9818 12838 9820
rect 12894 9818 12918 9820
rect 12974 9818 12998 9820
rect 13054 9818 13060 9820
rect 12814 9766 12816 9818
rect 12996 9766 12998 9818
rect 12752 9764 12758 9766
rect 12814 9764 12838 9766
rect 12894 9764 12918 9766
rect 12974 9764 12998 9766
rect 13054 9764 13060 9766
rect 12752 9755 13060 9764
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 9178 12664 9318
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12728 9058 12756 9386
rect 13096 9110 13124 9998
rect 13280 9722 13308 14214
rect 13464 13852 13492 14894
rect 13556 14414 13584 14962
rect 13832 14822 13860 15098
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14906 14044 14962
rect 13924 14878 14044 14906
rect 14292 14890 14320 16526
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14384 15570 14412 16118
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14280 14884 14332 14890
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13544 13864 13596 13870
rect 13464 13824 13544 13852
rect 13544 13806 13596 13812
rect 13556 12306 13584 13806
rect 13648 13394 13676 14758
rect 13924 13938 13952 14878
rect 14280 14826 14332 14832
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10810 13400 11494
rect 13464 11218 13492 11698
rect 13556 11558 13584 12242
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11286 13584 11494
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 11082 13492 11154
rect 13648 11150 13676 13330
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13832 10674 13860 10950
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13556 10266 13584 10610
rect 13924 10538 13952 12922
rect 14108 12646 14136 13806
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14200 12442 14228 14350
rect 14660 14278 14688 15302
rect 14752 15026 14780 17614
rect 14844 17338 14872 18226
rect 15028 18154 15056 20742
rect 15120 19310 15148 26710
rect 15212 26246 15240 26930
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15200 26240 15252 26246
rect 15200 26182 15252 26188
rect 15212 25294 15240 26182
rect 15396 25906 15424 26726
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15488 25498 15516 26930
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15580 25294 15608 26182
rect 16224 26042 16252 26318
rect 16212 26036 16264 26042
rect 16212 25978 16264 25984
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15488 24274 15516 24754
rect 16408 24274 16436 29106
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 17144 26586 17172 26726
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16776 25906 16804 26318
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16960 25974 16988 26182
rect 16948 25968 17000 25974
rect 16948 25910 17000 25916
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16776 24818 16804 25842
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 17972 24886 18000 25094
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 15488 23730 15516 24210
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 15580 23866 15608 24074
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 16316 23798 16344 24006
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 16028 23656 16080 23662
rect 16028 23598 16080 23604
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15212 22030 15240 22510
rect 15672 22234 15700 23054
rect 16040 23050 16068 23598
rect 16028 23044 16080 23050
rect 16028 22986 16080 22992
rect 15752 22976 15804 22982
rect 15752 22918 15804 22924
rect 15764 22710 15792 22918
rect 15752 22704 15804 22710
rect 15752 22646 15804 22652
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21486 15240 21966
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 21690 15332 21898
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15120 18766 15148 19246
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 15212 16794 15240 20266
rect 15304 16794 15332 20878
rect 15580 20466 15608 20946
rect 15672 20602 15700 20946
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15948 20602 15976 20810
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16046 14872 16390
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 15028 15706 15056 16526
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15396 14822 15424 18702
rect 15672 17746 15700 20538
rect 16040 20534 16068 22986
rect 16408 21146 16436 24210
rect 16776 24206 16804 24754
rect 18064 24410 18092 29106
rect 19520 28860 19828 28869
rect 19520 28858 19526 28860
rect 19582 28858 19606 28860
rect 19662 28858 19686 28860
rect 19742 28858 19766 28860
rect 19822 28858 19828 28860
rect 19582 28806 19584 28858
rect 19764 28806 19766 28858
rect 19520 28804 19526 28806
rect 19582 28804 19606 28806
rect 19662 28804 19686 28806
rect 19742 28804 19766 28806
rect 19822 28804 19828 28806
rect 19520 28795 19828 28804
rect 20180 28316 20488 28325
rect 20180 28314 20186 28316
rect 20242 28314 20266 28316
rect 20322 28314 20346 28316
rect 20402 28314 20426 28316
rect 20482 28314 20488 28316
rect 20242 28262 20244 28314
rect 20424 28262 20426 28314
rect 20180 28260 20186 28262
rect 20242 28260 20266 28262
rect 20322 28260 20346 28262
rect 20402 28260 20426 28262
rect 20482 28260 20488 28262
rect 20180 28251 20488 28260
rect 19520 27772 19828 27781
rect 19520 27770 19526 27772
rect 19582 27770 19606 27772
rect 19662 27770 19686 27772
rect 19742 27770 19766 27772
rect 19822 27770 19828 27772
rect 19582 27718 19584 27770
rect 19764 27718 19766 27770
rect 19520 27716 19526 27718
rect 19582 27716 19606 27718
rect 19662 27716 19686 27718
rect 19742 27716 19766 27718
rect 19822 27716 19828 27718
rect 19520 27707 19828 27716
rect 20640 27690 20668 31200
rect 27608 29404 27916 29413
rect 27608 29402 27614 29404
rect 27670 29402 27694 29404
rect 27750 29402 27774 29404
rect 27830 29402 27854 29404
rect 27910 29402 27916 29404
rect 27670 29350 27672 29402
rect 27852 29350 27854 29402
rect 27608 29348 27614 29350
rect 27670 29348 27694 29350
rect 27750 29348 27774 29350
rect 27830 29348 27854 29350
rect 27910 29348 27916 29350
rect 27608 29339 27916 29348
rect 26948 28860 27256 28869
rect 26948 28858 26954 28860
rect 27010 28858 27034 28860
rect 27090 28858 27114 28860
rect 27170 28858 27194 28860
rect 27250 28858 27256 28860
rect 27010 28806 27012 28858
rect 27192 28806 27194 28858
rect 26948 28804 26954 28806
rect 27010 28804 27034 28806
rect 27090 28804 27114 28806
rect 27170 28804 27194 28806
rect 27250 28804 27256 28806
rect 26948 28795 27256 28804
rect 27608 28316 27916 28325
rect 27608 28314 27614 28316
rect 27670 28314 27694 28316
rect 27750 28314 27774 28316
rect 27830 28314 27854 28316
rect 27910 28314 27916 28316
rect 27670 28262 27672 28314
rect 27852 28262 27854 28314
rect 27608 28260 27614 28262
rect 27670 28260 27694 28262
rect 27750 28260 27774 28262
rect 27830 28260 27854 28262
rect 27910 28260 27916 28262
rect 27608 28251 27916 28260
rect 26948 27772 27256 27781
rect 26948 27770 26954 27772
rect 27010 27770 27034 27772
rect 27090 27770 27114 27772
rect 27170 27770 27194 27772
rect 27250 27770 27256 27772
rect 27010 27718 27012 27770
rect 27192 27718 27194 27770
rect 26948 27716 26954 27718
rect 27010 27716 27034 27718
rect 27090 27716 27114 27718
rect 27170 27716 27194 27718
rect 27250 27716 27256 27718
rect 26948 27707 27256 27716
rect 20640 27662 20760 27690
rect 20180 27228 20488 27237
rect 20180 27226 20186 27228
rect 20242 27226 20266 27228
rect 20322 27226 20346 27228
rect 20402 27226 20426 27228
rect 20482 27226 20488 27228
rect 20242 27174 20244 27226
rect 20424 27174 20426 27226
rect 20180 27172 20186 27174
rect 20242 27172 20266 27174
rect 20322 27172 20346 27174
rect 20402 27172 20426 27174
rect 20482 27172 20488 27174
rect 20180 27163 20488 27172
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18708 26042 18736 26862
rect 19892 26852 19944 26858
rect 19892 26794 19944 26800
rect 19520 26684 19828 26693
rect 19520 26682 19526 26684
rect 19582 26682 19606 26684
rect 19662 26682 19686 26684
rect 19742 26682 19766 26684
rect 19822 26682 19828 26684
rect 19582 26630 19584 26682
rect 19764 26630 19766 26682
rect 19520 26628 19526 26630
rect 19582 26628 19606 26630
rect 19662 26628 19686 26630
rect 19742 26628 19766 26630
rect 19822 26628 19828 26630
rect 19520 26619 19828 26628
rect 19904 26586 19932 26794
rect 19892 26580 19944 26586
rect 19892 26522 19944 26528
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 19904 25702 19932 26522
rect 20180 26140 20488 26149
rect 20180 26138 20186 26140
rect 20242 26138 20266 26140
rect 20322 26138 20346 26140
rect 20402 26138 20426 26140
rect 20482 26138 20488 26140
rect 20242 26086 20244 26138
rect 20424 26086 20426 26138
rect 20180 26084 20186 26086
rect 20242 26084 20266 26086
rect 20322 26084 20346 26086
rect 20402 26084 20426 26086
rect 20482 26084 20488 26086
rect 20180 26075 20488 26084
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 18524 25498 18552 25638
rect 19520 25596 19828 25605
rect 19520 25594 19526 25596
rect 19582 25594 19606 25596
rect 19662 25594 19686 25596
rect 19742 25594 19766 25596
rect 19822 25594 19828 25596
rect 19582 25542 19584 25594
rect 19764 25542 19766 25594
rect 19520 25540 19526 25542
rect 19582 25540 19606 25542
rect 19662 25540 19686 25542
rect 19742 25540 19766 25542
rect 19822 25540 19828 25542
rect 19520 25531 19828 25540
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16776 22438 16804 24142
rect 18156 24138 18184 24550
rect 18524 24410 18552 24618
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18800 24342 18828 25094
rect 20180 25052 20488 25061
rect 20180 25050 20186 25052
rect 20242 25050 20266 25052
rect 20322 25050 20346 25052
rect 20402 25050 20426 25052
rect 20482 25050 20488 25052
rect 20242 24998 20244 25050
rect 20424 24998 20426 25050
rect 20180 24996 20186 24998
rect 20242 24996 20266 24998
rect 20322 24996 20346 24998
rect 20402 24996 20426 24998
rect 20482 24996 20488 24998
rect 20180 24987 20488 24996
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 18788 24336 18840 24342
rect 18788 24278 18840 24284
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23866 16896 24006
rect 18892 23866 18920 24550
rect 19076 24410 19104 24754
rect 19520 24508 19828 24517
rect 19520 24506 19526 24508
rect 19582 24506 19606 24508
rect 19662 24506 19686 24508
rect 19742 24506 19766 24508
rect 19822 24506 19828 24508
rect 19582 24454 19584 24506
rect 19764 24454 19766 24506
rect 19520 24452 19526 24454
rect 19582 24452 19606 24454
rect 19662 24452 19686 24454
rect 19742 24452 19766 24454
rect 19822 24452 19828 24454
rect 19520 24443 19828 24452
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19248 24200 19300 24206
rect 19300 24148 19380 24154
rect 19248 24142 19380 24148
rect 19260 24126 19380 24142
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 19248 23520 19300 23526
rect 19352 23474 19380 24126
rect 20180 23964 20488 23973
rect 20180 23962 20186 23964
rect 20242 23962 20266 23964
rect 20322 23962 20346 23964
rect 20402 23962 20426 23964
rect 20482 23962 20488 23964
rect 20242 23910 20244 23962
rect 20424 23910 20426 23962
rect 20180 23908 20186 23910
rect 20242 23908 20266 23910
rect 20322 23908 20346 23910
rect 20402 23908 20426 23910
rect 20482 23908 20488 23910
rect 20180 23899 20488 23908
rect 19300 23468 19380 23474
rect 19248 23462 19380 23468
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 19260 23446 19380 23462
rect 19352 23186 19380 23446
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19444 22794 19472 23462
rect 19520 23420 19828 23429
rect 19520 23418 19526 23420
rect 19582 23418 19606 23420
rect 19662 23418 19686 23420
rect 19742 23418 19766 23420
rect 19822 23418 19828 23420
rect 19582 23366 19584 23418
rect 19764 23366 19766 23418
rect 19520 23364 19526 23366
rect 19582 23364 19606 23366
rect 19662 23364 19686 23366
rect 19742 23364 19766 23366
rect 19822 23364 19828 23366
rect 19520 23355 19828 23364
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 19352 22766 19472 22794
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16776 22094 16804 22374
rect 16960 22234 16988 22510
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 17880 22166 17908 22714
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 16684 22066 16804 22094
rect 17776 22092 17828 22098
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16592 20874 16620 21286
rect 16684 21010 16712 22066
rect 17776 22034 17828 22040
rect 16764 21956 16816 21962
rect 16764 21898 16816 21904
rect 16776 21622 16804 21898
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 21690 17724 21830
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 16764 21616 16816 21622
rect 16816 21576 16896 21604
rect 16764 21558 16816 21564
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16776 20466 16804 20742
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16040 19514 16068 19654
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16224 19378 16252 19790
rect 16776 19514 16804 20402
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16224 18766 16252 19314
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16776 18970 16804 19246
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16868 18630 16896 21576
rect 17788 20398 17816 22034
rect 17972 22030 18000 22374
rect 18064 22234 18092 22578
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 18696 22092 18748 22098
rect 18984 22094 19012 22374
rect 18696 22034 18748 22040
rect 18800 22066 19288 22094
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18512 21956 18564 21962
rect 18512 21898 18564 21904
rect 18524 21690 18552 21898
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21690 18644 21830
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15580 16658 15608 17138
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15856 16590 15884 17138
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16114 15884 16526
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15366 15700 15846
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14568 13326 14596 14010
rect 14660 13870 14688 14214
rect 15672 13870 15700 14758
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12918 14596 13262
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 15212 12850 15240 13330
rect 15304 13326 15332 13670
rect 15292 13320 15344 13326
rect 15344 13280 15424 13308
rect 15292 13262 15344 13268
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 14188 12436 14240 12442
rect 15212 12434 15240 12786
rect 15396 12434 15424 13280
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15212 12406 15332 12434
rect 15396 12406 15516 12434
rect 14188 12378 14240 12384
rect 14200 11830 14228 12378
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11898 15240 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 11354 14964 11494
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 14844 10062 14872 10950
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10062 14964 10542
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13372 9586 13400 9998
rect 14200 9586 14228 9998
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 9178 13216 9318
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12636 9030 12756 9058
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8634 12572 8774
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12092 8188 12400 8197
rect 12092 8186 12098 8188
rect 12154 8186 12178 8188
rect 12234 8186 12258 8188
rect 12314 8186 12338 8188
rect 12394 8186 12400 8188
rect 12154 8134 12156 8186
rect 12336 8134 12338 8186
rect 12092 8132 12098 8134
rect 12154 8132 12178 8134
rect 12234 8132 12258 8134
rect 12314 8132 12338 8134
rect 12394 8132 12400 8134
rect 12092 8123 12400 8132
rect 12452 8090 12480 8434
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12636 7954 12664 9030
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12728 8838 12756 8910
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12752 8732 13060 8741
rect 12752 8730 12758 8732
rect 12814 8730 12838 8732
rect 12894 8730 12918 8732
rect 12974 8730 12998 8732
rect 13054 8730 13060 8732
rect 12814 8678 12816 8730
rect 12996 8678 12998 8730
rect 12752 8676 12758 8678
rect 12814 8676 12838 8678
rect 12894 8676 12918 8678
rect 12974 8676 12998 8678
rect 13054 8676 13060 8678
rect 12752 8667 13060 8676
rect 13372 8514 13400 9522
rect 14200 8974 14228 9522
rect 14936 9178 14964 9998
rect 15028 9586 15056 11154
rect 15304 10810 15332 12406
rect 15488 12238 15516 12406
rect 15580 12306 15608 12582
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 10810 15424 12038
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15120 10606 15148 10746
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10062 15148 10542
rect 15396 10266 15424 10746
rect 15488 10674 15516 11290
rect 15856 11286 15884 15506
rect 15948 15473 15976 18158
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17746 16620 18022
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16868 17338 16896 18566
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16868 16182 16896 17274
rect 16856 16176 16908 16182
rect 16856 16118 16908 16124
rect 15934 15464 15990 15473
rect 15934 15399 15990 15408
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15948 15026 15976 15302
rect 16316 15162 16344 15370
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 16960 14770 16988 19314
rect 17052 18766 17080 19858
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 17236 19242 17264 19722
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17236 18834 17264 19178
rect 17328 18970 17356 19994
rect 17420 19514 17448 20266
rect 17880 20244 17908 21558
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17788 20216 17908 20244
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17328 18766 17356 18906
rect 17512 18766 17540 19790
rect 17696 19378 17724 19926
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17788 19310 17816 20216
rect 17868 20052 17920 20058
rect 17972 20040 18000 20742
rect 17920 20012 18000 20040
rect 17868 19994 17920 20000
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17604 18970 17632 19246
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 17052 17338 17080 17546
rect 17236 17338 17264 18226
rect 17604 18222 17632 18702
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17776 18148 17828 18154
rect 17776 18090 17828 18096
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17224 17332 17276 17338
rect 17224 17274 17276 17280
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16182 17080 16934
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17788 16114 17816 18090
rect 17880 17338 17908 19314
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17972 17814 18000 18022
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17972 17338 18000 17750
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15434 17080 15846
rect 17788 15620 17816 16050
rect 17868 15632 17920 15638
rect 17788 15592 17868 15620
rect 17868 15574 17920 15580
rect 17972 15502 18000 16662
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 18064 15162 18092 21422
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18156 19174 18184 19314
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18902 18184 19110
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18156 16182 18184 16458
rect 18248 16250 18276 21490
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18340 21321 18368 21354
rect 18604 21344 18656 21350
rect 18326 21312 18382 21321
rect 18604 21286 18656 21292
rect 18326 21247 18382 21256
rect 18616 19854 18644 21286
rect 18708 21078 18736 22034
rect 18800 21554 18828 22066
rect 19260 22030 19288 22066
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19076 21690 19104 21966
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 18708 20330 18736 21014
rect 18800 20942 18828 21490
rect 19352 21418 19380 22766
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19352 21026 19380 21354
rect 19444 21146 19472 22374
rect 19520 22332 19828 22341
rect 19520 22330 19526 22332
rect 19582 22330 19606 22332
rect 19662 22330 19686 22332
rect 19742 22330 19766 22332
rect 19822 22330 19828 22332
rect 19582 22278 19584 22330
rect 19764 22278 19766 22330
rect 19520 22276 19526 22278
rect 19582 22276 19606 22278
rect 19662 22276 19686 22278
rect 19742 22276 19766 22278
rect 19822 22276 19828 22278
rect 19520 22267 19828 22276
rect 19904 22094 19932 22374
rect 19628 22066 19932 22094
rect 19628 22030 19656 22066
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19812 21894 19840 21966
rect 19800 21888 19852 21894
rect 19800 21830 19852 21836
rect 19904 21554 19932 22066
rect 19996 21690 20024 23122
rect 20548 23050 20576 23462
rect 20640 23186 20668 25230
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20180 22876 20488 22885
rect 20180 22874 20186 22876
rect 20242 22874 20266 22876
rect 20322 22874 20346 22876
rect 20402 22874 20426 22876
rect 20482 22874 20488 22876
rect 20242 22822 20244 22874
rect 20424 22822 20426 22874
rect 20180 22820 20186 22822
rect 20242 22820 20266 22822
rect 20322 22820 20346 22822
rect 20402 22820 20426 22822
rect 20482 22820 20488 22822
rect 20180 22811 20488 22820
rect 20168 22500 20220 22506
rect 20168 22442 20220 22448
rect 20180 22030 20208 22442
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20168 22024 20220 22030
rect 20088 21984 20168 22012
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20088 21604 20116 21984
rect 20168 21966 20220 21972
rect 20180 21788 20488 21797
rect 20180 21786 20186 21788
rect 20242 21786 20266 21788
rect 20322 21786 20346 21788
rect 20402 21786 20426 21788
rect 20482 21786 20488 21788
rect 20242 21734 20244 21786
rect 20424 21734 20426 21786
rect 20180 21732 20186 21734
rect 20242 21732 20266 21734
rect 20322 21732 20346 21734
rect 20402 21732 20426 21734
rect 20482 21732 20488 21734
rect 20180 21723 20488 21732
rect 20168 21616 20220 21622
rect 20088 21576 20168 21604
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19520 21244 19828 21253
rect 19520 21242 19526 21244
rect 19582 21242 19606 21244
rect 19662 21242 19686 21244
rect 19742 21242 19766 21244
rect 19822 21242 19828 21244
rect 19582 21190 19584 21242
rect 19764 21190 19766 21242
rect 19520 21188 19526 21190
rect 19582 21188 19606 21190
rect 19662 21188 19686 21190
rect 19742 21188 19766 21190
rect 19822 21188 19828 21190
rect 19520 21179 19828 21188
rect 19432 21140 19484 21146
rect 19484 21100 19656 21128
rect 19432 21082 19484 21088
rect 19352 20998 19564 21026
rect 19628 21010 19656 21100
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 18800 20398 18828 20878
rect 18892 20466 18920 20878
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18984 20466 19012 20810
rect 19352 20534 19380 20878
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 19536 20482 19564 20998
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 20088 20890 20116 21576
rect 20168 21558 20220 21564
rect 20352 21548 20404 21554
rect 20548 21536 20576 22102
rect 20404 21508 20576 21536
rect 20352 21490 20404 21496
rect 20364 21146 20392 21490
rect 20444 21344 20496 21350
rect 20628 21344 20680 21350
rect 20496 21292 20628 21298
rect 20444 21286 20680 21292
rect 20456 21270 20668 21286
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20732 21010 20760 27662
rect 27608 27228 27916 27237
rect 27608 27226 27614 27228
rect 27670 27226 27694 27228
rect 27750 27226 27774 27228
rect 27830 27226 27854 27228
rect 27910 27226 27916 27228
rect 27670 27174 27672 27226
rect 27852 27174 27854 27226
rect 27608 27172 27614 27174
rect 27670 27172 27694 27174
rect 27750 27172 27774 27174
rect 27830 27172 27854 27174
rect 27910 27172 27916 27174
rect 27608 27163 27916 27172
rect 26948 26684 27256 26693
rect 26948 26682 26954 26684
rect 27010 26682 27034 26684
rect 27090 26682 27114 26684
rect 27170 26682 27194 26684
rect 27250 26682 27256 26684
rect 27010 26630 27012 26682
rect 27192 26630 27194 26682
rect 26948 26628 26954 26630
rect 27010 26628 27034 26630
rect 27090 26628 27114 26630
rect 27170 26628 27194 26630
rect 27250 26628 27256 26630
rect 26948 26619 27256 26628
rect 27608 26140 27916 26149
rect 27608 26138 27614 26140
rect 27670 26138 27694 26140
rect 27750 26138 27774 26140
rect 27830 26138 27854 26140
rect 27910 26138 27916 26140
rect 27670 26086 27672 26138
rect 27852 26086 27854 26138
rect 27608 26084 27614 26086
rect 27670 26084 27694 26086
rect 27750 26084 27774 26086
rect 27830 26084 27854 26086
rect 27910 26084 27916 26086
rect 27608 26075 27916 26084
rect 26948 25596 27256 25605
rect 26948 25594 26954 25596
rect 27010 25594 27034 25596
rect 27090 25594 27114 25596
rect 27170 25594 27194 25596
rect 27250 25594 27256 25596
rect 27010 25542 27012 25594
rect 27192 25542 27194 25594
rect 26948 25540 26954 25542
rect 27010 25540 27034 25542
rect 27090 25540 27114 25542
rect 27170 25540 27194 25542
rect 27250 25540 27256 25542
rect 26948 25531 27256 25540
rect 27608 25052 27916 25061
rect 27608 25050 27614 25052
rect 27670 25050 27694 25052
rect 27750 25050 27774 25052
rect 27830 25050 27854 25052
rect 27910 25050 27916 25052
rect 27670 24998 27672 25050
rect 27852 24998 27854 25050
rect 27608 24996 27614 24998
rect 27670 24996 27694 24998
rect 27750 24996 27774 24998
rect 27830 24996 27854 24998
rect 27910 24996 27916 24998
rect 27608 24987 27916 24996
rect 26948 24508 27256 24517
rect 26948 24506 26954 24508
rect 27010 24506 27034 24508
rect 27090 24506 27114 24508
rect 27170 24506 27194 24508
rect 27250 24506 27256 24508
rect 27010 24454 27012 24506
rect 27192 24454 27194 24506
rect 26948 24452 26954 24454
rect 27010 24452 27034 24454
rect 27090 24452 27114 24454
rect 27170 24452 27194 24454
rect 27250 24452 27256 24454
rect 26948 24443 27256 24452
rect 27608 23964 27916 23973
rect 27608 23962 27614 23964
rect 27670 23962 27694 23964
rect 27750 23962 27774 23964
rect 27830 23962 27854 23964
rect 27910 23962 27916 23964
rect 27670 23910 27672 23962
rect 27852 23910 27854 23962
rect 27608 23908 27614 23910
rect 27670 23908 27694 23910
rect 27750 23908 27774 23910
rect 27830 23908 27854 23910
rect 27910 23908 27916 23910
rect 27608 23899 27916 23908
rect 25412 23792 25464 23798
rect 25412 23734 25464 23740
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20824 22778 20852 23666
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24400 23588 24452 23594
rect 24400 23530 24452 23536
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23492 23050 23520 23462
rect 23940 23180 23992 23186
rect 23940 23122 23992 23128
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21928 22778 21956 22918
rect 22756 22778 22784 22986
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21192 22234 21220 22510
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21928 22166 21956 22714
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21916 22160 21968 22166
rect 21916 22102 21968 22108
rect 21822 21992 21878 22001
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 21548 21956 21600 21962
rect 21822 21927 21824 21936
rect 21548 21898 21600 21904
rect 21876 21927 21878 21936
rect 21824 21898 21876 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20824 21486 20852 21830
rect 21192 21690 21220 21898
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21560 21554 21588 21898
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20824 21010 20852 21422
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 19996 20862 20116 20890
rect 19892 20800 19944 20806
rect 19996 20788 20024 20862
rect 19944 20760 20024 20788
rect 19892 20742 19944 20748
rect 19996 20602 20024 20760
rect 20076 20800 20128 20806
rect 20076 20742 20128 20748
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 19352 20058 19380 20470
rect 19536 20454 20024 20482
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19444 19938 19472 20198
rect 19520 20156 19828 20165
rect 19520 20154 19526 20156
rect 19582 20154 19606 20156
rect 19662 20154 19686 20156
rect 19742 20154 19766 20156
rect 19822 20154 19828 20156
rect 19582 20102 19584 20154
rect 19764 20102 19766 20154
rect 19520 20100 19526 20102
rect 19582 20100 19606 20102
rect 19662 20100 19686 20102
rect 19742 20100 19766 20102
rect 19822 20100 19828 20102
rect 19520 20091 19828 20100
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19352 19910 19472 19938
rect 18604 19848 18656 19854
rect 18656 19808 18828 19836
rect 18604 19790 18656 19796
rect 18696 19712 18748 19718
rect 18340 19638 18552 19666
rect 18696 19654 18748 19660
rect 18340 18970 18368 19638
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18340 17066 18368 17138
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18156 15706 18184 16118
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17224 14816 17276 14822
rect 16960 14742 17172 14770
rect 17224 14758 17276 14764
rect 16960 14618 16988 14742
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16132 13938 16160 14350
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15580 10538 15608 10950
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15856 10452 15884 11222
rect 15936 10464 15988 10470
rect 15856 10424 15936 10452
rect 15936 10406 15988 10412
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14200 8634 14228 8910
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 13280 8486 13400 8514
rect 14384 8498 14412 8910
rect 13636 8492 13688 8498
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11992 7410 12020 7754
rect 12752 7644 13060 7653
rect 12752 7642 12758 7644
rect 12814 7642 12838 7644
rect 12894 7642 12918 7644
rect 12974 7642 12998 7644
rect 13054 7642 13060 7644
rect 12814 7590 12816 7642
rect 12996 7590 12998 7642
rect 12752 7588 12758 7590
rect 12814 7588 12838 7590
rect 12894 7588 12918 7590
rect 12974 7588 12998 7590
rect 13054 7588 13060 7590
rect 12752 7579 13060 7588
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 8390 0 8446 800
rect 11992 762 12020 7346
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12092 7100 12400 7109
rect 12092 7098 12098 7100
rect 12154 7098 12178 7100
rect 12234 7098 12258 7100
rect 12314 7098 12338 7100
rect 12394 7098 12400 7100
rect 12154 7046 12156 7098
rect 12336 7046 12338 7098
rect 12092 7044 12098 7046
rect 12154 7044 12178 7046
rect 12234 7044 12258 7046
rect 12314 7044 12338 7046
rect 12394 7044 12400 7046
rect 12092 7035 12400 7044
rect 12728 7002 12756 7142
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12820 6730 12848 7142
rect 12912 6798 12940 7142
rect 13096 7002 13124 7346
rect 13188 7206 13216 7346
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13280 7002 13308 8486
rect 13636 8434 13688 8440
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13268 6996 13320 7002
rect 13268 6938 13320 6944
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 12752 6556 13060 6565
rect 12752 6554 12758 6556
rect 12814 6554 12838 6556
rect 12894 6554 12918 6556
rect 12974 6554 12998 6556
rect 13054 6554 13060 6556
rect 12814 6502 12816 6554
rect 12996 6502 12998 6554
rect 12752 6500 12758 6502
rect 12814 6500 12838 6502
rect 12894 6500 12918 6502
rect 12974 6500 12998 6502
rect 13054 6500 13060 6502
rect 12752 6491 13060 6500
rect 12092 6012 12400 6021
rect 12092 6010 12098 6012
rect 12154 6010 12178 6012
rect 12234 6010 12258 6012
rect 12314 6010 12338 6012
rect 12394 6010 12400 6012
rect 12154 5958 12156 6010
rect 12336 5958 12338 6010
rect 12092 5956 12098 5958
rect 12154 5956 12178 5958
rect 12234 5956 12258 5958
rect 12314 5956 12338 5958
rect 12394 5956 12400 5958
rect 12092 5947 12400 5956
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12268 5234 12296 5510
rect 12544 5370 12572 5646
rect 13280 5642 13308 6666
rect 13372 5914 13400 7346
rect 13464 6662 13492 7822
rect 13648 6730 13676 8434
rect 14568 8430 14596 9114
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15212 8634 15240 8910
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 8294 14596 8366
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 7336 13780 7342
rect 13832 7290 13860 7686
rect 14568 7410 14596 8230
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 13780 7284 13860 7290
rect 13728 7278 13860 7284
rect 13740 7262 13860 7278
rect 13832 7002 13860 7262
rect 13924 7290 13952 7346
rect 15304 7342 15332 8026
rect 15396 7818 15424 8774
rect 15488 8566 15516 9046
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15856 8430 15884 9522
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 8498 16068 9454
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15292 7336 15344 7342
rect 13924 7274 14136 7290
rect 15292 7278 15344 7284
rect 13924 7268 14148 7274
rect 13924 7262 14096 7268
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6934 13952 7262
rect 14096 7210 14148 7216
rect 14464 7200 14516 7206
rect 15292 7200 15344 7206
rect 14516 7148 14872 7154
rect 14464 7142 14872 7148
rect 15292 7142 15344 7148
rect 14476 7126 14872 7142
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 14844 6798 14872 7126
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14936 6798 14964 6938
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13464 5846 13492 6598
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 12752 5468 13060 5477
rect 12752 5466 12758 5468
rect 12814 5466 12838 5468
rect 12894 5466 12918 5468
rect 12974 5466 12998 5468
rect 13054 5466 13060 5468
rect 12814 5414 12816 5466
rect 12996 5414 12998 5466
rect 12752 5412 12758 5414
rect 12814 5412 12838 5414
rect 12894 5412 12918 5414
rect 12974 5412 12998 5414
rect 13054 5412 13060 5414
rect 12752 5403 13060 5412
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 13280 5166 13308 5578
rect 13464 5574 13492 5782
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 5302 13492 5510
rect 13648 5370 13676 6666
rect 13740 6458 13768 6734
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 14292 5914 14320 6734
rect 14844 6254 14872 6734
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14108 5370 14136 5646
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13452 5296 13504 5302
rect 13452 5238 13504 5244
rect 14752 5166 14780 5510
rect 14844 5234 14872 5510
rect 15212 5370 15240 6802
rect 15304 6798 15332 7142
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15396 6458 15424 6734
rect 15488 6730 15516 7346
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15580 6322 15608 7210
rect 15672 6322 15700 7346
rect 15856 6866 15884 8366
rect 15948 7546 15976 8434
rect 16040 8090 16068 8434
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 16040 6458 16068 7890
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5778 15332 6190
rect 16040 5778 16068 6394
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 12092 4924 12400 4933
rect 12092 4922 12098 4924
rect 12154 4922 12178 4924
rect 12234 4922 12258 4924
rect 12314 4922 12338 4924
rect 12394 4922 12400 4924
rect 12154 4870 12156 4922
rect 12336 4870 12338 4922
rect 12092 4868 12098 4870
rect 12154 4868 12178 4870
rect 12234 4868 12258 4870
rect 12314 4868 12338 4870
rect 12394 4868 12400 4870
rect 12092 4859 12400 4868
rect 12752 4380 13060 4389
rect 12752 4378 12758 4380
rect 12814 4378 12838 4380
rect 12894 4378 12918 4380
rect 12974 4378 12998 4380
rect 13054 4378 13060 4380
rect 12814 4326 12816 4378
rect 12996 4326 12998 4378
rect 12752 4324 12758 4326
rect 12814 4324 12838 4326
rect 12894 4324 12918 4326
rect 12974 4324 12998 4326
rect 13054 4324 13060 4326
rect 12752 4315 13060 4324
rect 16132 4146 16160 13874
rect 16224 13394 16252 14214
rect 16592 13530 16620 14282
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 13870 16896 14214
rect 16856 13864 16908 13870
rect 16776 13824 16856 13852
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16224 12646 16252 13330
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16684 12986 16712 13262
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12238 16252 12582
rect 16776 12434 16804 13824
rect 16856 13806 16908 13812
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12986 16896 13126
rect 16960 12986 16988 13194
rect 17052 12986 17080 13262
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12782 17172 14742
rect 17236 14618 17264 14758
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17696 14074 17724 14282
rect 17788 14074 17816 14350
rect 17684 14068 17736 14074
rect 17684 14010 17736 14016
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17788 13394 17816 14010
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17144 12434 17172 12718
rect 16684 12406 16804 12434
rect 16960 12406 17172 12434
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10606 16528 11018
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16500 9994 16528 10542
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9654 16620 9862
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16408 8498 16436 9386
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16408 7002 16436 8434
rect 16592 8294 16620 8774
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16592 7546 16620 8230
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6322 16436 6598
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16316 5778 16344 6054
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 12092 3836 12400 3845
rect 12092 3834 12098 3836
rect 12154 3834 12178 3836
rect 12234 3834 12258 3836
rect 12314 3834 12338 3836
rect 12394 3834 12400 3836
rect 12154 3782 12156 3834
rect 12336 3782 12338 3834
rect 12092 3780 12098 3782
rect 12154 3780 12178 3782
rect 12234 3780 12258 3782
rect 12314 3780 12338 3782
rect 12394 3780 12400 3782
rect 12092 3771 12400 3780
rect 12752 3292 13060 3301
rect 12752 3290 12758 3292
rect 12814 3290 12838 3292
rect 12894 3290 12918 3292
rect 12974 3290 12998 3292
rect 13054 3290 13060 3292
rect 12814 3238 12816 3290
rect 12996 3238 12998 3290
rect 12752 3236 12758 3238
rect 12814 3236 12838 3238
rect 12894 3236 12918 3238
rect 12974 3236 12998 3238
rect 13054 3236 13060 3238
rect 12752 3227 13060 3236
rect 12092 2748 12400 2757
rect 12092 2746 12098 2748
rect 12154 2746 12178 2748
rect 12234 2746 12258 2748
rect 12314 2746 12338 2748
rect 12394 2746 12400 2748
rect 12154 2694 12156 2746
rect 12336 2694 12338 2746
rect 12092 2692 12098 2694
rect 12154 2692 12178 2694
rect 12234 2692 12258 2694
rect 12314 2692 12338 2694
rect 12394 2692 12400 2694
rect 12092 2683 12400 2692
rect 12752 2204 13060 2213
rect 12752 2202 12758 2204
rect 12814 2202 12838 2204
rect 12894 2202 12918 2204
rect 12974 2202 12998 2204
rect 13054 2202 13060 2204
rect 12814 2150 12816 2202
rect 12996 2150 12998 2202
rect 12752 2148 12758 2150
rect 12814 2148 12838 2150
rect 12894 2148 12918 2150
rect 12974 2148 12998 2150
rect 13054 2148 13060 2150
rect 12752 2139 13060 2148
rect 12176 870 12296 898
rect 12176 762 12204 870
rect 12268 800 12296 870
rect 14844 800 14872 4082
rect 16684 2774 16712 12406
rect 16960 11830 16988 12406
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16960 11082 16988 11290
rect 17144 11150 17172 12242
rect 17236 11694 17264 12718
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17420 12434 17448 12650
rect 17420 12406 17540 12434
rect 17512 12238 17540 12406
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11762 17356 12038
rect 17696 11762 17724 12922
rect 17788 12434 17816 13330
rect 17880 13326 17908 14350
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 18064 12434 18092 15098
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 13326 18184 14214
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 18248 12918 18276 16186
rect 18340 16046 18368 17002
rect 18432 16794 18460 19450
rect 18524 19360 18552 19638
rect 18708 19514 18736 19654
rect 18800 19514 18828 19808
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18892 19378 18920 19654
rect 19168 19378 19196 19858
rect 19352 19378 19380 19910
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 19514 19472 19790
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 18604 19372 18656 19378
rect 18524 19332 18604 19360
rect 18604 19314 18656 19320
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 18892 19258 18920 19314
rect 18892 19230 19012 19258
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18426 18920 19110
rect 18984 18902 19012 19230
rect 19076 18970 19104 19314
rect 19168 18970 19196 19314
rect 19520 19068 19828 19077
rect 19520 19066 19526 19068
rect 19582 19066 19606 19068
rect 19662 19066 19686 19068
rect 19742 19066 19766 19068
rect 19822 19066 19828 19068
rect 19582 19014 19584 19066
rect 19764 19014 19766 19066
rect 19520 19012 19526 19014
rect 19582 19012 19606 19014
rect 19662 19012 19686 19014
rect 19742 19012 19766 19014
rect 19822 19012 19828 19014
rect 19520 19003 19828 19012
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18984 18766 19012 18838
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18892 16946 18920 18362
rect 18984 17882 19012 18702
rect 19260 18086 19288 18770
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19156 17876 19208 17882
rect 19156 17818 19208 17824
rect 18892 16918 19012 16946
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18432 15162 18460 15642
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18524 14958 18552 16458
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18616 16046 18644 16186
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15638 18644 15846
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18708 15502 18736 16118
rect 18800 16046 18828 16526
rect 18892 16522 18920 16730
rect 18880 16516 18932 16522
rect 18880 16458 18932 16464
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18800 15026 18828 15982
rect 18892 15706 18920 16458
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18328 13252 18380 13258
rect 18380 13212 18460 13240
rect 18328 13194 18380 13200
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 17788 12406 17908 12434
rect 18064 12406 18184 12434
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16960 10674 16988 11018
rect 17144 10810 17172 11086
rect 17420 11082 17448 11698
rect 17788 11558 17816 12038
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 11218 17816 11494
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17880 11150 17908 12406
rect 17868 11144 17920 11150
rect 17920 11104 18000 11132
rect 17868 11086 17920 11092
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9722 16804 9862
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16868 9586 16896 10066
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16960 9518 16988 10610
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17144 9586 17172 10474
rect 17328 10266 17356 10610
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9674 17356 10066
rect 17236 9646 17356 9674
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 8906 16804 9318
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 16776 8566 16804 8842
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 7886 16804 8230
rect 17144 8090 17172 8366
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17236 7954 17264 9646
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 8362 17356 9522
rect 17420 9518 17448 11018
rect 17972 10674 18000 11104
rect 17960 10668 18012 10674
rect 18012 10628 18092 10656
rect 17960 10610 18012 10616
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 9994 17540 10406
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17972 8090 18000 8502
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18064 7954 18092 10628
rect 18156 9586 18184 12406
rect 18432 11558 18460 13212
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18248 9926 18276 11494
rect 18340 11082 18368 11494
rect 18432 11150 18460 11494
rect 18524 11150 18552 13330
rect 18708 12850 18736 14758
rect 18800 14550 18828 14962
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18984 14414 19012 16918
rect 19168 16726 19196 17818
rect 19260 17678 19288 18022
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 17338 19380 17478
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19352 15094 19380 16186
rect 19444 15978 19472 18022
rect 19520 17980 19828 17989
rect 19520 17978 19526 17980
rect 19582 17978 19606 17980
rect 19662 17978 19686 17980
rect 19742 17978 19766 17980
rect 19822 17978 19828 17980
rect 19582 17926 19584 17978
rect 19764 17926 19766 17978
rect 19520 17924 19526 17926
rect 19582 17924 19606 17926
rect 19662 17924 19686 17926
rect 19742 17924 19766 17926
rect 19822 17924 19828 17926
rect 19520 17915 19828 17924
rect 19904 17882 19932 18702
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19904 17270 19932 17478
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19520 16892 19828 16901
rect 19520 16890 19526 16892
rect 19582 16890 19606 16892
rect 19662 16890 19686 16892
rect 19742 16890 19766 16892
rect 19822 16890 19828 16892
rect 19582 16838 19584 16890
rect 19764 16838 19766 16890
rect 19520 16836 19526 16838
rect 19582 16836 19606 16838
rect 19662 16836 19686 16838
rect 19742 16836 19766 16838
rect 19822 16836 19828 16838
rect 19520 16827 19828 16836
rect 19904 16794 19932 16934
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19996 16658 20024 20454
rect 20088 20058 20116 20742
rect 20180 20700 20488 20709
rect 20180 20698 20186 20700
rect 20242 20698 20266 20700
rect 20322 20698 20346 20700
rect 20402 20698 20426 20700
rect 20482 20698 20488 20700
rect 20242 20646 20244 20698
rect 20424 20646 20426 20698
rect 20180 20644 20186 20646
rect 20242 20644 20266 20646
rect 20322 20644 20346 20646
rect 20402 20644 20426 20646
rect 20482 20644 20488 20646
rect 20180 20635 20488 20644
rect 20732 20602 20760 20946
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 21008 19922 21036 20810
rect 21836 20754 21864 21898
rect 21928 20874 21956 22102
rect 22112 22030 22140 22374
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21836 20726 22048 20754
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20088 19514 20116 19790
rect 20180 19612 20488 19621
rect 20180 19610 20186 19612
rect 20242 19610 20266 19612
rect 20322 19610 20346 19612
rect 20402 19610 20426 19612
rect 20482 19610 20488 19612
rect 20242 19558 20244 19610
rect 20424 19558 20426 19610
rect 20180 19556 20186 19558
rect 20242 19556 20266 19558
rect 20322 19556 20346 19558
rect 20402 19556 20426 19558
rect 20482 19556 20488 19558
rect 20180 19547 20488 19556
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20088 18222 20116 19450
rect 20548 19446 20576 19790
rect 20536 19440 20588 19446
rect 20536 19382 20588 19388
rect 20732 19310 20760 19790
rect 20824 19378 20852 19790
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20824 19258 20852 19314
rect 20824 19230 21036 19258
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20916 18698 20944 19110
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20180 18524 20488 18533
rect 20180 18522 20186 18524
rect 20242 18522 20266 18524
rect 20322 18522 20346 18524
rect 20402 18522 20426 18524
rect 20482 18522 20488 18524
rect 20242 18470 20244 18522
rect 20424 18470 20426 18522
rect 20180 18468 20186 18470
rect 20242 18468 20266 18470
rect 20322 18468 20346 18470
rect 20402 18468 20426 18470
rect 20482 18468 20488 18470
rect 20180 18459 20488 18468
rect 20916 18290 20944 18634
rect 21008 18290 21036 19230
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20088 17202 20116 18158
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 20180 17542 20208 17750
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20180 17436 20488 17445
rect 20180 17434 20186 17436
rect 20242 17434 20266 17436
rect 20322 17434 20346 17436
rect 20402 17434 20426 17436
rect 20482 17434 20488 17436
rect 20242 17382 20244 17434
rect 20424 17382 20426 17434
rect 20180 17380 20186 17382
rect 20242 17380 20266 17382
rect 20322 17380 20346 17382
rect 20402 17380 20426 17382
rect 20482 17380 20488 17382
rect 20180 17371 20488 17380
rect 20548 17202 20576 18226
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20536 16788 20588 16794
rect 20536 16730 20588 16736
rect 20076 16720 20128 16726
rect 20076 16662 20128 16668
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19260 14906 19288 14962
rect 19064 14884 19116 14890
rect 19260 14878 19380 14906
rect 19064 14826 19116 14832
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18892 13938 18920 14282
rect 19076 14074 19104 14826
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19168 13938 19196 14282
rect 19260 14278 19288 14418
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 13938 19288 14214
rect 19352 13954 19380 14878
rect 19444 14396 19472 15914
rect 19520 15804 19828 15813
rect 19520 15802 19526 15804
rect 19582 15802 19606 15804
rect 19662 15802 19686 15804
rect 19742 15802 19766 15804
rect 19822 15802 19828 15804
rect 19582 15750 19584 15802
rect 19764 15750 19766 15802
rect 19520 15748 19526 15750
rect 19582 15748 19606 15750
rect 19662 15748 19686 15750
rect 19742 15748 19766 15750
rect 19822 15748 19828 15750
rect 19520 15739 19828 15748
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 15162 19748 15302
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19520 14716 19828 14725
rect 19520 14714 19526 14716
rect 19582 14714 19606 14716
rect 19662 14714 19686 14716
rect 19742 14714 19766 14716
rect 19822 14714 19828 14716
rect 19582 14662 19584 14714
rect 19764 14662 19766 14714
rect 19520 14660 19526 14662
rect 19582 14660 19606 14662
rect 19662 14660 19686 14662
rect 19742 14660 19766 14662
rect 19822 14660 19828 14662
rect 19520 14651 19828 14660
rect 19524 14408 19576 14414
rect 19444 14368 19524 14396
rect 19524 14350 19576 14356
rect 19352 13938 19656 13954
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19352 13932 19668 13938
rect 19352 13926 19616 13932
rect 18892 13326 18920 13874
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18708 11694 18736 12038
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 18328 11076 18380 11082
rect 18328 11018 18380 11024
rect 18524 10810 18552 11086
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 8430 18184 8774
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 18064 7546 18092 7890
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17972 6934 18000 7142
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 5914 17816 6598
rect 18064 6322 18092 6802
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 16684 2746 16804 2774
rect 16776 800 16804 2746
rect 17420 800 17448 4082
rect 18064 800 18092 6258
rect 18156 4146 18184 8366
rect 18248 5710 18276 9318
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8362 18460 8910
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18340 7410 18368 7686
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18432 6322 18460 8298
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18708 800 18736 11630
rect 18892 11150 18920 13262
rect 19352 12434 19380 13926
rect 19616 13874 19668 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13462 19472 13806
rect 19520 13628 19828 13637
rect 19520 13626 19526 13628
rect 19582 13626 19606 13628
rect 19662 13626 19686 13628
rect 19742 13626 19766 13628
rect 19822 13626 19828 13628
rect 19582 13574 19584 13626
rect 19764 13574 19766 13626
rect 19520 13572 19526 13574
rect 19582 13572 19606 13574
rect 19662 13572 19686 13574
rect 19742 13572 19766 13574
rect 19822 13572 19828 13574
rect 19520 13563 19828 13572
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19996 12986 20024 15506
rect 20088 14414 20116 16662
rect 20180 16348 20488 16357
rect 20180 16346 20186 16348
rect 20242 16346 20266 16348
rect 20322 16346 20346 16348
rect 20402 16346 20426 16348
rect 20482 16346 20488 16348
rect 20242 16294 20244 16346
rect 20424 16294 20426 16346
rect 20180 16292 20186 16294
rect 20242 16292 20266 16294
rect 20322 16292 20346 16294
rect 20402 16292 20426 16294
rect 20482 16292 20488 16294
rect 20180 16283 20488 16292
rect 20548 16114 20576 16730
rect 20640 16522 20668 18022
rect 20916 17202 20944 18226
rect 21008 17202 21036 18226
rect 21100 17338 21128 20334
rect 21180 19916 21232 19922
rect 21180 19858 21232 19864
rect 21192 19310 21220 19858
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21100 16794 21128 17274
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15434 20208 15846
rect 20168 15428 20220 15434
rect 20168 15370 20220 15376
rect 20180 15260 20488 15269
rect 20180 15258 20186 15260
rect 20242 15258 20266 15260
rect 20322 15258 20346 15260
rect 20402 15258 20426 15260
rect 20482 15258 20488 15260
rect 20242 15206 20244 15258
rect 20424 15206 20426 15258
rect 20180 15204 20186 15206
rect 20242 15204 20266 15206
rect 20322 15204 20346 15206
rect 20402 15204 20426 15206
rect 20482 15204 20488 15206
rect 20180 15195 20488 15204
rect 20548 14618 20576 16050
rect 21008 15706 21036 16594
rect 21088 16516 21140 16522
rect 21088 16458 21140 16464
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21008 15366 21036 15642
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 15162 21036 15302
rect 21100 15162 21128 16458
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 20180 14172 20488 14181
rect 20180 14170 20186 14172
rect 20242 14170 20266 14172
rect 20322 14170 20346 14172
rect 20402 14170 20426 14172
rect 20482 14170 20488 14172
rect 20242 14118 20244 14170
rect 20424 14118 20426 14170
rect 20180 14116 20186 14118
rect 20242 14116 20266 14118
rect 20322 14116 20346 14118
rect 20402 14116 20426 14118
rect 20482 14116 20488 14118
rect 20180 14107 20488 14116
rect 20824 13394 20852 14894
rect 21100 14822 21128 15098
rect 21192 14890 21220 15302
rect 21376 14958 21404 15438
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 13938 21128 14758
rect 21376 14618 21404 14894
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21468 14006 21496 20334
rect 21836 16454 21864 20538
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21928 19378 21956 19450
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21824 16448 21876 16454
rect 21824 16390 21876 16396
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21652 15706 21680 15846
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21652 15570 21680 15642
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21836 15162 21864 16390
rect 21928 15978 21956 16594
rect 22020 16538 22048 20726
rect 22112 20602 22140 21966
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22204 20942 22232 21830
rect 22296 21486 22324 21830
rect 22572 21690 22600 21898
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22848 21554 22876 21898
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22296 21078 22324 21422
rect 23032 21078 23060 21490
rect 23124 21146 23152 21490
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22848 20602 22876 21014
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22848 19854 22876 20198
rect 22940 19922 22968 20334
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22940 19310 22968 19858
rect 23032 19786 23060 20402
rect 23400 19854 23428 20402
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23020 19780 23072 19786
rect 23020 19722 23072 19728
rect 23032 19378 23060 19722
rect 23400 19446 23428 19790
rect 23492 19718 23520 20334
rect 23860 20330 23888 21422
rect 23848 20324 23900 20330
rect 23848 20266 23900 20272
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 22928 19304 22980 19310
rect 22928 19246 22980 19252
rect 22940 18834 22968 19246
rect 22928 18828 22980 18834
rect 22928 18770 22980 18776
rect 22940 18290 22968 18770
rect 23032 18766 23060 19314
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23020 18760 23072 18766
rect 23020 18702 23072 18708
rect 23032 18290 23060 18702
rect 22928 18284 22980 18290
rect 22928 18226 22980 18232
rect 23020 18284 23072 18290
rect 23020 18226 23072 18232
rect 22940 17746 22968 18226
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 23032 17678 23060 18226
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23020 16992 23072 16998
rect 23020 16934 23072 16940
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23032 16726 23060 16934
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 23124 16590 23152 16934
rect 23112 16584 23164 16590
rect 22020 16522 22140 16538
rect 23112 16526 23164 16532
rect 22008 16516 22140 16522
rect 22060 16510 22140 16516
rect 22008 16458 22060 16464
rect 22112 16046 22140 16510
rect 23216 16250 23244 17002
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23308 16096 23336 19110
rect 23400 18698 23428 19382
rect 23492 19378 23520 19654
rect 23952 19378 23980 23122
rect 24412 23050 24440 23530
rect 24504 23186 24532 23598
rect 24872 23322 24900 23598
rect 25424 23322 25452 23734
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 26948 23420 27256 23429
rect 26948 23418 26954 23420
rect 27010 23418 27034 23420
rect 27090 23418 27114 23420
rect 27170 23418 27194 23420
rect 27250 23418 27256 23420
rect 27010 23366 27012 23418
rect 27192 23366 27194 23418
rect 26948 23364 26954 23366
rect 27010 23364 27034 23366
rect 27090 23364 27114 23366
rect 27170 23364 27194 23366
rect 27250 23364 27256 23366
rect 26948 23355 27256 23364
rect 27448 23322 27476 23462
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24228 22710 24256 22918
rect 25148 22778 25176 23054
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 25136 22772 25188 22778
rect 25136 22714 25188 22720
rect 24216 22704 24268 22710
rect 24216 22646 24268 22652
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 24044 21486 24072 21966
rect 24228 21622 24256 22646
rect 24780 22506 24808 22646
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24768 22500 24820 22506
rect 24768 22442 24820 22448
rect 25056 22234 25084 22578
rect 25044 22228 25096 22234
rect 25044 22170 25096 22176
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21690 24440 21830
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23492 18766 23520 19314
rect 23848 18896 23900 18902
rect 23848 18838 23900 18844
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18290 23428 18634
rect 23492 18578 23520 18702
rect 23492 18550 23612 18578
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23400 17610 23428 18226
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23388 17604 23440 17610
rect 23388 17546 23440 17552
rect 23492 17270 23520 18022
rect 23584 17678 23612 18550
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23676 16590 23704 17138
rect 23768 16726 23796 17138
rect 23756 16720 23808 16726
rect 23756 16662 23808 16668
rect 23664 16584 23716 16590
rect 23664 16526 23716 16532
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23216 16068 23336 16096
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21732 15020 21784 15026
rect 21836 15008 21864 15098
rect 21928 15026 21956 15370
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 21784 14980 21864 15008
rect 21916 15020 21968 15026
rect 21732 14962 21784 14968
rect 21916 14962 21968 14968
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21928 14414 21956 14962
rect 21916 14408 21968 14414
rect 21836 14368 21916 14396
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 21008 13326 21036 13874
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20180 13084 20488 13093
rect 20180 13082 20186 13084
rect 20242 13082 20266 13084
rect 20322 13082 20346 13084
rect 20402 13082 20426 13084
rect 20482 13082 20488 13084
rect 20242 13030 20244 13082
rect 20424 13030 20426 13082
rect 20180 13028 20186 13030
rect 20242 13028 20266 13030
rect 20322 13028 20346 13030
rect 20402 13028 20426 13030
rect 20482 13028 20488 13030
rect 20180 13019 20488 13028
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19520 12540 19828 12549
rect 19520 12538 19526 12540
rect 19582 12538 19606 12540
rect 19662 12538 19686 12540
rect 19742 12538 19766 12540
rect 19822 12538 19828 12540
rect 19582 12486 19584 12538
rect 19764 12486 19766 12538
rect 19520 12484 19526 12486
rect 19582 12484 19606 12486
rect 19662 12484 19686 12486
rect 19742 12484 19766 12486
rect 19822 12484 19828 12486
rect 19520 12475 19828 12484
rect 19260 12406 19380 12434
rect 19260 12238 19288 12406
rect 19996 12306 20024 12922
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19984 12300 20036 12306
rect 20036 12260 20116 12288
rect 19984 12242 20036 12248
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 19260 10538 19288 12174
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 19352 10130 19380 12242
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19996 11898 20024 12106
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11762 20116 12260
rect 20180 11996 20488 12005
rect 20180 11994 20186 11996
rect 20242 11994 20266 11996
rect 20322 11994 20346 11996
rect 20402 11994 20426 11996
rect 20482 11994 20488 11996
rect 20242 11942 20244 11994
rect 20424 11942 20426 11994
rect 20180 11940 20186 11942
rect 20242 11940 20266 11942
rect 20322 11940 20346 11942
rect 20402 11940 20426 11942
rect 20482 11940 20488 11942
rect 20180 11931 20488 11940
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19444 10674 19472 11494
rect 19520 11452 19828 11461
rect 19520 11450 19526 11452
rect 19582 11450 19606 11452
rect 19662 11450 19686 11452
rect 19742 11450 19766 11452
rect 19822 11450 19828 11452
rect 19582 11398 19584 11450
rect 19764 11398 19766 11450
rect 19520 11396 19526 11398
rect 19582 11396 19606 11398
rect 19662 11396 19686 11398
rect 19742 11396 19766 11398
rect 19822 11396 19828 11398
rect 19520 11387 19828 11396
rect 19996 11218 20024 11494
rect 19984 11212 20036 11218
rect 19984 11154 20036 11160
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19904 10742 19932 11018
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19892 10736 19944 10742
rect 19892 10678 19944 10684
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 19168 9722 19196 9862
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18800 7954 18828 8026
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18800 7410 18828 7890
rect 19444 7886 19472 10610
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19520 10364 19828 10373
rect 19520 10362 19526 10364
rect 19582 10362 19606 10364
rect 19662 10362 19686 10364
rect 19742 10362 19766 10364
rect 19822 10362 19828 10364
rect 19582 10310 19584 10362
rect 19764 10310 19766 10362
rect 19520 10308 19526 10310
rect 19582 10308 19606 10310
rect 19662 10308 19686 10310
rect 19742 10308 19766 10310
rect 19822 10308 19828 10310
rect 19520 10299 19828 10308
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19536 9382 19564 9998
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19520 9276 19828 9285
rect 19520 9274 19526 9276
rect 19582 9274 19606 9276
rect 19662 9274 19686 9276
rect 19742 9274 19766 9276
rect 19822 9274 19828 9276
rect 19582 9222 19584 9274
rect 19764 9222 19766 9274
rect 19520 9220 19526 9222
rect 19582 9220 19606 9222
rect 19662 9220 19686 9222
rect 19742 9220 19766 9222
rect 19822 9220 19828 9222
rect 19520 9211 19828 9220
rect 19904 9058 19932 10406
rect 19812 9030 19932 9058
rect 19812 8294 19840 9030
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19520 8188 19828 8197
rect 19520 8186 19526 8188
rect 19582 8186 19606 8188
rect 19662 8186 19686 8188
rect 19742 8186 19766 8188
rect 19822 8186 19828 8188
rect 19582 8134 19584 8186
rect 19764 8134 19766 8186
rect 19520 8132 19526 8134
rect 19582 8132 19606 8134
rect 19662 8132 19686 8134
rect 19742 8132 19766 8134
rect 19822 8132 19828 8134
rect 19520 8123 19828 8132
rect 19904 8090 19932 8366
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19444 7410 19472 7822
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 7410 19748 7686
rect 19812 7410 19840 7890
rect 19996 7886 20024 10746
rect 20088 10674 20116 10950
rect 20180 10908 20488 10917
rect 20180 10906 20186 10908
rect 20242 10906 20266 10908
rect 20322 10906 20346 10908
rect 20402 10906 20426 10908
rect 20482 10906 20488 10908
rect 20242 10854 20244 10906
rect 20424 10854 20426 10906
rect 20180 10852 20186 10854
rect 20242 10852 20266 10854
rect 20322 10852 20346 10854
rect 20402 10852 20426 10854
rect 20482 10852 20488 10854
rect 20180 10843 20488 10852
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 7886 20116 10610
rect 20548 10130 20576 12854
rect 20640 11762 20668 13126
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 21100 11694 21128 13330
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21376 12442 21404 13194
rect 21548 12640 21600 12646
rect 21548 12582 21600 12588
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21560 12238 21588 12582
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21744 11898 21772 12174
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20640 10010 20668 10950
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 21008 10146 21036 11630
rect 21192 11354 21220 11630
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21100 10606 21128 11290
rect 21836 11286 21864 14368
rect 21916 14350 21968 14356
rect 22020 14346 22048 14962
rect 22112 14482 22140 15302
rect 22296 14822 22324 15438
rect 22480 15094 22508 15642
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22652 15156 22704 15162
rect 22652 15098 22704 15104
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22480 14550 22508 15030
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22020 13802 22048 14282
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 22112 13274 22140 13874
rect 22204 13394 22232 14214
rect 22296 13394 22324 14282
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 22112 13246 22232 13274
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11898 21956 12038
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 22204 11778 22232 13246
rect 22296 12986 22324 13330
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12986 22508 13262
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22296 11880 22324 12922
rect 22296 11852 22508 11880
rect 22204 11750 22416 11778
rect 21824 11280 21876 11286
rect 21824 11222 21876 11228
rect 22388 11150 22416 11750
rect 22192 11144 22244 11150
rect 21822 11112 21878 11121
rect 22192 11086 22244 11092
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 21822 11047 21824 11056
rect 21876 11047 21878 11056
rect 21824 11018 21876 11024
rect 21836 10742 21864 11018
rect 22204 10810 22232 11086
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 20548 9982 20668 10010
rect 20180 9820 20488 9829
rect 20180 9818 20186 9820
rect 20242 9818 20266 9820
rect 20322 9818 20346 9820
rect 20402 9818 20426 9820
rect 20482 9818 20488 9820
rect 20242 9766 20244 9818
rect 20424 9766 20426 9818
rect 20180 9764 20186 9766
rect 20242 9764 20266 9766
rect 20322 9764 20346 9766
rect 20402 9764 20426 9766
rect 20482 9764 20488 9766
rect 20180 9755 20488 9764
rect 20548 9382 20576 9982
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20180 8732 20488 8741
rect 20180 8730 20186 8732
rect 20242 8730 20266 8732
rect 20322 8730 20346 8732
rect 20402 8730 20426 8732
rect 20482 8730 20488 8732
rect 20242 8678 20244 8730
rect 20424 8678 20426 8730
rect 20180 8676 20186 8678
rect 20242 8676 20266 8678
rect 20322 8676 20346 8678
rect 20402 8676 20426 8678
rect 20482 8676 20488 8678
rect 20180 8667 20488 8676
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 7954 20300 8230
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 18800 6866 18828 7346
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 19444 6798 19472 7346
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19520 7100 19828 7109
rect 19520 7098 19526 7100
rect 19582 7098 19606 7100
rect 19662 7098 19686 7100
rect 19742 7098 19766 7100
rect 19822 7098 19828 7100
rect 19582 7046 19584 7098
rect 19764 7046 19766 7098
rect 19520 7044 19526 7046
rect 19582 7044 19606 7046
rect 19662 7044 19686 7046
rect 19742 7044 19766 7046
rect 19822 7044 19828 7046
rect 19520 7035 19828 7044
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19444 5914 19472 6190
rect 19520 6012 19828 6021
rect 19520 6010 19526 6012
rect 19582 6010 19606 6012
rect 19662 6010 19686 6012
rect 19742 6010 19766 6012
rect 19822 6010 19828 6012
rect 19582 5958 19584 6010
rect 19764 5958 19766 6010
rect 19520 5956 19526 5958
rect 19582 5956 19606 5958
rect 19662 5956 19686 5958
rect 19742 5956 19766 5958
rect 19822 5956 19828 5958
rect 19520 5947 19828 5956
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19904 5710 19932 7142
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19520 4924 19828 4933
rect 19520 4922 19526 4924
rect 19582 4922 19606 4924
rect 19662 4922 19686 4924
rect 19742 4922 19766 4924
rect 19822 4922 19828 4924
rect 19582 4870 19584 4922
rect 19764 4870 19766 4922
rect 19520 4868 19526 4870
rect 19582 4868 19606 4870
rect 19662 4868 19686 4870
rect 19742 4868 19766 4870
rect 19822 4868 19828 4870
rect 19520 4859 19828 4868
rect 19520 3836 19828 3845
rect 19520 3834 19526 3836
rect 19582 3834 19606 3836
rect 19662 3834 19686 3836
rect 19742 3834 19766 3836
rect 19822 3834 19828 3836
rect 19582 3782 19584 3834
rect 19764 3782 19766 3834
rect 19520 3780 19526 3782
rect 19582 3780 19606 3782
rect 19662 3780 19686 3782
rect 19742 3780 19766 3782
rect 19822 3780 19828 3782
rect 19520 3771 19828 3780
rect 19520 2748 19828 2757
rect 19520 2746 19526 2748
rect 19582 2746 19606 2748
rect 19662 2746 19686 2748
rect 19742 2746 19766 2748
rect 19822 2746 19828 2748
rect 19582 2694 19584 2746
rect 19764 2694 19766 2746
rect 19520 2692 19526 2694
rect 19582 2692 19606 2694
rect 19662 2692 19686 2694
rect 19742 2692 19766 2694
rect 19822 2692 19828 2694
rect 19520 2683 19828 2692
rect 19996 800 20024 7686
rect 20180 7644 20488 7653
rect 20180 7642 20186 7644
rect 20242 7642 20266 7644
rect 20322 7642 20346 7644
rect 20402 7642 20426 7644
rect 20482 7642 20488 7644
rect 20242 7590 20244 7642
rect 20424 7590 20426 7642
rect 20180 7588 20186 7590
rect 20242 7588 20266 7590
rect 20322 7588 20346 7590
rect 20402 7588 20426 7590
rect 20482 7588 20488 7590
rect 20180 7579 20488 7588
rect 20548 7546 20576 8502
rect 20640 7546 20668 9862
rect 20824 9042 20852 10134
rect 20916 9994 20944 10134
rect 21008 10118 21220 10146
rect 22020 10130 22048 10610
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 10266 22324 10406
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 21192 10062 21220 10118
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 22020 9042 22048 10066
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21744 8634 21772 8910
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20824 7886 20852 8366
rect 22020 8294 22048 8978
rect 22388 8974 22416 9998
rect 22480 9450 22508 11852
rect 22664 11150 22692 15098
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 14074 22784 14214
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22848 13802 22876 15438
rect 23216 15366 23244 16068
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23308 15706 23336 15846
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23400 15586 23428 16390
rect 23492 16114 23520 16390
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23492 15586 23520 15642
rect 23296 15564 23348 15570
rect 23400 15558 23520 15586
rect 23400 15552 23428 15558
rect 23348 15524 23428 15552
rect 23296 15506 23348 15512
rect 23204 15360 23256 15366
rect 23124 15320 23204 15348
rect 23124 14618 23152 15320
rect 23204 15302 23256 15308
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23204 14272 23256 14278
rect 23204 14214 23256 14220
rect 23216 13938 23244 14214
rect 23204 13932 23256 13938
rect 23480 13932 23532 13938
rect 23256 13892 23480 13920
rect 23204 13874 23256 13880
rect 23480 13874 23532 13880
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22756 13394 22784 13670
rect 22848 13394 22876 13738
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23492 13394 23520 13466
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23584 12850 23612 16050
rect 23768 15638 23796 16662
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23860 15434 23888 18838
rect 23952 18290 23980 19314
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24044 17542 24072 21422
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 20058 24164 20810
rect 25240 20534 25268 22986
rect 25504 22636 25556 22642
rect 25504 22578 25556 22584
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25320 21956 25372 21962
rect 25320 21898 25372 21904
rect 25332 21486 25360 21898
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25044 20528 25096 20534
rect 25044 20470 25096 20476
rect 25228 20528 25280 20534
rect 25228 20470 25280 20476
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24228 19446 24256 19722
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 24504 19514 24532 19654
rect 24492 19508 24544 19514
rect 24492 19450 24544 19456
rect 24964 19446 24992 20198
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 18426 24440 18566
rect 24596 18426 24624 18702
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24872 17882 24900 18294
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 25056 17678 25084 20470
rect 25424 19990 25452 22510
rect 25516 22166 25544 22578
rect 26056 22432 26108 22438
rect 26056 22374 26108 22380
rect 27344 22432 27396 22438
rect 27344 22374 27396 22380
rect 25504 22160 25556 22166
rect 25504 22102 25556 22108
rect 25516 21010 25544 22102
rect 26068 22080 26096 22374
rect 26948 22332 27256 22341
rect 26948 22330 26954 22332
rect 27010 22330 27034 22332
rect 27090 22330 27114 22332
rect 27170 22330 27194 22332
rect 27250 22330 27256 22332
rect 27010 22278 27012 22330
rect 27192 22278 27194 22330
rect 26948 22276 26954 22278
rect 27010 22276 27034 22278
rect 27090 22276 27114 22278
rect 27170 22276 27194 22278
rect 27250 22276 27256 22278
rect 26948 22267 27256 22276
rect 26240 22092 26292 22098
rect 27356 22094 27384 22374
rect 27448 22234 27476 23258
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 27608 22876 27916 22885
rect 27608 22874 27614 22876
rect 27670 22874 27694 22876
rect 27750 22874 27774 22876
rect 27830 22874 27854 22876
rect 27910 22874 27916 22876
rect 27670 22822 27672 22874
rect 27852 22822 27854 22874
rect 27608 22820 27614 22822
rect 27670 22820 27694 22822
rect 27750 22820 27774 22822
rect 27830 22820 27854 22822
rect 27910 22820 27916 22822
rect 27608 22811 27916 22820
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 26068 22052 26240 22080
rect 26068 21570 26096 22052
rect 26240 22034 26292 22040
rect 27264 22066 27384 22094
rect 27264 22030 27292 22066
rect 26332 22024 26384 22030
rect 26330 21992 26332 22001
rect 26884 22024 26936 22030
rect 26384 21992 26386 22001
rect 26804 21984 26884 22012
rect 26240 21956 26292 21962
rect 26386 21950 26556 21978
rect 26330 21927 26386 21936
rect 26240 21898 26292 21904
rect 26252 21706 26280 21898
rect 26160 21690 26372 21706
rect 26148 21684 26372 21690
rect 26200 21678 26372 21684
rect 26148 21626 26200 21632
rect 25872 21548 25924 21554
rect 26068 21542 26280 21570
rect 25872 21490 25924 21496
rect 25884 21049 25912 21490
rect 25870 21040 25926 21049
rect 25504 21004 25556 21010
rect 25870 20975 25926 20984
rect 25504 20946 25556 20952
rect 25412 19984 25464 19990
rect 25412 19926 25464 19932
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19514 25268 19654
rect 25228 19508 25280 19514
rect 25228 19450 25280 19456
rect 25424 18222 25452 19926
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25792 19446 25820 19858
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 26252 19310 26280 21542
rect 26344 21536 26372 21678
rect 26424 21548 26476 21554
rect 26344 21508 26424 21536
rect 26424 21490 26476 21496
rect 26528 19446 26556 21950
rect 26804 21622 26832 21984
rect 26884 21966 26936 21972
rect 27252 22024 27304 22030
rect 27252 21966 27304 21972
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 26792 21616 26844 21622
rect 26792 21558 26844 21564
rect 26608 21412 26660 21418
rect 26608 21354 26660 21360
rect 26620 21010 26648 21354
rect 26804 21146 26832 21558
rect 26896 21486 26924 21830
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26884 21480 26936 21486
rect 26884 21422 26936 21428
rect 26988 21350 27016 21490
rect 27264 21350 27292 21966
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 26948 21244 27256 21253
rect 26948 21242 26954 21244
rect 27010 21242 27034 21244
rect 27090 21242 27114 21244
rect 27170 21242 27194 21244
rect 27250 21242 27256 21244
rect 27010 21190 27012 21242
rect 27192 21190 27194 21242
rect 26948 21188 26954 21190
rect 27010 21188 27034 21190
rect 27090 21188 27114 21190
rect 27170 21188 27194 21190
rect 27250 21188 27256 21190
rect 26948 21179 27256 21188
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26792 21140 26844 21146
rect 26792 21082 26844 21088
rect 26608 21004 26660 21010
rect 26608 20946 26660 20952
rect 26712 20534 26740 21082
rect 27158 21040 27214 21049
rect 27158 20975 27160 20984
rect 27212 20975 27214 20984
rect 27160 20946 27212 20952
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26804 20602 26832 20878
rect 27160 20868 27212 20874
rect 27160 20810 27212 20816
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26700 20528 26752 20534
rect 26700 20470 26752 20476
rect 26804 19514 26832 20538
rect 27172 20482 27200 20810
rect 27356 20602 27384 21490
rect 27540 21146 27568 22714
rect 27896 22228 27948 22234
rect 28000 22216 28028 23054
rect 28908 22976 28960 22982
rect 28908 22918 28960 22924
rect 28920 22778 28948 22918
rect 28908 22772 28960 22778
rect 28908 22714 28960 22720
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 27948 22188 28028 22216
rect 27896 22170 27948 22176
rect 27608 21788 27916 21797
rect 27608 21786 27614 21788
rect 27670 21786 27694 21788
rect 27750 21786 27774 21788
rect 27830 21786 27854 21788
rect 27910 21786 27916 21788
rect 27670 21734 27672 21786
rect 27852 21734 27854 21786
rect 27608 21732 27614 21734
rect 27670 21732 27694 21734
rect 27750 21732 27774 21734
rect 27830 21732 27854 21734
rect 27910 21732 27916 21734
rect 27608 21723 27916 21732
rect 28000 21622 28028 22188
rect 28184 22166 28212 22578
rect 28816 22500 28868 22506
rect 28816 22442 28868 22448
rect 28632 22432 28684 22438
rect 28632 22374 28684 22380
rect 28172 22160 28224 22166
rect 28172 22102 28224 22108
rect 28644 22094 28672 22374
rect 28828 22166 28856 22442
rect 29092 22432 29144 22438
rect 29092 22374 29144 22380
rect 29276 22432 29328 22438
rect 29276 22374 29328 22380
rect 28816 22160 28868 22166
rect 28816 22102 28868 22108
rect 28460 22066 28672 22094
rect 28080 21888 28132 21894
rect 28078 21856 28080 21865
rect 28132 21856 28134 21865
rect 28078 21791 28134 21800
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27988 21072 28040 21078
rect 27988 21014 28040 21020
rect 27608 20700 27916 20709
rect 27608 20698 27614 20700
rect 27670 20698 27694 20700
rect 27750 20698 27774 20700
rect 27830 20698 27854 20700
rect 27910 20698 27916 20700
rect 27670 20646 27672 20698
rect 27852 20646 27854 20698
rect 27608 20644 27614 20646
rect 27670 20644 27694 20646
rect 27750 20644 27774 20646
rect 27830 20644 27854 20646
rect 27910 20644 27916 20646
rect 27608 20635 27916 20644
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27618 20496 27674 20505
rect 27172 20454 27384 20482
rect 26948 20156 27256 20165
rect 26948 20154 26954 20156
rect 27010 20154 27034 20156
rect 27090 20154 27114 20156
rect 27170 20154 27194 20156
rect 27250 20154 27256 20156
rect 27010 20102 27012 20154
rect 27192 20102 27194 20154
rect 26948 20100 26954 20102
rect 27010 20100 27034 20102
rect 27090 20100 27114 20102
rect 27170 20100 27194 20102
rect 27250 20100 27256 20102
rect 26948 20091 27256 20100
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26516 19440 26568 19446
rect 26516 19382 26568 19388
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 26424 19372 26476 19378
rect 26424 19314 26476 19320
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26344 18970 26372 19314
rect 26332 18964 26384 18970
rect 26332 18906 26384 18912
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24032 17536 24084 17542
rect 24032 17478 24084 17484
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23952 15706 23980 16390
rect 24872 16250 24900 16594
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23676 14074 23704 14554
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23768 13530 23796 14962
rect 23860 14346 23888 15370
rect 23952 14618 23980 15438
rect 24320 15026 24348 15506
rect 24964 15502 24992 17274
rect 25056 16130 25084 17614
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25148 16250 25176 17138
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 16250 25452 16458
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25056 16114 25360 16130
rect 25044 16108 25372 16114
rect 25096 16102 25320 16108
rect 25044 16050 25096 16056
rect 25320 16050 25372 16056
rect 25976 15586 26004 18566
rect 26252 18426 26280 18566
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 26068 17354 26096 18158
rect 26160 17542 26188 18226
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26068 17326 26188 17354
rect 26436 17338 26464 19314
rect 26884 19304 26936 19310
rect 26884 19246 26936 19252
rect 26896 19122 26924 19246
rect 27356 19174 27384 20454
rect 27618 20431 27674 20440
rect 27632 20058 27660 20431
rect 27620 20052 27672 20058
rect 28000 20040 28028 21014
rect 28460 20942 28488 22066
rect 28828 22030 28856 22102
rect 29104 22030 29132 22374
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 29092 22024 29144 22030
rect 29092 21966 29144 21972
rect 28644 21078 28672 21966
rect 29288 21962 29316 22374
rect 29276 21956 29328 21962
rect 29276 21898 29328 21904
rect 28632 21072 28684 21078
rect 28632 21014 28684 21020
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28552 20398 28580 20878
rect 28644 20602 28672 21014
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 28816 20596 28868 20602
rect 28816 20538 28868 20544
rect 28540 20392 28592 20398
rect 28540 20334 28592 20340
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 20058 28212 20198
rect 28172 20052 28224 20058
rect 28000 20012 28120 20040
rect 27620 19994 27672 20000
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 27608 19612 27916 19621
rect 27608 19610 27614 19612
rect 27670 19610 27694 19612
rect 27750 19610 27774 19612
rect 27830 19610 27854 19612
rect 27910 19610 27916 19612
rect 27670 19558 27672 19610
rect 27852 19558 27854 19610
rect 27608 19556 27614 19558
rect 27670 19556 27694 19558
rect 27750 19556 27774 19558
rect 27830 19556 27854 19558
rect 27910 19556 27916 19558
rect 27608 19547 27916 19556
rect 28000 19378 28028 19858
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 26804 19094 26924 19122
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 27896 19168 27948 19174
rect 27948 19128 28028 19156
rect 27896 19110 27948 19116
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26160 16522 26188 17326
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26528 16522 26556 18770
rect 26804 18290 26832 19094
rect 26948 19068 27256 19077
rect 26948 19066 26954 19068
rect 27010 19066 27034 19068
rect 27090 19066 27114 19068
rect 27170 19066 27194 19068
rect 27250 19066 27256 19068
rect 27010 19014 27012 19066
rect 27192 19014 27194 19066
rect 26948 19012 26954 19014
rect 27010 19012 27034 19014
rect 27090 19012 27114 19014
rect 27170 19012 27194 19014
rect 27250 19012 27256 19014
rect 26948 19003 27256 19012
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27344 18352 27396 18358
rect 27344 18294 27396 18300
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26804 16794 26832 18226
rect 26948 17980 27256 17989
rect 26948 17978 26954 17980
rect 27010 17978 27034 17980
rect 27090 17978 27114 17980
rect 27170 17978 27194 17980
rect 27250 17978 27256 17980
rect 27010 17926 27012 17978
rect 27192 17926 27194 17978
rect 26948 17924 26954 17926
rect 27010 17924 27034 17926
rect 27090 17924 27114 17926
rect 27170 17924 27194 17926
rect 27250 17924 27256 17926
rect 26948 17915 27256 17924
rect 27356 17746 27384 18294
rect 27448 18068 27476 18702
rect 27608 18524 27916 18533
rect 27608 18522 27614 18524
rect 27670 18522 27694 18524
rect 27750 18522 27774 18524
rect 27830 18522 27854 18524
rect 27910 18522 27916 18524
rect 27670 18470 27672 18522
rect 27852 18470 27854 18522
rect 27608 18468 27614 18470
rect 27670 18468 27694 18470
rect 27750 18468 27774 18470
rect 27830 18468 27854 18470
rect 27910 18468 27916 18470
rect 27608 18459 27916 18468
rect 28000 18358 28028 19128
rect 28092 18970 28120 20012
rect 28172 19994 28224 20000
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28276 19174 28304 19994
rect 28630 19816 28686 19825
rect 28828 19802 28856 20538
rect 29000 20528 29052 20534
rect 29288 20482 29316 21898
rect 29368 21888 29420 21894
rect 29368 21830 29420 21836
rect 29380 20942 29408 21830
rect 29368 20936 29420 20942
rect 29368 20878 29420 20884
rect 29052 20476 29316 20482
rect 29000 20470 29316 20476
rect 29012 20454 29316 20470
rect 28998 20360 29054 20369
rect 28998 20295 29000 20304
rect 29052 20295 29054 20304
rect 29092 20324 29144 20330
rect 29000 20266 29052 20272
rect 29092 20266 29144 20272
rect 28908 20256 28960 20262
rect 28908 20198 28960 20204
rect 28920 19922 28948 20198
rect 29104 20074 29132 20266
rect 29104 20046 29224 20074
rect 29092 19984 29144 19990
rect 29092 19926 29144 19932
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 28828 19774 28948 19802
rect 28630 19751 28632 19760
rect 28684 19751 28686 19760
rect 28632 19722 28684 19728
rect 28920 19174 28948 19774
rect 29104 19718 29132 19926
rect 29196 19768 29224 20046
rect 29288 19922 29316 20454
rect 29276 19916 29328 19922
rect 29276 19858 29328 19864
rect 29276 19780 29328 19786
rect 29196 19740 29276 19768
rect 29276 19722 29328 19728
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 29288 19242 29316 19722
rect 29380 19378 29408 20878
rect 29644 20800 29696 20806
rect 29644 20742 29696 20748
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29472 20058 29500 20402
rect 29552 20392 29604 20398
rect 29550 20360 29552 20369
rect 29604 20360 29606 20369
rect 29550 20295 29606 20304
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29656 19718 29684 20742
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 29644 19712 29696 19718
rect 29644 19654 29696 19660
rect 30116 19378 30144 20402
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30300 20058 30328 20198
rect 30288 20052 30340 20058
rect 30288 19994 30340 20000
rect 30300 19514 30328 19994
rect 30288 19508 30340 19514
rect 30288 19450 30340 19456
rect 29368 19372 29420 19378
rect 29368 19314 29420 19320
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 29276 19236 29328 19242
rect 29276 19178 29328 19184
rect 28264 19168 28316 19174
rect 28264 19110 28316 19116
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28908 19168 28960 19174
rect 28908 19110 28960 19116
rect 29184 19168 29236 19174
rect 29184 19110 29236 19116
rect 28080 18964 28132 18970
rect 28080 18906 28132 18912
rect 28092 18748 28120 18906
rect 28172 18760 28224 18766
rect 28092 18720 28172 18748
rect 28172 18702 28224 18708
rect 28276 18630 28304 19110
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 27988 18352 28040 18358
rect 27988 18294 28040 18300
rect 28172 18352 28224 18358
rect 28172 18294 28224 18300
rect 27528 18080 27580 18086
rect 27448 18040 27528 18068
rect 27448 17882 27476 18040
rect 27528 18022 27580 18028
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 27632 17785 27660 17818
rect 27618 17776 27674 17785
rect 27344 17740 27396 17746
rect 27618 17711 27674 17720
rect 27344 17682 27396 17688
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 27608 17436 27916 17445
rect 27608 17434 27614 17436
rect 27670 17434 27694 17436
rect 27750 17434 27774 17436
rect 27830 17434 27854 17436
rect 27910 17434 27916 17436
rect 27670 17382 27672 17434
rect 27852 17382 27854 17434
rect 27608 17380 27614 17382
rect 27670 17380 27694 17382
rect 27750 17380 27774 17382
rect 27830 17380 27854 17382
rect 27910 17380 27916 17382
rect 27608 17371 27916 17380
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 26948 16892 27256 16901
rect 26948 16890 26954 16892
rect 27010 16890 27034 16892
rect 27090 16890 27114 16892
rect 27170 16890 27194 16892
rect 27250 16890 27256 16892
rect 27010 16838 27012 16890
rect 27192 16838 27194 16890
rect 26948 16836 26954 16838
rect 27010 16836 27034 16838
rect 27090 16836 27114 16838
rect 27170 16836 27194 16838
rect 27250 16836 27256 16838
rect 26948 16827 27256 16836
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26148 16516 26200 16522
rect 26148 16458 26200 16464
rect 26516 16516 26568 16522
rect 26516 16458 26568 16464
rect 26160 16046 26188 16458
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26252 16114 26280 16390
rect 26804 16114 26832 16730
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27448 16182 27476 16594
rect 27540 16522 27568 17138
rect 27802 17096 27858 17105
rect 27802 17031 27804 17040
rect 27856 17031 27858 17040
rect 27804 17002 27856 17008
rect 28000 16794 28028 17614
rect 28092 17610 28120 18022
rect 28184 17882 28212 18294
rect 28172 17876 28224 17882
rect 28172 17818 28224 17824
rect 28080 17604 28132 17610
rect 28080 17546 28132 17552
rect 28092 16998 28120 17546
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 27528 16516 27580 16522
rect 27528 16458 27580 16464
rect 27436 16176 27488 16182
rect 27436 16118 27488 16124
rect 27540 16130 27568 16458
rect 27608 16348 27916 16357
rect 27608 16346 27614 16348
rect 27670 16346 27694 16348
rect 27750 16346 27774 16348
rect 27830 16346 27854 16348
rect 27910 16346 27916 16348
rect 27670 16294 27672 16346
rect 27852 16294 27854 16346
rect 27608 16292 27614 16294
rect 27670 16292 27694 16294
rect 27750 16292 27774 16294
rect 27830 16292 27854 16294
rect 27910 16292 27916 16294
rect 27608 16283 27916 16292
rect 27540 16114 27660 16130
rect 28000 16114 28028 16730
rect 28184 16504 28212 17138
rect 28276 17134 28304 18566
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28264 16516 28316 16522
rect 28184 16476 28264 16504
rect 28264 16458 28316 16464
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 27540 16108 27672 16114
rect 27540 16102 27620 16108
rect 26056 16040 26108 16046
rect 26056 15982 26108 15988
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26068 15706 26096 15982
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25976 15558 26096 15586
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24320 14618 24348 14962
rect 25056 14618 25084 15302
rect 25608 15162 25636 15302
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 24044 13802 24072 14350
rect 24780 13938 24808 14350
rect 24964 14278 24992 14554
rect 25884 14550 25912 14962
rect 25976 14890 26004 15438
rect 26068 15026 26096 15558
rect 26344 15502 26372 15846
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26332 15496 26384 15502
rect 26332 15438 26384 15444
rect 26252 15162 26280 15438
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26712 15026 26740 16050
rect 26948 15804 27256 15813
rect 26948 15802 26954 15804
rect 27010 15802 27034 15804
rect 27090 15802 27114 15804
rect 27170 15802 27194 15804
rect 27250 15802 27256 15804
rect 27010 15750 27012 15802
rect 27192 15750 27194 15802
rect 26948 15748 26954 15750
rect 27010 15748 27034 15750
rect 27090 15748 27114 15750
rect 27170 15748 27194 15750
rect 27250 15748 27256 15750
rect 26948 15739 27256 15748
rect 27540 15502 27568 16102
rect 27620 16050 27672 16056
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 27620 15972 27672 15978
rect 27620 15914 27672 15920
rect 27632 15745 27660 15914
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 27618 15736 27674 15745
rect 27618 15671 27674 15680
rect 28184 15570 28212 15846
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28276 15502 28304 16458
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26700 15020 26752 15026
rect 26700 14962 26752 14968
rect 25964 14884 26016 14890
rect 25964 14826 26016 14832
rect 25872 14544 25924 14550
rect 25872 14486 25924 14492
rect 25044 14408 25096 14414
rect 25228 14408 25280 14414
rect 25096 14356 25228 14362
rect 25044 14350 25280 14356
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25056 14334 25268 14350
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24872 14074 24900 14214
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 23848 13796 23900 13802
rect 23848 13738 23900 13744
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23860 13394 23888 13738
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 24044 13326 24072 13738
rect 24768 13388 24820 13394
rect 24872 13376 24900 14010
rect 25056 14006 25084 14334
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 25332 13938 25360 14350
rect 25504 14340 25556 14346
rect 25504 14282 25556 14288
rect 25516 14074 25544 14282
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 24820 13348 24900 13376
rect 24768 13330 24820 13336
rect 25148 13326 25176 13670
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 24044 12850 24072 13262
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 24688 12850 24716 13126
rect 25516 12850 25544 13126
rect 25608 12986 25636 14350
rect 25884 14074 25912 14486
rect 26160 14414 26188 14962
rect 27540 14958 27568 15438
rect 27608 15260 27916 15269
rect 27608 15258 27614 15260
rect 27670 15258 27694 15260
rect 27750 15258 27774 15260
rect 27830 15258 27854 15260
rect 27910 15258 27916 15260
rect 27670 15206 27672 15258
rect 27852 15206 27854 15258
rect 27608 15204 27614 15206
rect 27670 15204 27694 15206
rect 27750 15204 27774 15206
rect 27830 15204 27854 15206
rect 27910 15204 27916 15206
rect 27608 15195 27916 15204
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 26948 14716 27256 14725
rect 26948 14714 26954 14716
rect 27010 14714 27034 14716
rect 27090 14714 27114 14716
rect 27170 14714 27194 14716
rect 27250 14714 27256 14716
rect 27010 14662 27012 14714
rect 27192 14662 27194 14714
rect 26948 14660 26954 14662
rect 27010 14660 27034 14662
rect 27090 14660 27114 14662
rect 27170 14660 27194 14662
rect 27250 14660 27256 14662
rect 26948 14651 27256 14660
rect 27724 14618 27752 14758
rect 28276 14618 28304 14758
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 26148 14408 26200 14414
rect 26148 14350 26200 14356
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26160 13734 26188 14214
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26252 13530 26280 13806
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26344 13326 26372 14214
rect 27608 14172 27916 14181
rect 27608 14170 27614 14172
rect 27670 14170 27694 14172
rect 27750 14170 27774 14172
rect 27830 14170 27854 14172
rect 27910 14170 27916 14172
rect 27670 14118 27672 14170
rect 27852 14118 27854 14170
rect 27608 14116 27614 14118
rect 27670 14116 27694 14118
rect 27750 14116 27774 14118
rect 27830 14116 27854 14118
rect 27910 14116 27916 14118
rect 27608 14107 27916 14116
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 27342 13696 27398 13705
rect 26528 13462 26556 13670
rect 26948 13628 27256 13637
rect 27342 13631 27398 13640
rect 26948 13626 26954 13628
rect 27010 13626 27034 13628
rect 27090 13626 27114 13628
rect 27170 13626 27194 13628
rect 27250 13626 27256 13628
rect 27010 13574 27012 13626
rect 27192 13574 27194 13626
rect 26948 13572 26954 13574
rect 27010 13572 27034 13574
rect 27090 13572 27114 13574
rect 27170 13572 27194 13574
rect 27250 13572 27256 13574
rect 26948 13563 27256 13572
rect 26516 13456 26568 13462
rect 26516 13398 26568 13404
rect 27356 13394 27384 13631
rect 28368 13530 28396 18566
rect 28460 18426 28488 18702
rect 28828 18698 28856 19110
rect 29196 18698 29224 19110
rect 29288 18902 29316 19178
rect 29276 18896 29328 18902
rect 29276 18838 29328 18844
rect 28816 18692 28868 18698
rect 28816 18634 28868 18640
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 28630 18456 28686 18465
rect 28448 18420 28500 18426
rect 29196 18426 29224 18634
rect 28630 18391 28686 18400
rect 29184 18420 29236 18426
rect 28448 18362 28500 18368
rect 28644 18358 28672 18391
rect 29184 18362 29236 18368
rect 30116 18358 30144 19314
rect 28632 18352 28684 18358
rect 28632 18294 28684 18300
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 29184 18284 29236 18290
rect 29184 18226 29236 18232
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 29196 17882 29224 18226
rect 30024 17882 30052 18226
rect 29184 17876 29236 17882
rect 29184 17818 29236 17824
rect 30012 17876 30064 17882
rect 30012 17818 30064 17824
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 16425 30420 16458
rect 30378 16416 30434 16425
rect 30378 16351 30434 16360
rect 28356 13524 28408 13530
rect 28356 13466 28408 13472
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23032 12238 23060 12718
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11830 23060 12038
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 23216 11014 23244 12786
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23860 11150 23888 11630
rect 23952 11286 23980 11698
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24320 11354 24348 11494
rect 25148 11354 25176 12718
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22572 10062 22600 10406
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22664 9722 22692 9862
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22572 9450 22600 9658
rect 22756 9586 22784 10542
rect 23032 10266 23060 10610
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23032 9926 23060 10202
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22756 8634 22784 9522
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22020 8090 22048 8230
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22388 8022 22416 8366
rect 22664 8022 22692 8434
rect 22376 8016 22428 8022
rect 22376 7958 22428 7964
rect 22652 8016 22704 8022
rect 22652 7958 22704 7964
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 7546 20760 7754
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20088 6730 20116 7482
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20180 6798 20208 7278
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 7002 20300 7142
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 20180 6556 20488 6565
rect 20180 6554 20186 6556
rect 20242 6554 20266 6556
rect 20322 6554 20346 6556
rect 20402 6554 20426 6556
rect 20482 6554 20488 6556
rect 20242 6502 20244 6554
rect 20424 6502 20426 6554
rect 20180 6500 20186 6502
rect 20242 6500 20266 6502
rect 20322 6500 20346 6502
rect 20402 6500 20426 6502
rect 20482 6500 20488 6502
rect 20180 6491 20488 6500
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20180 5914 20208 6326
rect 20548 6186 20576 7482
rect 22388 7478 22416 7958
rect 22376 7472 22428 7478
rect 22376 7414 22428 7420
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22020 7290 22048 7346
rect 21928 7262 22048 7290
rect 21928 6866 21956 7262
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21376 6746 21404 6802
rect 21284 6718 21404 6746
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20180 5468 20488 5477
rect 20180 5466 20186 5468
rect 20242 5466 20266 5468
rect 20322 5466 20346 5468
rect 20402 5466 20426 5468
rect 20482 5466 20488 5468
rect 20242 5414 20244 5466
rect 20424 5414 20426 5466
rect 20180 5412 20186 5414
rect 20242 5412 20266 5414
rect 20322 5412 20346 5414
rect 20402 5412 20426 5414
rect 20482 5412 20488 5414
rect 20180 5403 20488 5412
rect 20180 4380 20488 4389
rect 20180 4378 20186 4380
rect 20242 4378 20266 4380
rect 20322 4378 20346 4380
rect 20402 4378 20426 4380
rect 20482 4378 20488 4380
rect 20242 4326 20244 4378
rect 20424 4326 20426 4378
rect 20180 4324 20186 4326
rect 20242 4324 20266 4326
rect 20322 4324 20346 4326
rect 20402 4324 20426 4326
rect 20482 4324 20488 4326
rect 20180 4315 20488 4324
rect 20180 3292 20488 3301
rect 20180 3290 20186 3292
rect 20242 3290 20266 3292
rect 20322 3290 20346 3292
rect 20402 3290 20426 3292
rect 20482 3290 20488 3292
rect 20242 3238 20244 3290
rect 20424 3238 20426 3290
rect 20180 3236 20186 3238
rect 20242 3236 20266 3238
rect 20322 3236 20346 3238
rect 20402 3236 20426 3238
rect 20482 3236 20488 3238
rect 20180 3227 20488 3236
rect 20180 2204 20488 2213
rect 20180 2202 20186 2204
rect 20242 2202 20266 2204
rect 20322 2202 20346 2204
rect 20402 2202 20426 2204
rect 20482 2202 20488 2204
rect 20242 2150 20244 2202
rect 20424 2150 20426 2202
rect 20180 2148 20186 2150
rect 20242 2148 20266 2150
rect 20322 2148 20346 2150
rect 20402 2148 20426 2150
rect 20482 2148 20488 2150
rect 20180 2139 20488 2148
rect 21284 800 21312 6718
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6322 21404 6598
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 22572 5914 22600 6326
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22664 2774 22692 7958
rect 22848 6866 22876 9590
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22940 9178 22968 9454
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23032 9058 23060 9862
rect 23492 9654 23520 11086
rect 23860 11014 23888 11086
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10674 23888 10950
rect 23952 10810 23980 11222
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24320 10674 24348 11290
rect 25056 11218 25084 11290
rect 24860 11212 24912 11218
rect 25044 11212 25096 11218
rect 24912 11172 24992 11200
rect 24860 11154 24912 11160
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24676 11144 24728 11150
rect 24728 11092 24900 11098
rect 24676 11086 24900 11092
rect 24504 10810 24532 11086
rect 24688 11070 24900 11086
rect 24872 10810 24900 11070
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 9994 24624 10610
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 22940 9030 23060 9058
rect 22940 8906 22968 9030
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 22940 7274 22968 8842
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23400 8430 23428 8570
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 24228 7546 24256 9318
rect 24596 8634 24624 9930
rect 24780 9654 24808 10134
rect 24872 10062 24900 10746
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24964 9654 24992 11172
rect 25044 11154 25096 11160
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10810 25452 10950
rect 25412 10804 25464 10810
rect 25412 10746 25464 10752
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 24780 8634 24808 9590
rect 25332 9586 25360 10542
rect 25516 10266 25544 11154
rect 25976 10266 26004 12854
rect 26160 12850 26188 13194
rect 26436 12986 26464 13262
rect 27608 13084 27916 13093
rect 27608 13082 27614 13084
rect 27670 13082 27694 13084
rect 27750 13082 27774 13084
rect 27830 13082 27854 13084
rect 27910 13082 27916 13084
rect 27670 13030 27672 13082
rect 27852 13030 27854 13082
rect 27608 13028 27614 13030
rect 27670 13028 27694 13030
rect 27750 13028 27774 13030
rect 27830 13028 27854 13030
rect 27910 13028 27916 13030
rect 27608 13019 27916 13028
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26160 12434 26188 12786
rect 26948 12540 27256 12549
rect 26948 12538 26954 12540
rect 27010 12538 27034 12540
rect 27090 12538 27114 12540
rect 27170 12538 27194 12540
rect 27250 12538 27256 12540
rect 27010 12486 27012 12538
rect 27192 12486 27194 12538
rect 26948 12484 26954 12486
rect 27010 12484 27034 12486
rect 27090 12484 27114 12486
rect 27170 12484 27194 12486
rect 27250 12484 27256 12486
rect 26948 12475 27256 12484
rect 26068 12406 26188 12434
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 26068 10146 26096 12406
rect 27608 11996 27916 12005
rect 27608 11994 27614 11996
rect 27670 11994 27694 11996
rect 27750 11994 27774 11996
rect 27830 11994 27854 11996
rect 27910 11994 27916 11996
rect 27670 11942 27672 11994
rect 27852 11942 27854 11994
rect 27608 11940 27614 11942
rect 27670 11940 27694 11942
rect 27750 11940 27774 11942
rect 27830 11940 27854 11942
rect 27910 11940 27916 11942
rect 27608 11931 27916 11940
rect 26948 11452 27256 11461
rect 26948 11450 26954 11452
rect 27010 11450 27034 11452
rect 27090 11450 27114 11452
rect 27170 11450 27194 11452
rect 27250 11450 27256 11452
rect 27010 11398 27012 11450
rect 27192 11398 27194 11450
rect 26948 11396 26954 11398
rect 27010 11396 27034 11398
rect 27090 11396 27114 11398
rect 27170 11396 27194 11398
rect 27250 11396 27256 11398
rect 26948 11387 27256 11396
rect 27608 10908 27916 10917
rect 27608 10906 27614 10908
rect 27670 10906 27694 10908
rect 27750 10906 27774 10908
rect 27830 10906 27854 10908
rect 27910 10906 27916 10908
rect 27670 10854 27672 10906
rect 27852 10854 27854 10906
rect 27608 10852 27614 10854
rect 27670 10852 27694 10854
rect 27750 10852 27774 10854
rect 27830 10852 27854 10854
rect 27910 10852 27916 10854
rect 27608 10843 27916 10852
rect 26948 10364 27256 10373
rect 26948 10362 26954 10364
rect 27010 10362 27034 10364
rect 27090 10362 27114 10364
rect 27170 10362 27194 10364
rect 27250 10362 27256 10364
rect 27010 10310 27012 10362
rect 27192 10310 27194 10362
rect 26948 10308 26954 10310
rect 27010 10308 27034 10310
rect 27090 10308 27114 10310
rect 27170 10308 27194 10310
rect 27250 10308 27256 10310
rect 26948 10299 27256 10308
rect 25792 10130 26096 10146
rect 25780 10124 26096 10130
rect 25832 10118 26096 10124
rect 25780 10066 25832 10072
rect 25412 9988 25464 9994
rect 25412 9930 25464 9936
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25056 9178 25084 9522
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24584 8628 24636 8634
rect 24584 8570 24636 8576
rect 24768 8628 24820 8634
rect 24768 8570 24820 8576
rect 25148 8498 25176 8774
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 7886 24716 8298
rect 25332 8294 25360 9522
rect 25424 9110 25452 9930
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25412 9104 25464 9110
rect 25412 9046 25464 9052
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7546 24716 7822
rect 25424 7818 25452 8434
rect 25608 8022 25636 8570
rect 25700 8362 25728 9522
rect 25792 8974 25820 10066
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25976 9586 26004 9862
rect 27608 9820 27916 9829
rect 27608 9818 27614 9820
rect 27670 9818 27694 9820
rect 27750 9818 27774 9820
rect 27830 9818 27854 9820
rect 27910 9818 27916 9820
rect 27670 9766 27672 9818
rect 27852 9766 27854 9818
rect 27608 9764 27614 9766
rect 27670 9764 27694 9766
rect 27750 9764 27774 9766
rect 27830 9764 27854 9766
rect 27910 9764 27916 9766
rect 27608 9755 27916 9764
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 25884 8498 25912 8842
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25976 8090 26004 9522
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26160 9178 26188 9454
rect 26948 9276 27256 9285
rect 26948 9274 26954 9276
rect 27010 9274 27034 9276
rect 27090 9274 27114 9276
rect 27170 9274 27194 9276
rect 27250 9274 27256 9276
rect 27010 9222 27012 9274
rect 27192 9222 27194 9274
rect 26948 9220 26954 9222
rect 27010 9220 27034 9222
rect 27090 9220 27114 9222
rect 27170 9220 27194 9222
rect 27250 9220 27256 9222
rect 26948 9211 27256 9220
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 27608 8732 27916 8741
rect 27608 8730 27614 8732
rect 27670 8730 27694 8732
rect 27750 8730 27774 8732
rect 27830 8730 27854 8732
rect 27910 8730 27916 8732
rect 27670 8678 27672 8730
rect 27852 8678 27854 8730
rect 27608 8676 27614 8678
rect 27670 8676 27694 8678
rect 27750 8676 27774 8678
rect 27830 8676 27854 8678
rect 27910 8676 27916 8678
rect 27608 8667 27916 8676
rect 26948 8188 27256 8197
rect 26948 8186 26954 8188
rect 27010 8186 27034 8188
rect 27090 8186 27114 8188
rect 27170 8186 27194 8188
rect 27250 8186 27256 8188
rect 27010 8134 27012 8186
rect 27192 8134 27194 8186
rect 26948 8132 26954 8134
rect 27010 8132 27034 8134
rect 27090 8132 27114 8134
rect 27170 8132 27194 8134
rect 27250 8132 27256 8134
rect 26948 8123 27256 8132
rect 25964 8084 26016 8090
rect 25964 8026 26016 8032
rect 25596 8016 25648 8022
rect 25596 7958 25648 7964
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 25412 7812 25464 7818
rect 25412 7754 25464 7760
rect 25056 7546 25084 7754
rect 25608 7546 25636 7958
rect 27608 7644 27916 7653
rect 27608 7642 27614 7644
rect 27670 7642 27694 7644
rect 27750 7642 27774 7644
rect 27830 7642 27854 7644
rect 27910 7642 27916 7644
rect 27670 7590 27672 7642
rect 27852 7590 27854 7642
rect 27608 7588 27614 7590
rect 27670 7588 27694 7590
rect 27750 7588 27774 7590
rect 27830 7588 27854 7590
rect 27910 7588 27916 7590
rect 27608 7579 27916 7588
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 22928 7268 22980 7274
rect 22928 7210 22980 7216
rect 23032 6866 23060 7278
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 23676 6798 23704 7142
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23584 6186 23612 6598
rect 23860 6458 23888 6598
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 23572 6180 23624 6186
rect 23572 6122 23624 6128
rect 24412 5914 24440 6326
rect 24596 6254 24624 7346
rect 24688 6458 24716 7482
rect 26948 7100 27256 7109
rect 26948 7098 26954 7100
rect 27010 7098 27034 7100
rect 27090 7098 27114 7100
rect 27170 7098 27194 7100
rect 27250 7098 27256 7100
rect 27010 7046 27012 7098
rect 27192 7046 27194 7098
rect 26948 7044 26954 7046
rect 27010 7044 27034 7046
rect 27090 7044 27114 7046
rect 27170 7044 27194 7046
rect 27250 7044 27256 7046
rect 26948 7035 27256 7044
rect 27608 6556 27916 6565
rect 27608 6554 27614 6556
rect 27670 6554 27694 6556
rect 27750 6554 27774 6556
rect 27830 6554 27854 6556
rect 27910 6554 27916 6556
rect 27670 6502 27672 6554
rect 27852 6502 27854 6554
rect 27608 6500 27614 6502
rect 27670 6500 27694 6502
rect 27750 6500 27774 6502
rect 27830 6500 27854 6502
rect 27910 6500 27916 6502
rect 27608 6491 27916 6500
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 26948 6012 27256 6021
rect 26948 6010 26954 6012
rect 27010 6010 27034 6012
rect 27090 6010 27114 6012
rect 27170 6010 27194 6012
rect 27250 6010 27256 6012
rect 27010 5958 27012 6010
rect 27192 5958 27194 6010
rect 26948 5956 26954 5958
rect 27010 5956 27034 5958
rect 27090 5956 27114 5958
rect 27170 5956 27194 5958
rect 27250 5956 27256 5958
rect 26948 5947 27256 5956
rect 24400 5908 24452 5914
rect 24400 5850 24452 5856
rect 27608 5468 27916 5477
rect 27608 5466 27614 5468
rect 27670 5466 27694 5468
rect 27750 5466 27774 5468
rect 27830 5466 27854 5468
rect 27910 5466 27916 5468
rect 27670 5414 27672 5466
rect 27852 5414 27854 5466
rect 27608 5412 27614 5414
rect 27670 5412 27694 5414
rect 27750 5412 27774 5414
rect 27830 5412 27854 5414
rect 27910 5412 27916 5414
rect 27608 5403 27916 5412
rect 26948 4924 27256 4933
rect 26948 4922 26954 4924
rect 27010 4922 27034 4924
rect 27090 4922 27114 4924
rect 27170 4922 27194 4924
rect 27250 4922 27256 4924
rect 27010 4870 27012 4922
rect 27192 4870 27194 4922
rect 26948 4868 26954 4870
rect 27010 4868 27034 4870
rect 27090 4868 27114 4870
rect 27170 4868 27194 4870
rect 27250 4868 27256 4870
rect 26948 4859 27256 4868
rect 27608 4380 27916 4389
rect 27608 4378 27614 4380
rect 27670 4378 27694 4380
rect 27750 4378 27774 4380
rect 27830 4378 27854 4380
rect 27910 4378 27916 4380
rect 27670 4326 27672 4378
rect 27852 4326 27854 4378
rect 27608 4324 27614 4326
rect 27670 4324 27694 4326
rect 27750 4324 27774 4326
rect 27830 4324 27854 4326
rect 27910 4324 27916 4326
rect 27608 4315 27916 4324
rect 26948 3836 27256 3845
rect 26948 3834 26954 3836
rect 27010 3834 27034 3836
rect 27090 3834 27114 3836
rect 27170 3834 27194 3836
rect 27250 3834 27256 3836
rect 27010 3782 27012 3834
rect 27192 3782 27194 3834
rect 26948 3780 26954 3782
rect 27010 3780 27034 3782
rect 27090 3780 27114 3782
rect 27170 3780 27194 3782
rect 27250 3780 27256 3782
rect 26948 3771 27256 3780
rect 27608 3292 27916 3301
rect 27608 3290 27614 3292
rect 27670 3290 27694 3292
rect 27750 3290 27774 3292
rect 27830 3290 27854 3292
rect 27910 3290 27916 3292
rect 27670 3238 27672 3290
rect 27852 3238 27854 3290
rect 27608 3236 27614 3238
rect 27670 3236 27694 3238
rect 27750 3236 27774 3238
rect 27830 3236 27854 3238
rect 27910 3236 27916 3238
rect 27608 3227 27916 3236
rect 22572 2746 22692 2774
rect 26948 2748 27256 2757
rect 26948 2746 26954 2748
rect 27010 2746 27034 2748
rect 27090 2746 27114 2748
rect 27170 2746 27194 2748
rect 27250 2746 27256 2748
rect 22572 800 22600 2746
rect 27010 2694 27012 2746
rect 27192 2694 27194 2746
rect 26948 2692 26954 2694
rect 27010 2692 27034 2694
rect 27090 2692 27114 2694
rect 27170 2692 27194 2694
rect 27250 2692 27256 2694
rect 26948 2683 27256 2692
rect 27608 2204 27916 2213
rect 27608 2202 27614 2204
rect 27670 2202 27694 2204
rect 27750 2202 27774 2204
rect 27830 2202 27854 2204
rect 27910 2202 27916 2204
rect 27670 2150 27672 2202
rect 27852 2150 27854 2202
rect 27608 2148 27614 2150
rect 27670 2148 27694 2150
rect 27750 2148 27774 2150
rect 27830 2148 27854 2150
rect 27910 2148 27916 2150
rect 27608 2139 27916 2148
rect 11992 734 12204 762
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
<< via2 >>
rect 5330 29402 5386 29404
rect 5410 29402 5466 29404
rect 5490 29402 5546 29404
rect 5570 29402 5626 29404
rect 5330 29350 5376 29402
rect 5376 29350 5386 29402
rect 5410 29350 5440 29402
rect 5440 29350 5452 29402
rect 5452 29350 5466 29402
rect 5490 29350 5504 29402
rect 5504 29350 5516 29402
rect 5516 29350 5546 29402
rect 5570 29350 5580 29402
rect 5580 29350 5626 29402
rect 5330 29348 5386 29350
rect 5410 29348 5466 29350
rect 5490 29348 5546 29350
rect 5570 29348 5626 29350
rect 12758 29402 12814 29404
rect 12838 29402 12894 29404
rect 12918 29402 12974 29404
rect 12998 29402 13054 29404
rect 12758 29350 12804 29402
rect 12804 29350 12814 29402
rect 12838 29350 12868 29402
rect 12868 29350 12880 29402
rect 12880 29350 12894 29402
rect 12918 29350 12932 29402
rect 12932 29350 12944 29402
rect 12944 29350 12974 29402
rect 12998 29350 13008 29402
rect 13008 29350 13054 29402
rect 12758 29348 12814 29350
rect 12838 29348 12894 29350
rect 12918 29348 12974 29350
rect 12998 29348 13054 29350
rect 4670 28858 4726 28860
rect 4750 28858 4806 28860
rect 4830 28858 4886 28860
rect 4910 28858 4966 28860
rect 4670 28806 4716 28858
rect 4716 28806 4726 28858
rect 4750 28806 4780 28858
rect 4780 28806 4792 28858
rect 4792 28806 4806 28858
rect 4830 28806 4844 28858
rect 4844 28806 4856 28858
rect 4856 28806 4886 28858
rect 4910 28806 4920 28858
rect 4920 28806 4966 28858
rect 4670 28804 4726 28806
rect 4750 28804 4806 28806
rect 4830 28804 4886 28806
rect 4910 28804 4966 28806
rect 12098 28858 12154 28860
rect 12178 28858 12234 28860
rect 12258 28858 12314 28860
rect 12338 28858 12394 28860
rect 12098 28806 12144 28858
rect 12144 28806 12154 28858
rect 12178 28806 12208 28858
rect 12208 28806 12220 28858
rect 12220 28806 12234 28858
rect 12258 28806 12272 28858
rect 12272 28806 12284 28858
rect 12284 28806 12314 28858
rect 12338 28806 12348 28858
rect 12348 28806 12394 28858
rect 12098 28804 12154 28806
rect 12178 28804 12234 28806
rect 12258 28804 12314 28806
rect 12338 28804 12394 28806
rect 5330 28314 5386 28316
rect 5410 28314 5466 28316
rect 5490 28314 5546 28316
rect 5570 28314 5626 28316
rect 5330 28262 5376 28314
rect 5376 28262 5386 28314
rect 5410 28262 5440 28314
rect 5440 28262 5452 28314
rect 5452 28262 5466 28314
rect 5490 28262 5504 28314
rect 5504 28262 5516 28314
rect 5516 28262 5546 28314
rect 5570 28262 5580 28314
rect 5580 28262 5626 28314
rect 5330 28260 5386 28262
rect 5410 28260 5466 28262
rect 5490 28260 5546 28262
rect 5570 28260 5626 28262
rect 12758 28314 12814 28316
rect 12838 28314 12894 28316
rect 12918 28314 12974 28316
rect 12998 28314 13054 28316
rect 12758 28262 12804 28314
rect 12804 28262 12814 28314
rect 12838 28262 12868 28314
rect 12868 28262 12880 28314
rect 12880 28262 12894 28314
rect 12918 28262 12932 28314
rect 12932 28262 12944 28314
rect 12944 28262 12974 28314
rect 12998 28262 13008 28314
rect 13008 28262 13054 28314
rect 12758 28260 12814 28262
rect 12838 28260 12894 28262
rect 12918 28260 12974 28262
rect 12998 28260 13054 28262
rect 4670 27770 4726 27772
rect 4750 27770 4806 27772
rect 4830 27770 4886 27772
rect 4910 27770 4966 27772
rect 4670 27718 4716 27770
rect 4716 27718 4726 27770
rect 4750 27718 4780 27770
rect 4780 27718 4792 27770
rect 4792 27718 4806 27770
rect 4830 27718 4844 27770
rect 4844 27718 4856 27770
rect 4856 27718 4886 27770
rect 4910 27718 4920 27770
rect 4920 27718 4966 27770
rect 4670 27716 4726 27718
rect 4750 27716 4806 27718
rect 4830 27716 4886 27718
rect 4910 27716 4966 27718
rect 12098 27770 12154 27772
rect 12178 27770 12234 27772
rect 12258 27770 12314 27772
rect 12338 27770 12394 27772
rect 12098 27718 12144 27770
rect 12144 27718 12154 27770
rect 12178 27718 12208 27770
rect 12208 27718 12220 27770
rect 12220 27718 12234 27770
rect 12258 27718 12272 27770
rect 12272 27718 12284 27770
rect 12284 27718 12314 27770
rect 12338 27718 12348 27770
rect 12348 27718 12394 27770
rect 12098 27716 12154 27718
rect 12178 27716 12234 27718
rect 12258 27716 12314 27718
rect 12338 27716 12394 27718
rect 5330 27226 5386 27228
rect 5410 27226 5466 27228
rect 5490 27226 5546 27228
rect 5570 27226 5626 27228
rect 5330 27174 5376 27226
rect 5376 27174 5386 27226
rect 5410 27174 5440 27226
rect 5440 27174 5452 27226
rect 5452 27174 5466 27226
rect 5490 27174 5504 27226
rect 5504 27174 5516 27226
rect 5516 27174 5546 27226
rect 5570 27174 5580 27226
rect 5580 27174 5626 27226
rect 5330 27172 5386 27174
rect 5410 27172 5466 27174
rect 5490 27172 5546 27174
rect 5570 27172 5626 27174
rect 12758 27226 12814 27228
rect 12838 27226 12894 27228
rect 12918 27226 12974 27228
rect 12998 27226 13054 27228
rect 12758 27174 12804 27226
rect 12804 27174 12814 27226
rect 12838 27174 12868 27226
rect 12868 27174 12880 27226
rect 12880 27174 12894 27226
rect 12918 27174 12932 27226
rect 12932 27174 12944 27226
rect 12944 27174 12974 27226
rect 12998 27174 13008 27226
rect 13008 27174 13054 27226
rect 12758 27172 12814 27174
rect 12838 27172 12894 27174
rect 12918 27172 12974 27174
rect 12998 27172 13054 27174
rect 4670 26682 4726 26684
rect 4750 26682 4806 26684
rect 4830 26682 4886 26684
rect 4910 26682 4966 26684
rect 4670 26630 4716 26682
rect 4716 26630 4726 26682
rect 4750 26630 4780 26682
rect 4780 26630 4792 26682
rect 4792 26630 4806 26682
rect 4830 26630 4844 26682
rect 4844 26630 4856 26682
rect 4856 26630 4886 26682
rect 4910 26630 4920 26682
rect 4920 26630 4966 26682
rect 4670 26628 4726 26630
rect 4750 26628 4806 26630
rect 4830 26628 4886 26630
rect 4910 26628 4966 26630
rect 12098 26682 12154 26684
rect 12178 26682 12234 26684
rect 12258 26682 12314 26684
rect 12338 26682 12394 26684
rect 12098 26630 12144 26682
rect 12144 26630 12154 26682
rect 12178 26630 12208 26682
rect 12208 26630 12220 26682
rect 12220 26630 12234 26682
rect 12258 26630 12272 26682
rect 12272 26630 12284 26682
rect 12284 26630 12314 26682
rect 12338 26630 12348 26682
rect 12348 26630 12394 26682
rect 12098 26628 12154 26630
rect 12178 26628 12234 26630
rect 12258 26628 12314 26630
rect 12338 26628 12394 26630
rect 5330 26138 5386 26140
rect 5410 26138 5466 26140
rect 5490 26138 5546 26140
rect 5570 26138 5626 26140
rect 5330 26086 5376 26138
rect 5376 26086 5386 26138
rect 5410 26086 5440 26138
rect 5440 26086 5452 26138
rect 5452 26086 5466 26138
rect 5490 26086 5504 26138
rect 5504 26086 5516 26138
rect 5516 26086 5546 26138
rect 5570 26086 5580 26138
rect 5580 26086 5626 26138
rect 5330 26084 5386 26086
rect 5410 26084 5466 26086
rect 5490 26084 5546 26086
rect 5570 26084 5626 26086
rect 12758 26138 12814 26140
rect 12838 26138 12894 26140
rect 12918 26138 12974 26140
rect 12998 26138 13054 26140
rect 12758 26086 12804 26138
rect 12804 26086 12814 26138
rect 12838 26086 12868 26138
rect 12868 26086 12880 26138
rect 12880 26086 12894 26138
rect 12918 26086 12932 26138
rect 12932 26086 12944 26138
rect 12944 26086 12974 26138
rect 12998 26086 13008 26138
rect 13008 26086 13054 26138
rect 12758 26084 12814 26086
rect 12838 26084 12894 26086
rect 12918 26084 12974 26086
rect 12998 26084 13054 26086
rect 3974 25880 4030 25936
rect 938 21120 994 21176
rect 1490 20576 1546 20632
rect 938 19760 994 19816
rect 1490 19116 1492 19136
rect 1492 19116 1544 19136
rect 1544 19116 1546 19136
rect 1490 19080 1546 19116
rect 938 18400 994 18456
rect 4670 25594 4726 25596
rect 4750 25594 4806 25596
rect 4830 25594 4886 25596
rect 4910 25594 4966 25596
rect 4670 25542 4716 25594
rect 4716 25542 4726 25594
rect 4750 25542 4780 25594
rect 4780 25542 4792 25594
rect 4792 25542 4806 25594
rect 4830 25542 4844 25594
rect 4844 25542 4856 25594
rect 4856 25542 4886 25594
rect 4910 25542 4920 25594
rect 4920 25542 4966 25594
rect 4670 25540 4726 25542
rect 4750 25540 4806 25542
rect 4830 25540 4886 25542
rect 4910 25540 4966 25542
rect 12098 25594 12154 25596
rect 12178 25594 12234 25596
rect 12258 25594 12314 25596
rect 12338 25594 12394 25596
rect 12098 25542 12144 25594
rect 12144 25542 12154 25594
rect 12178 25542 12208 25594
rect 12208 25542 12220 25594
rect 12220 25542 12234 25594
rect 12258 25542 12272 25594
rect 12272 25542 12284 25594
rect 12284 25542 12314 25594
rect 12338 25542 12348 25594
rect 12348 25542 12394 25594
rect 12098 25540 12154 25542
rect 12178 25540 12234 25542
rect 12258 25540 12314 25542
rect 12338 25540 12394 25542
rect 5330 25050 5386 25052
rect 5410 25050 5466 25052
rect 5490 25050 5546 25052
rect 5570 25050 5626 25052
rect 5330 24998 5376 25050
rect 5376 24998 5386 25050
rect 5410 24998 5440 25050
rect 5440 24998 5452 25050
rect 5452 24998 5466 25050
rect 5490 24998 5504 25050
rect 5504 24998 5516 25050
rect 5516 24998 5546 25050
rect 5570 24998 5580 25050
rect 5580 24998 5626 25050
rect 5330 24996 5386 24998
rect 5410 24996 5466 24998
rect 5490 24996 5546 24998
rect 5570 24996 5626 24998
rect 4670 24506 4726 24508
rect 4750 24506 4806 24508
rect 4830 24506 4886 24508
rect 4910 24506 4966 24508
rect 4670 24454 4716 24506
rect 4716 24454 4726 24506
rect 4750 24454 4780 24506
rect 4780 24454 4792 24506
rect 4792 24454 4806 24506
rect 4830 24454 4844 24506
rect 4844 24454 4856 24506
rect 4856 24454 4886 24506
rect 4910 24454 4920 24506
rect 4920 24454 4966 24506
rect 4670 24452 4726 24454
rect 4750 24452 4806 24454
rect 4830 24452 4886 24454
rect 4910 24452 4966 24454
rect 12758 25050 12814 25052
rect 12838 25050 12894 25052
rect 12918 25050 12974 25052
rect 12998 25050 13054 25052
rect 12758 24998 12804 25050
rect 12804 24998 12814 25050
rect 12838 24998 12868 25050
rect 12868 24998 12880 25050
rect 12880 24998 12894 25050
rect 12918 24998 12932 25050
rect 12932 24998 12944 25050
rect 12944 24998 12974 25050
rect 12998 24998 13008 25050
rect 13008 24998 13054 25050
rect 12758 24996 12814 24998
rect 12838 24996 12894 24998
rect 12918 24996 12974 24998
rect 12998 24996 13054 24998
rect 5330 23962 5386 23964
rect 5410 23962 5466 23964
rect 5490 23962 5546 23964
rect 5570 23962 5626 23964
rect 5330 23910 5376 23962
rect 5376 23910 5386 23962
rect 5410 23910 5440 23962
rect 5440 23910 5452 23962
rect 5452 23910 5466 23962
rect 5490 23910 5504 23962
rect 5504 23910 5516 23962
rect 5516 23910 5546 23962
rect 5570 23910 5580 23962
rect 5580 23910 5626 23962
rect 5330 23908 5386 23910
rect 5410 23908 5466 23910
rect 5490 23908 5546 23910
rect 5570 23908 5626 23910
rect 4670 23418 4726 23420
rect 4750 23418 4806 23420
rect 4830 23418 4886 23420
rect 4910 23418 4966 23420
rect 4670 23366 4716 23418
rect 4716 23366 4726 23418
rect 4750 23366 4780 23418
rect 4780 23366 4792 23418
rect 4792 23366 4806 23418
rect 4830 23366 4844 23418
rect 4844 23366 4856 23418
rect 4856 23366 4886 23418
rect 4910 23366 4920 23418
rect 4920 23366 4966 23418
rect 4670 23364 4726 23366
rect 4750 23364 4806 23366
rect 4830 23364 4886 23366
rect 4910 23364 4966 23366
rect 5330 22874 5386 22876
rect 5410 22874 5466 22876
rect 5490 22874 5546 22876
rect 5570 22874 5626 22876
rect 5330 22822 5376 22874
rect 5376 22822 5386 22874
rect 5410 22822 5440 22874
rect 5440 22822 5452 22874
rect 5452 22822 5466 22874
rect 5490 22822 5504 22874
rect 5504 22822 5516 22874
rect 5516 22822 5546 22874
rect 5570 22822 5580 22874
rect 5580 22822 5626 22874
rect 5330 22820 5386 22822
rect 5410 22820 5466 22822
rect 5490 22820 5546 22822
rect 5570 22820 5626 22822
rect 4670 22330 4726 22332
rect 4750 22330 4806 22332
rect 4830 22330 4886 22332
rect 4910 22330 4966 22332
rect 4670 22278 4716 22330
rect 4716 22278 4726 22330
rect 4750 22278 4780 22330
rect 4780 22278 4792 22330
rect 4792 22278 4806 22330
rect 4830 22278 4844 22330
rect 4844 22278 4856 22330
rect 4856 22278 4886 22330
rect 4910 22278 4920 22330
rect 4920 22278 4966 22330
rect 4670 22276 4726 22278
rect 4750 22276 4806 22278
rect 4830 22276 4886 22278
rect 4910 22276 4966 22278
rect 938 14320 994 14376
rect 4066 15000 4122 15056
rect 4066 13676 4068 13696
rect 4068 13676 4120 13696
rect 4120 13676 4122 13696
rect 4066 13640 4122 13676
rect 4670 21242 4726 21244
rect 4750 21242 4806 21244
rect 4830 21242 4886 21244
rect 4910 21242 4966 21244
rect 4670 21190 4716 21242
rect 4716 21190 4726 21242
rect 4750 21190 4780 21242
rect 4780 21190 4792 21242
rect 4792 21190 4806 21242
rect 4830 21190 4844 21242
rect 4844 21190 4856 21242
rect 4856 21190 4886 21242
rect 4910 21190 4920 21242
rect 4920 21190 4966 21242
rect 4670 21188 4726 21190
rect 4750 21188 4806 21190
rect 4830 21188 4886 21190
rect 4910 21188 4966 21190
rect 4670 20154 4726 20156
rect 4750 20154 4806 20156
rect 4830 20154 4886 20156
rect 4910 20154 4966 20156
rect 4670 20102 4716 20154
rect 4716 20102 4726 20154
rect 4750 20102 4780 20154
rect 4780 20102 4792 20154
rect 4792 20102 4806 20154
rect 4830 20102 4844 20154
rect 4844 20102 4856 20154
rect 4856 20102 4886 20154
rect 4910 20102 4920 20154
rect 4920 20102 4966 20154
rect 4670 20100 4726 20102
rect 4750 20100 4806 20102
rect 4830 20100 4886 20102
rect 4910 20100 4966 20102
rect 5330 21786 5386 21788
rect 5410 21786 5466 21788
rect 5490 21786 5546 21788
rect 5570 21786 5626 21788
rect 5330 21734 5376 21786
rect 5376 21734 5386 21786
rect 5410 21734 5440 21786
rect 5440 21734 5452 21786
rect 5452 21734 5466 21786
rect 5490 21734 5504 21786
rect 5504 21734 5516 21786
rect 5516 21734 5546 21786
rect 5570 21734 5580 21786
rect 5580 21734 5626 21786
rect 5330 21732 5386 21734
rect 5410 21732 5466 21734
rect 5490 21732 5546 21734
rect 5570 21732 5626 21734
rect 5330 20698 5386 20700
rect 5410 20698 5466 20700
rect 5490 20698 5546 20700
rect 5570 20698 5626 20700
rect 5330 20646 5376 20698
rect 5376 20646 5386 20698
rect 5410 20646 5440 20698
rect 5440 20646 5452 20698
rect 5452 20646 5466 20698
rect 5490 20646 5504 20698
rect 5504 20646 5516 20698
rect 5516 20646 5546 20698
rect 5570 20646 5580 20698
rect 5580 20646 5626 20698
rect 5330 20644 5386 20646
rect 5410 20644 5466 20646
rect 5490 20644 5546 20646
rect 5570 20644 5626 20646
rect 4670 19066 4726 19068
rect 4750 19066 4806 19068
rect 4830 19066 4886 19068
rect 4910 19066 4966 19068
rect 4670 19014 4716 19066
rect 4716 19014 4726 19066
rect 4750 19014 4780 19066
rect 4780 19014 4792 19066
rect 4792 19014 4806 19066
rect 4830 19014 4844 19066
rect 4844 19014 4856 19066
rect 4856 19014 4886 19066
rect 4910 19014 4920 19066
rect 4920 19014 4966 19066
rect 4670 19012 4726 19014
rect 4750 19012 4806 19014
rect 4830 19012 4886 19014
rect 4910 19012 4966 19014
rect 5330 19610 5386 19612
rect 5410 19610 5466 19612
rect 5490 19610 5546 19612
rect 5570 19610 5626 19612
rect 5330 19558 5376 19610
rect 5376 19558 5386 19610
rect 5410 19558 5440 19610
rect 5440 19558 5452 19610
rect 5452 19558 5466 19610
rect 5490 19558 5504 19610
rect 5504 19558 5516 19610
rect 5516 19558 5546 19610
rect 5570 19558 5580 19610
rect 5580 19558 5626 19610
rect 5330 19556 5386 19558
rect 5410 19556 5466 19558
rect 5490 19556 5546 19558
rect 5570 19556 5626 19558
rect 5330 18522 5386 18524
rect 5410 18522 5466 18524
rect 5490 18522 5546 18524
rect 5570 18522 5626 18524
rect 5330 18470 5376 18522
rect 5376 18470 5386 18522
rect 5410 18470 5440 18522
rect 5440 18470 5452 18522
rect 5452 18470 5466 18522
rect 5490 18470 5504 18522
rect 5504 18470 5516 18522
rect 5516 18470 5546 18522
rect 5570 18470 5580 18522
rect 5580 18470 5626 18522
rect 5330 18468 5386 18470
rect 5410 18468 5466 18470
rect 5490 18468 5546 18470
rect 5570 18468 5626 18470
rect 4670 17978 4726 17980
rect 4750 17978 4806 17980
rect 4830 17978 4886 17980
rect 4910 17978 4966 17980
rect 4670 17926 4716 17978
rect 4716 17926 4726 17978
rect 4750 17926 4780 17978
rect 4780 17926 4792 17978
rect 4792 17926 4806 17978
rect 4830 17926 4844 17978
rect 4844 17926 4856 17978
rect 4856 17926 4886 17978
rect 4910 17926 4920 17978
rect 4920 17926 4966 17978
rect 4670 17924 4726 17926
rect 4750 17924 4806 17926
rect 4830 17924 4886 17926
rect 4910 17924 4966 17926
rect 4670 16890 4726 16892
rect 4750 16890 4806 16892
rect 4830 16890 4886 16892
rect 4910 16890 4966 16892
rect 4670 16838 4716 16890
rect 4716 16838 4726 16890
rect 4750 16838 4780 16890
rect 4780 16838 4792 16890
rect 4792 16838 4806 16890
rect 4830 16838 4844 16890
rect 4844 16838 4856 16890
rect 4856 16838 4886 16890
rect 4910 16838 4920 16890
rect 4920 16838 4966 16890
rect 4670 16836 4726 16838
rect 4750 16836 4806 16838
rect 4830 16836 4886 16838
rect 4910 16836 4966 16838
rect 4434 16360 4490 16416
rect 4342 15680 4398 15736
rect 5330 17434 5386 17436
rect 5410 17434 5466 17436
rect 5490 17434 5546 17436
rect 5570 17434 5626 17436
rect 5330 17382 5376 17434
rect 5376 17382 5386 17434
rect 5410 17382 5440 17434
rect 5440 17382 5452 17434
rect 5452 17382 5466 17434
rect 5490 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5546 17434
rect 5570 17382 5580 17434
rect 5580 17382 5626 17434
rect 5330 17380 5386 17382
rect 5410 17380 5466 17382
rect 5490 17380 5546 17382
rect 5570 17380 5626 17382
rect 5330 16346 5386 16348
rect 5410 16346 5466 16348
rect 5490 16346 5546 16348
rect 5570 16346 5626 16348
rect 5330 16294 5376 16346
rect 5376 16294 5386 16346
rect 5410 16294 5440 16346
rect 5440 16294 5452 16346
rect 5452 16294 5466 16346
rect 5490 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5546 16346
rect 5570 16294 5580 16346
rect 5580 16294 5626 16346
rect 5330 16292 5386 16294
rect 5410 16292 5466 16294
rect 5490 16292 5546 16294
rect 5570 16292 5626 16294
rect 4670 15802 4726 15804
rect 4750 15802 4806 15804
rect 4830 15802 4886 15804
rect 4910 15802 4966 15804
rect 4670 15750 4716 15802
rect 4716 15750 4726 15802
rect 4750 15750 4780 15802
rect 4780 15750 4792 15802
rect 4792 15750 4806 15802
rect 4830 15750 4844 15802
rect 4844 15750 4856 15802
rect 4856 15750 4886 15802
rect 4910 15750 4920 15802
rect 4920 15750 4966 15802
rect 4670 15748 4726 15750
rect 4750 15748 4806 15750
rect 4830 15748 4886 15750
rect 4910 15748 4966 15750
rect 7930 17040 7986 17096
rect 5330 15258 5386 15260
rect 5410 15258 5466 15260
rect 5490 15258 5546 15260
rect 5570 15258 5626 15260
rect 5330 15206 5376 15258
rect 5376 15206 5386 15258
rect 5410 15206 5440 15258
rect 5440 15206 5452 15258
rect 5452 15206 5466 15258
rect 5490 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5546 15258
rect 5570 15206 5580 15258
rect 5580 15206 5626 15258
rect 5330 15204 5386 15206
rect 5410 15204 5466 15206
rect 5490 15204 5546 15206
rect 5570 15204 5626 15206
rect 4670 14714 4726 14716
rect 4750 14714 4806 14716
rect 4830 14714 4886 14716
rect 4910 14714 4966 14716
rect 4670 14662 4716 14714
rect 4716 14662 4726 14714
rect 4750 14662 4780 14714
rect 4780 14662 4792 14714
rect 4792 14662 4806 14714
rect 4830 14662 4844 14714
rect 4844 14662 4856 14714
rect 4856 14662 4886 14714
rect 4910 14662 4920 14714
rect 4920 14662 4966 14714
rect 4670 14660 4726 14662
rect 4750 14660 4806 14662
rect 4830 14660 4886 14662
rect 4910 14660 4966 14662
rect 4670 13626 4726 13628
rect 4750 13626 4806 13628
rect 4830 13626 4886 13628
rect 4910 13626 4966 13628
rect 4670 13574 4716 13626
rect 4716 13574 4726 13626
rect 4750 13574 4780 13626
rect 4780 13574 4792 13626
rect 4792 13574 4806 13626
rect 4830 13574 4844 13626
rect 4844 13574 4856 13626
rect 4856 13574 4886 13626
rect 4910 13574 4920 13626
rect 4920 13574 4966 13626
rect 4670 13572 4726 13574
rect 4750 13572 4806 13574
rect 4830 13572 4886 13574
rect 4910 13572 4966 13574
rect 5330 14170 5386 14172
rect 5410 14170 5466 14172
rect 5490 14170 5546 14172
rect 5570 14170 5626 14172
rect 5330 14118 5376 14170
rect 5376 14118 5386 14170
rect 5410 14118 5440 14170
rect 5440 14118 5452 14170
rect 5452 14118 5466 14170
rect 5490 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5546 14170
rect 5570 14118 5580 14170
rect 5580 14118 5626 14170
rect 5330 14116 5386 14118
rect 5410 14116 5466 14118
rect 5490 14116 5546 14118
rect 5570 14116 5626 14118
rect 5330 13082 5386 13084
rect 5410 13082 5466 13084
rect 5490 13082 5546 13084
rect 5570 13082 5626 13084
rect 5330 13030 5376 13082
rect 5376 13030 5386 13082
rect 5410 13030 5440 13082
rect 5440 13030 5452 13082
rect 5452 13030 5466 13082
rect 5490 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5546 13082
rect 5570 13030 5580 13082
rect 5580 13030 5626 13082
rect 5330 13028 5386 13030
rect 5410 13028 5466 13030
rect 5490 13028 5546 13030
rect 5570 13028 5626 13030
rect 3974 12300 4030 12336
rect 3974 12280 3976 12300
rect 3976 12280 4028 12300
rect 4028 12280 4030 12300
rect 3974 10920 4030 10976
rect 4066 9596 4068 9616
rect 4068 9596 4120 9616
rect 4120 9596 4122 9616
rect 4066 9560 4122 9596
rect 4670 12538 4726 12540
rect 4750 12538 4806 12540
rect 4830 12538 4886 12540
rect 4910 12538 4966 12540
rect 4670 12486 4716 12538
rect 4716 12486 4726 12538
rect 4750 12486 4780 12538
rect 4780 12486 4792 12538
rect 4792 12486 4806 12538
rect 4830 12486 4844 12538
rect 4844 12486 4856 12538
rect 4856 12486 4886 12538
rect 4910 12486 4920 12538
rect 4920 12486 4966 12538
rect 4670 12484 4726 12486
rect 4750 12484 4806 12486
rect 4830 12484 4886 12486
rect 4910 12484 4966 12486
rect 4670 11450 4726 11452
rect 4750 11450 4806 11452
rect 4830 11450 4886 11452
rect 4910 11450 4966 11452
rect 4670 11398 4716 11450
rect 4716 11398 4726 11450
rect 4750 11398 4780 11450
rect 4780 11398 4792 11450
rect 4792 11398 4806 11450
rect 4830 11398 4844 11450
rect 4844 11398 4856 11450
rect 4856 11398 4886 11450
rect 4910 11398 4920 11450
rect 4920 11398 4966 11450
rect 4670 11396 4726 11398
rect 4750 11396 4806 11398
rect 4830 11396 4886 11398
rect 4910 11396 4966 11398
rect 5330 11994 5386 11996
rect 5410 11994 5466 11996
rect 5490 11994 5546 11996
rect 5570 11994 5626 11996
rect 5330 11942 5376 11994
rect 5376 11942 5386 11994
rect 5410 11942 5440 11994
rect 5440 11942 5452 11994
rect 5452 11942 5466 11994
rect 5490 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5546 11994
rect 5570 11942 5580 11994
rect 5580 11942 5626 11994
rect 5330 11940 5386 11942
rect 5410 11940 5466 11942
rect 5490 11940 5546 11942
rect 5570 11940 5626 11942
rect 4670 10362 4726 10364
rect 4750 10362 4806 10364
rect 4830 10362 4886 10364
rect 4910 10362 4966 10364
rect 4670 10310 4716 10362
rect 4716 10310 4726 10362
rect 4750 10310 4780 10362
rect 4780 10310 4792 10362
rect 4792 10310 4806 10362
rect 4830 10310 4844 10362
rect 4844 10310 4856 10362
rect 4856 10310 4886 10362
rect 4910 10310 4920 10362
rect 4920 10310 4966 10362
rect 4670 10308 4726 10310
rect 4750 10308 4806 10310
rect 4830 10308 4886 10310
rect 4910 10308 4966 10310
rect 4670 9274 4726 9276
rect 4750 9274 4806 9276
rect 4830 9274 4886 9276
rect 4910 9274 4966 9276
rect 4670 9222 4716 9274
rect 4716 9222 4726 9274
rect 4750 9222 4780 9274
rect 4780 9222 4792 9274
rect 4792 9222 4806 9274
rect 4830 9222 4844 9274
rect 4844 9222 4856 9274
rect 4856 9222 4886 9274
rect 4910 9222 4920 9274
rect 4920 9222 4966 9274
rect 4670 9220 4726 9222
rect 4750 9220 4806 9222
rect 4830 9220 4886 9222
rect 4910 9220 4966 9222
rect 5330 10906 5386 10908
rect 5410 10906 5466 10908
rect 5490 10906 5546 10908
rect 5570 10906 5626 10908
rect 5330 10854 5376 10906
rect 5376 10854 5386 10906
rect 5410 10854 5440 10906
rect 5440 10854 5452 10906
rect 5452 10854 5466 10906
rect 5490 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5546 10906
rect 5570 10854 5580 10906
rect 5580 10854 5626 10906
rect 5330 10852 5386 10854
rect 5410 10852 5466 10854
rect 5490 10852 5546 10854
rect 5570 10852 5626 10854
rect 5330 9818 5386 9820
rect 5410 9818 5466 9820
rect 5490 9818 5546 9820
rect 5570 9818 5626 9820
rect 5330 9766 5376 9818
rect 5376 9766 5386 9818
rect 5410 9766 5440 9818
rect 5440 9766 5452 9818
rect 5452 9766 5466 9818
rect 5490 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5546 9818
rect 5570 9766 5580 9818
rect 5580 9766 5626 9818
rect 5330 9764 5386 9766
rect 5410 9764 5466 9766
rect 5490 9764 5546 9766
rect 5570 9764 5626 9766
rect 4066 8200 4122 8256
rect 4670 8186 4726 8188
rect 4750 8186 4806 8188
rect 4830 8186 4886 8188
rect 4910 8186 4966 8188
rect 4670 8134 4716 8186
rect 4716 8134 4726 8186
rect 4750 8134 4780 8186
rect 4780 8134 4792 8186
rect 4792 8134 4806 8186
rect 4830 8134 4844 8186
rect 4844 8134 4856 8186
rect 4856 8134 4886 8186
rect 4910 8134 4920 8186
rect 4920 8134 4966 8186
rect 4670 8132 4726 8134
rect 4750 8132 4806 8134
rect 4830 8132 4886 8134
rect 4910 8132 4966 8134
rect 5330 8730 5386 8732
rect 5410 8730 5466 8732
rect 5490 8730 5546 8732
rect 5570 8730 5626 8732
rect 5330 8678 5376 8730
rect 5376 8678 5386 8730
rect 5410 8678 5440 8730
rect 5440 8678 5452 8730
rect 5452 8678 5466 8730
rect 5490 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5546 8730
rect 5570 8678 5580 8730
rect 5580 8678 5626 8730
rect 5330 8676 5386 8678
rect 5410 8676 5466 8678
rect 5490 8676 5546 8678
rect 5570 8676 5626 8678
rect 4670 7098 4726 7100
rect 4750 7098 4806 7100
rect 4830 7098 4886 7100
rect 4910 7098 4966 7100
rect 4670 7046 4716 7098
rect 4716 7046 4726 7098
rect 4750 7046 4780 7098
rect 4780 7046 4792 7098
rect 4792 7046 4806 7098
rect 4830 7046 4844 7098
rect 4844 7046 4856 7098
rect 4856 7046 4886 7098
rect 4910 7046 4920 7098
rect 4920 7046 4966 7098
rect 4670 7044 4726 7046
rect 4750 7044 4806 7046
rect 4830 7044 4886 7046
rect 4910 7044 4966 7046
rect 5330 7642 5386 7644
rect 5410 7642 5466 7644
rect 5490 7642 5546 7644
rect 5570 7642 5626 7644
rect 5330 7590 5376 7642
rect 5376 7590 5386 7642
rect 5410 7590 5440 7642
rect 5440 7590 5452 7642
rect 5452 7590 5466 7642
rect 5490 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5546 7642
rect 5570 7590 5580 7642
rect 5580 7590 5626 7642
rect 5330 7588 5386 7590
rect 5410 7588 5466 7590
rect 5490 7588 5546 7590
rect 5570 7588 5626 7590
rect 5330 6554 5386 6556
rect 5410 6554 5466 6556
rect 5490 6554 5546 6556
rect 5570 6554 5626 6556
rect 5330 6502 5376 6554
rect 5376 6502 5386 6554
rect 5410 6502 5440 6554
rect 5440 6502 5452 6554
rect 5452 6502 5466 6554
rect 5490 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5546 6554
rect 5570 6502 5580 6554
rect 5580 6502 5626 6554
rect 5330 6500 5386 6502
rect 5410 6500 5466 6502
rect 5490 6500 5546 6502
rect 5570 6500 5626 6502
rect 4670 6010 4726 6012
rect 4750 6010 4806 6012
rect 4830 6010 4886 6012
rect 4910 6010 4966 6012
rect 4670 5958 4716 6010
rect 4716 5958 4726 6010
rect 4750 5958 4780 6010
rect 4780 5958 4792 6010
rect 4792 5958 4806 6010
rect 4830 5958 4844 6010
rect 4844 5958 4856 6010
rect 4856 5958 4886 6010
rect 4910 5958 4920 6010
rect 4920 5958 4966 6010
rect 4670 5956 4726 5958
rect 4750 5956 4806 5958
rect 4830 5956 4886 5958
rect 4910 5956 4966 5958
rect 8666 13812 8668 13832
rect 8668 13812 8720 13832
rect 8720 13812 8722 13832
rect 8666 13776 8722 13812
rect 12098 24506 12154 24508
rect 12178 24506 12234 24508
rect 12258 24506 12314 24508
rect 12338 24506 12394 24508
rect 12098 24454 12144 24506
rect 12144 24454 12154 24506
rect 12178 24454 12208 24506
rect 12208 24454 12220 24506
rect 12220 24454 12234 24506
rect 12258 24454 12272 24506
rect 12272 24454 12284 24506
rect 12284 24454 12314 24506
rect 12338 24454 12348 24506
rect 12348 24454 12394 24506
rect 12098 24452 12154 24454
rect 12178 24452 12234 24454
rect 12258 24452 12314 24454
rect 12338 24452 12394 24454
rect 12758 23962 12814 23964
rect 12838 23962 12894 23964
rect 12918 23962 12974 23964
rect 12998 23962 13054 23964
rect 12758 23910 12804 23962
rect 12804 23910 12814 23962
rect 12838 23910 12868 23962
rect 12868 23910 12880 23962
rect 12880 23910 12894 23962
rect 12918 23910 12932 23962
rect 12932 23910 12944 23962
rect 12944 23910 12974 23962
rect 12998 23910 13008 23962
rect 13008 23910 13054 23962
rect 12758 23908 12814 23910
rect 12838 23908 12894 23910
rect 12918 23908 12974 23910
rect 12998 23908 13054 23910
rect 12098 23418 12154 23420
rect 12178 23418 12234 23420
rect 12258 23418 12314 23420
rect 12338 23418 12394 23420
rect 12098 23366 12144 23418
rect 12144 23366 12154 23418
rect 12178 23366 12208 23418
rect 12208 23366 12220 23418
rect 12220 23366 12234 23418
rect 12258 23366 12272 23418
rect 12272 23366 12284 23418
rect 12284 23366 12314 23418
rect 12338 23366 12348 23418
rect 12348 23366 12394 23418
rect 12098 23364 12154 23366
rect 12178 23364 12234 23366
rect 12258 23364 12314 23366
rect 12338 23364 12394 23366
rect 12098 22330 12154 22332
rect 12178 22330 12234 22332
rect 12258 22330 12314 22332
rect 12338 22330 12394 22332
rect 12098 22278 12144 22330
rect 12144 22278 12154 22330
rect 12178 22278 12208 22330
rect 12208 22278 12220 22330
rect 12220 22278 12234 22330
rect 12258 22278 12272 22330
rect 12272 22278 12284 22330
rect 12284 22278 12314 22330
rect 12338 22278 12348 22330
rect 12348 22278 12394 22330
rect 12098 22276 12154 22278
rect 12178 22276 12234 22278
rect 12258 22276 12314 22278
rect 12338 22276 12394 22278
rect 12098 21242 12154 21244
rect 12178 21242 12234 21244
rect 12258 21242 12314 21244
rect 12338 21242 12394 21244
rect 12098 21190 12144 21242
rect 12144 21190 12154 21242
rect 12178 21190 12208 21242
rect 12208 21190 12220 21242
rect 12220 21190 12234 21242
rect 12258 21190 12272 21242
rect 12272 21190 12284 21242
rect 12284 21190 12314 21242
rect 12338 21190 12348 21242
rect 12348 21190 12394 21242
rect 12098 21188 12154 21190
rect 12178 21188 12234 21190
rect 12258 21188 12314 21190
rect 12338 21188 12394 21190
rect 12758 22874 12814 22876
rect 12838 22874 12894 22876
rect 12918 22874 12974 22876
rect 12998 22874 13054 22876
rect 12758 22822 12804 22874
rect 12804 22822 12814 22874
rect 12838 22822 12868 22874
rect 12868 22822 12880 22874
rect 12880 22822 12894 22874
rect 12918 22822 12932 22874
rect 12932 22822 12944 22874
rect 12944 22822 12974 22874
rect 12998 22822 13008 22874
rect 13008 22822 13054 22874
rect 12758 22820 12814 22822
rect 12838 22820 12894 22822
rect 12918 22820 12974 22822
rect 12998 22820 13054 22822
rect 12098 20154 12154 20156
rect 12178 20154 12234 20156
rect 12258 20154 12314 20156
rect 12338 20154 12394 20156
rect 12098 20102 12144 20154
rect 12144 20102 12154 20154
rect 12178 20102 12208 20154
rect 12208 20102 12220 20154
rect 12220 20102 12234 20154
rect 12258 20102 12272 20154
rect 12272 20102 12284 20154
rect 12284 20102 12314 20154
rect 12338 20102 12348 20154
rect 12348 20102 12394 20154
rect 12098 20100 12154 20102
rect 12178 20100 12234 20102
rect 12258 20100 12314 20102
rect 12338 20100 12394 20102
rect 12758 21786 12814 21788
rect 12838 21786 12894 21788
rect 12918 21786 12974 21788
rect 12998 21786 13054 21788
rect 12758 21734 12804 21786
rect 12804 21734 12814 21786
rect 12838 21734 12868 21786
rect 12868 21734 12880 21786
rect 12880 21734 12894 21786
rect 12918 21734 12932 21786
rect 12932 21734 12944 21786
rect 12944 21734 12974 21786
rect 12998 21734 13008 21786
rect 13008 21734 13054 21786
rect 12758 21732 12814 21734
rect 12838 21732 12894 21734
rect 12918 21732 12974 21734
rect 12998 21732 13054 21734
rect 12758 20698 12814 20700
rect 12838 20698 12894 20700
rect 12918 20698 12974 20700
rect 12998 20698 13054 20700
rect 12758 20646 12804 20698
rect 12804 20646 12814 20698
rect 12838 20646 12868 20698
rect 12868 20646 12880 20698
rect 12880 20646 12894 20698
rect 12918 20646 12932 20698
rect 12932 20646 12944 20698
rect 12944 20646 12974 20698
rect 12998 20646 13008 20698
rect 13008 20646 13054 20698
rect 12758 20644 12814 20646
rect 12838 20644 12894 20646
rect 12918 20644 12974 20646
rect 12998 20644 13054 20646
rect 20186 29402 20242 29404
rect 20266 29402 20322 29404
rect 20346 29402 20402 29404
rect 20426 29402 20482 29404
rect 20186 29350 20232 29402
rect 20232 29350 20242 29402
rect 20266 29350 20296 29402
rect 20296 29350 20308 29402
rect 20308 29350 20322 29402
rect 20346 29350 20360 29402
rect 20360 29350 20372 29402
rect 20372 29350 20402 29402
rect 20426 29350 20436 29402
rect 20436 29350 20482 29402
rect 20186 29348 20242 29350
rect 20266 29348 20322 29350
rect 20346 29348 20402 29350
rect 20426 29348 20482 29350
rect 12758 19610 12814 19612
rect 12838 19610 12894 19612
rect 12918 19610 12974 19612
rect 12998 19610 13054 19612
rect 12758 19558 12804 19610
rect 12804 19558 12814 19610
rect 12838 19558 12868 19610
rect 12868 19558 12880 19610
rect 12880 19558 12894 19610
rect 12918 19558 12932 19610
rect 12932 19558 12944 19610
rect 12944 19558 12974 19610
rect 12998 19558 13008 19610
rect 13008 19558 13054 19610
rect 12758 19556 12814 19558
rect 12838 19556 12894 19558
rect 12918 19556 12974 19558
rect 12998 19556 13054 19558
rect 12098 19066 12154 19068
rect 12178 19066 12234 19068
rect 12258 19066 12314 19068
rect 12338 19066 12394 19068
rect 12098 19014 12144 19066
rect 12144 19014 12154 19066
rect 12178 19014 12208 19066
rect 12208 19014 12220 19066
rect 12220 19014 12234 19066
rect 12258 19014 12272 19066
rect 12272 19014 12284 19066
rect 12284 19014 12314 19066
rect 12338 19014 12348 19066
rect 12348 19014 12394 19066
rect 12098 19012 12154 19014
rect 12178 19012 12234 19014
rect 12258 19012 12314 19014
rect 12338 19012 12394 19014
rect 12758 18522 12814 18524
rect 12838 18522 12894 18524
rect 12918 18522 12974 18524
rect 12998 18522 13054 18524
rect 12758 18470 12804 18522
rect 12804 18470 12814 18522
rect 12838 18470 12868 18522
rect 12868 18470 12880 18522
rect 12880 18470 12894 18522
rect 12918 18470 12932 18522
rect 12932 18470 12944 18522
rect 12944 18470 12974 18522
rect 12998 18470 13008 18522
rect 13008 18470 13054 18522
rect 12758 18468 12814 18470
rect 12838 18468 12894 18470
rect 12918 18468 12974 18470
rect 12998 18468 13054 18470
rect 12098 17978 12154 17980
rect 12178 17978 12234 17980
rect 12258 17978 12314 17980
rect 12338 17978 12394 17980
rect 12098 17926 12144 17978
rect 12144 17926 12154 17978
rect 12178 17926 12208 17978
rect 12208 17926 12220 17978
rect 12220 17926 12234 17978
rect 12258 17926 12272 17978
rect 12272 17926 12284 17978
rect 12284 17926 12314 17978
rect 12338 17926 12348 17978
rect 12348 17926 12394 17978
rect 12098 17924 12154 17926
rect 12178 17924 12234 17926
rect 12258 17924 12314 17926
rect 12338 17924 12394 17926
rect 12758 17434 12814 17436
rect 12838 17434 12894 17436
rect 12918 17434 12974 17436
rect 12998 17434 13054 17436
rect 12758 17382 12804 17434
rect 12804 17382 12814 17434
rect 12838 17382 12868 17434
rect 12868 17382 12880 17434
rect 12880 17382 12894 17434
rect 12918 17382 12932 17434
rect 12932 17382 12944 17434
rect 12944 17382 12974 17434
rect 12998 17382 13008 17434
rect 13008 17382 13054 17434
rect 12758 17380 12814 17382
rect 12838 17380 12894 17382
rect 12918 17380 12974 17382
rect 12998 17380 13054 17382
rect 10782 13776 10838 13832
rect 11058 12416 11114 12472
rect 8850 7928 8906 7984
rect 5330 5466 5386 5468
rect 5410 5466 5466 5468
rect 5490 5466 5546 5468
rect 5570 5466 5626 5468
rect 5330 5414 5376 5466
rect 5376 5414 5386 5466
rect 5410 5414 5440 5466
rect 5440 5414 5452 5466
rect 5452 5414 5466 5466
rect 5490 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5546 5466
rect 5570 5414 5580 5466
rect 5580 5414 5626 5466
rect 5330 5412 5386 5414
rect 5410 5412 5466 5414
rect 5490 5412 5546 5414
rect 5570 5412 5626 5414
rect 4670 4922 4726 4924
rect 4750 4922 4806 4924
rect 4830 4922 4886 4924
rect 4910 4922 4966 4924
rect 4670 4870 4716 4922
rect 4716 4870 4726 4922
rect 4750 4870 4780 4922
rect 4780 4870 4792 4922
rect 4792 4870 4806 4922
rect 4830 4870 4844 4922
rect 4844 4870 4856 4922
rect 4856 4870 4886 4922
rect 4910 4870 4920 4922
rect 4920 4870 4966 4922
rect 4670 4868 4726 4870
rect 4750 4868 4806 4870
rect 4830 4868 4886 4870
rect 4910 4868 4966 4870
rect 5330 4378 5386 4380
rect 5410 4378 5466 4380
rect 5490 4378 5546 4380
rect 5570 4378 5626 4380
rect 5330 4326 5376 4378
rect 5376 4326 5386 4378
rect 5410 4326 5440 4378
rect 5440 4326 5452 4378
rect 5452 4326 5466 4378
rect 5490 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5546 4378
rect 5570 4326 5580 4378
rect 5580 4326 5626 4378
rect 5330 4324 5386 4326
rect 5410 4324 5466 4326
rect 5490 4324 5546 4326
rect 5570 4324 5626 4326
rect 4670 3834 4726 3836
rect 4750 3834 4806 3836
rect 4830 3834 4886 3836
rect 4910 3834 4966 3836
rect 4670 3782 4716 3834
rect 4716 3782 4726 3834
rect 4750 3782 4780 3834
rect 4780 3782 4792 3834
rect 4792 3782 4806 3834
rect 4830 3782 4844 3834
rect 4844 3782 4856 3834
rect 4856 3782 4886 3834
rect 4910 3782 4920 3834
rect 4920 3782 4966 3834
rect 4670 3780 4726 3782
rect 4750 3780 4806 3782
rect 4830 3780 4886 3782
rect 4910 3780 4966 3782
rect 5330 3290 5386 3292
rect 5410 3290 5466 3292
rect 5490 3290 5546 3292
rect 5570 3290 5626 3292
rect 5330 3238 5376 3290
rect 5376 3238 5386 3290
rect 5410 3238 5440 3290
rect 5440 3238 5452 3290
rect 5452 3238 5466 3290
rect 5490 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5546 3290
rect 5570 3238 5580 3290
rect 5580 3238 5626 3290
rect 5330 3236 5386 3238
rect 5410 3236 5466 3238
rect 5490 3236 5546 3238
rect 5570 3236 5626 3238
rect 4670 2746 4726 2748
rect 4750 2746 4806 2748
rect 4830 2746 4886 2748
rect 4910 2746 4966 2748
rect 4670 2694 4716 2746
rect 4716 2694 4726 2746
rect 4750 2694 4780 2746
rect 4780 2694 4792 2746
rect 4792 2694 4806 2746
rect 4830 2694 4844 2746
rect 4844 2694 4856 2746
rect 4856 2694 4886 2746
rect 4910 2694 4920 2746
rect 4920 2694 4966 2746
rect 4670 2692 4726 2694
rect 4750 2692 4806 2694
rect 4830 2692 4886 2694
rect 4910 2692 4966 2694
rect 5330 2202 5386 2204
rect 5410 2202 5466 2204
rect 5490 2202 5546 2204
rect 5570 2202 5626 2204
rect 5330 2150 5376 2202
rect 5376 2150 5386 2202
rect 5410 2150 5440 2202
rect 5440 2150 5452 2202
rect 5452 2150 5466 2202
rect 5490 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5546 2202
rect 5570 2150 5580 2202
rect 5580 2150 5626 2202
rect 5330 2148 5386 2150
rect 5410 2148 5466 2150
rect 5490 2148 5546 2150
rect 5570 2148 5626 2150
rect 12098 16890 12154 16892
rect 12178 16890 12234 16892
rect 12258 16890 12314 16892
rect 12338 16890 12394 16892
rect 12098 16838 12144 16890
rect 12144 16838 12154 16890
rect 12178 16838 12208 16890
rect 12208 16838 12220 16890
rect 12220 16838 12234 16890
rect 12258 16838 12272 16890
rect 12272 16838 12284 16890
rect 12284 16838 12314 16890
rect 12338 16838 12348 16890
rect 12348 16838 12394 16890
rect 12098 16836 12154 16838
rect 12178 16836 12234 16838
rect 12258 16836 12314 16838
rect 12338 16836 12394 16838
rect 12758 16346 12814 16348
rect 12838 16346 12894 16348
rect 12918 16346 12974 16348
rect 12998 16346 13054 16348
rect 12758 16294 12804 16346
rect 12804 16294 12814 16346
rect 12838 16294 12868 16346
rect 12868 16294 12880 16346
rect 12880 16294 12894 16346
rect 12918 16294 12932 16346
rect 12932 16294 12944 16346
rect 12944 16294 12974 16346
rect 12998 16294 13008 16346
rect 13008 16294 13054 16346
rect 12758 16292 12814 16294
rect 12838 16292 12894 16294
rect 12918 16292 12974 16294
rect 12998 16292 13054 16294
rect 12098 15802 12154 15804
rect 12178 15802 12234 15804
rect 12258 15802 12314 15804
rect 12338 15802 12394 15804
rect 12098 15750 12144 15802
rect 12144 15750 12154 15802
rect 12178 15750 12208 15802
rect 12208 15750 12220 15802
rect 12220 15750 12234 15802
rect 12258 15750 12272 15802
rect 12272 15750 12284 15802
rect 12284 15750 12314 15802
rect 12338 15750 12348 15802
rect 12348 15750 12394 15802
rect 12098 15748 12154 15750
rect 12178 15748 12234 15750
rect 12258 15748 12314 15750
rect 12338 15748 12394 15750
rect 12530 15408 12586 15464
rect 12098 14714 12154 14716
rect 12178 14714 12234 14716
rect 12258 14714 12314 14716
rect 12338 14714 12394 14716
rect 12098 14662 12144 14714
rect 12144 14662 12154 14714
rect 12178 14662 12208 14714
rect 12208 14662 12220 14714
rect 12220 14662 12234 14714
rect 12258 14662 12272 14714
rect 12272 14662 12284 14714
rect 12284 14662 12314 14714
rect 12338 14662 12348 14714
rect 12348 14662 12394 14714
rect 12098 14660 12154 14662
rect 12178 14660 12234 14662
rect 12258 14660 12314 14662
rect 12338 14660 12394 14662
rect 11610 12416 11666 12472
rect 9586 7928 9642 7984
rect 12098 13626 12154 13628
rect 12178 13626 12234 13628
rect 12258 13626 12314 13628
rect 12338 13626 12394 13628
rect 12098 13574 12144 13626
rect 12144 13574 12154 13626
rect 12178 13574 12208 13626
rect 12208 13574 12220 13626
rect 12220 13574 12234 13626
rect 12258 13574 12272 13626
rect 12272 13574 12284 13626
rect 12284 13574 12314 13626
rect 12338 13574 12348 13626
rect 12348 13574 12394 13626
rect 12098 13572 12154 13574
rect 12178 13572 12234 13574
rect 12258 13572 12314 13574
rect 12338 13572 12394 13574
rect 12098 12538 12154 12540
rect 12178 12538 12234 12540
rect 12258 12538 12314 12540
rect 12338 12538 12394 12540
rect 12098 12486 12144 12538
rect 12144 12486 12154 12538
rect 12178 12486 12208 12538
rect 12208 12486 12220 12538
rect 12220 12486 12234 12538
rect 12258 12486 12272 12538
rect 12272 12486 12284 12538
rect 12284 12486 12314 12538
rect 12338 12486 12348 12538
rect 12348 12486 12394 12538
rect 12098 12484 12154 12486
rect 12178 12484 12234 12486
rect 12258 12484 12314 12486
rect 12338 12484 12394 12486
rect 12098 11450 12154 11452
rect 12178 11450 12234 11452
rect 12258 11450 12314 11452
rect 12338 11450 12394 11452
rect 12098 11398 12144 11450
rect 12144 11398 12154 11450
rect 12178 11398 12208 11450
rect 12208 11398 12220 11450
rect 12220 11398 12234 11450
rect 12258 11398 12272 11450
rect 12272 11398 12284 11450
rect 12284 11398 12314 11450
rect 12338 11398 12348 11450
rect 12348 11398 12394 11450
rect 12098 11396 12154 11398
rect 12178 11396 12234 11398
rect 12258 11396 12314 11398
rect 12338 11396 12394 11398
rect 12098 10362 12154 10364
rect 12178 10362 12234 10364
rect 12258 10362 12314 10364
rect 12338 10362 12394 10364
rect 12098 10310 12144 10362
rect 12144 10310 12154 10362
rect 12178 10310 12208 10362
rect 12208 10310 12220 10362
rect 12220 10310 12234 10362
rect 12258 10310 12272 10362
rect 12272 10310 12284 10362
rect 12284 10310 12314 10362
rect 12338 10310 12348 10362
rect 12348 10310 12394 10362
rect 12098 10308 12154 10310
rect 12178 10308 12234 10310
rect 12258 10308 12314 10310
rect 12338 10308 12394 10310
rect 12758 15258 12814 15260
rect 12838 15258 12894 15260
rect 12918 15258 12974 15260
rect 12998 15258 13054 15260
rect 12758 15206 12804 15258
rect 12804 15206 12814 15258
rect 12838 15206 12868 15258
rect 12868 15206 12880 15258
rect 12880 15206 12894 15258
rect 12918 15206 12932 15258
rect 12932 15206 12944 15258
rect 12944 15206 12974 15258
rect 12998 15206 13008 15258
rect 13008 15206 13054 15258
rect 12758 15204 12814 15206
rect 12838 15204 12894 15206
rect 12918 15204 12974 15206
rect 12998 15204 13054 15206
rect 12758 14170 12814 14172
rect 12838 14170 12894 14172
rect 12918 14170 12974 14172
rect 12998 14170 13054 14172
rect 12758 14118 12804 14170
rect 12804 14118 12814 14170
rect 12838 14118 12868 14170
rect 12868 14118 12880 14170
rect 12880 14118 12894 14170
rect 12918 14118 12932 14170
rect 12932 14118 12944 14170
rect 12944 14118 12974 14170
rect 12998 14118 13008 14170
rect 13008 14118 13054 14170
rect 12758 14116 12814 14118
rect 12838 14116 12894 14118
rect 12918 14116 12974 14118
rect 12998 14116 13054 14118
rect 14554 21256 14610 21312
rect 13726 15444 13728 15464
rect 13728 15444 13780 15464
rect 13780 15444 13782 15464
rect 13726 15408 13782 15444
rect 12758 13082 12814 13084
rect 12838 13082 12894 13084
rect 12918 13082 12974 13084
rect 12998 13082 13054 13084
rect 12758 13030 12804 13082
rect 12804 13030 12814 13082
rect 12838 13030 12868 13082
rect 12868 13030 12880 13082
rect 12880 13030 12894 13082
rect 12918 13030 12932 13082
rect 12932 13030 12944 13082
rect 12944 13030 12974 13082
rect 12998 13030 13008 13082
rect 13008 13030 13054 13082
rect 12758 13028 12814 13030
rect 12838 13028 12894 13030
rect 12918 13028 12974 13030
rect 12998 13028 13054 13030
rect 12758 11994 12814 11996
rect 12838 11994 12894 11996
rect 12918 11994 12974 11996
rect 12998 11994 13054 11996
rect 12758 11942 12804 11994
rect 12804 11942 12814 11994
rect 12838 11942 12868 11994
rect 12868 11942 12880 11994
rect 12880 11942 12894 11994
rect 12918 11942 12932 11994
rect 12932 11942 12944 11994
rect 12944 11942 12974 11994
rect 12998 11942 13008 11994
rect 13008 11942 13054 11994
rect 12758 11940 12814 11942
rect 12838 11940 12894 11942
rect 12918 11940 12974 11942
rect 12998 11940 13054 11942
rect 12758 10906 12814 10908
rect 12838 10906 12894 10908
rect 12918 10906 12974 10908
rect 12998 10906 13054 10908
rect 12758 10854 12804 10906
rect 12804 10854 12814 10906
rect 12838 10854 12868 10906
rect 12868 10854 12880 10906
rect 12880 10854 12894 10906
rect 12918 10854 12932 10906
rect 12932 10854 12944 10906
rect 12944 10854 12974 10906
rect 12998 10854 13008 10906
rect 13008 10854 13054 10906
rect 12758 10852 12814 10854
rect 12838 10852 12894 10854
rect 12918 10852 12974 10854
rect 12998 10852 13054 10854
rect 12098 9274 12154 9276
rect 12178 9274 12234 9276
rect 12258 9274 12314 9276
rect 12338 9274 12394 9276
rect 12098 9222 12144 9274
rect 12144 9222 12154 9274
rect 12178 9222 12208 9274
rect 12208 9222 12220 9274
rect 12220 9222 12234 9274
rect 12258 9222 12272 9274
rect 12272 9222 12284 9274
rect 12284 9222 12314 9274
rect 12338 9222 12348 9274
rect 12348 9222 12394 9274
rect 12098 9220 12154 9222
rect 12178 9220 12234 9222
rect 12258 9220 12314 9222
rect 12338 9220 12394 9222
rect 12758 9818 12814 9820
rect 12838 9818 12894 9820
rect 12918 9818 12974 9820
rect 12998 9818 13054 9820
rect 12758 9766 12804 9818
rect 12804 9766 12814 9818
rect 12838 9766 12868 9818
rect 12868 9766 12880 9818
rect 12880 9766 12894 9818
rect 12918 9766 12932 9818
rect 12932 9766 12944 9818
rect 12944 9766 12974 9818
rect 12998 9766 13008 9818
rect 13008 9766 13054 9818
rect 12758 9764 12814 9766
rect 12838 9764 12894 9766
rect 12918 9764 12974 9766
rect 12998 9764 13054 9766
rect 19526 28858 19582 28860
rect 19606 28858 19662 28860
rect 19686 28858 19742 28860
rect 19766 28858 19822 28860
rect 19526 28806 19572 28858
rect 19572 28806 19582 28858
rect 19606 28806 19636 28858
rect 19636 28806 19648 28858
rect 19648 28806 19662 28858
rect 19686 28806 19700 28858
rect 19700 28806 19712 28858
rect 19712 28806 19742 28858
rect 19766 28806 19776 28858
rect 19776 28806 19822 28858
rect 19526 28804 19582 28806
rect 19606 28804 19662 28806
rect 19686 28804 19742 28806
rect 19766 28804 19822 28806
rect 20186 28314 20242 28316
rect 20266 28314 20322 28316
rect 20346 28314 20402 28316
rect 20426 28314 20482 28316
rect 20186 28262 20232 28314
rect 20232 28262 20242 28314
rect 20266 28262 20296 28314
rect 20296 28262 20308 28314
rect 20308 28262 20322 28314
rect 20346 28262 20360 28314
rect 20360 28262 20372 28314
rect 20372 28262 20402 28314
rect 20426 28262 20436 28314
rect 20436 28262 20482 28314
rect 20186 28260 20242 28262
rect 20266 28260 20322 28262
rect 20346 28260 20402 28262
rect 20426 28260 20482 28262
rect 19526 27770 19582 27772
rect 19606 27770 19662 27772
rect 19686 27770 19742 27772
rect 19766 27770 19822 27772
rect 19526 27718 19572 27770
rect 19572 27718 19582 27770
rect 19606 27718 19636 27770
rect 19636 27718 19648 27770
rect 19648 27718 19662 27770
rect 19686 27718 19700 27770
rect 19700 27718 19712 27770
rect 19712 27718 19742 27770
rect 19766 27718 19776 27770
rect 19776 27718 19822 27770
rect 19526 27716 19582 27718
rect 19606 27716 19662 27718
rect 19686 27716 19742 27718
rect 19766 27716 19822 27718
rect 27614 29402 27670 29404
rect 27694 29402 27750 29404
rect 27774 29402 27830 29404
rect 27854 29402 27910 29404
rect 27614 29350 27660 29402
rect 27660 29350 27670 29402
rect 27694 29350 27724 29402
rect 27724 29350 27736 29402
rect 27736 29350 27750 29402
rect 27774 29350 27788 29402
rect 27788 29350 27800 29402
rect 27800 29350 27830 29402
rect 27854 29350 27864 29402
rect 27864 29350 27910 29402
rect 27614 29348 27670 29350
rect 27694 29348 27750 29350
rect 27774 29348 27830 29350
rect 27854 29348 27910 29350
rect 26954 28858 27010 28860
rect 27034 28858 27090 28860
rect 27114 28858 27170 28860
rect 27194 28858 27250 28860
rect 26954 28806 27000 28858
rect 27000 28806 27010 28858
rect 27034 28806 27064 28858
rect 27064 28806 27076 28858
rect 27076 28806 27090 28858
rect 27114 28806 27128 28858
rect 27128 28806 27140 28858
rect 27140 28806 27170 28858
rect 27194 28806 27204 28858
rect 27204 28806 27250 28858
rect 26954 28804 27010 28806
rect 27034 28804 27090 28806
rect 27114 28804 27170 28806
rect 27194 28804 27250 28806
rect 27614 28314 27670 28316
rect 27694 28314 27750 28316
rect 27774 28314 27830 28316
rect 27854 28314 27910 28316
rect 27614 28262 27660 28314
rect 27660 28262 27670 28314
rect 27694 28262 27724 28314
rect 27724 28262 27736 28314
rect 27736 28262 27750 28314
rect 27774 28262 27788 28314
rect 27788 28262 27800 28314
rect 27800 28262 27830 28314
rect 27854 28262 27864 28314
rect 27864 28262 27910 28314
rect 27614 28260 27670 28262
rect 27694 28260 27750 28262
rect 27774 28260 27830 28262
rect 27854 28260 27910 28262
rect 26954 27770 27010 27772
rect 27034 27770 27090 27772
rect 27114 27770 27170 27772
rect 27194 27770 27250 27772
rect 26954 27718 27000 27770
rect 27000 27718 27010 27770
rect 27034 27718 27064 27770
rect 27064 27718 27076 27770
rect 27076 27718 27090 27770
rect 27114 27718 27128 27770
rect 27128 27718 27140 27770
rect 27140 27718 27170 27770
rect 27194 27718 27204 27770
rect 27204 27718 27250 27770
rect 26954 27716 27010 27718
rect 27034 27716 27090 27718
rect 27114 27716 27170 27718
rect 27194 27716 27250 27718
rect 20186 27226 20242 27228
rect 20266 27226 20322 27228
rect 20346 27226 20402 27228
rect 20426 27226 20482 27228
rect 20186 27174 20232 27226
rect 20232 27174 20242 27226
rect 20266 27174 20296 27226
rect 20296 27174 20308 27226
rect 20308 27174 20322 27226
rect 20346 27174 20360 27226
rect 20360 27174 20372 27226
rect 20372 27174 20402 27226
rect 20426 27174 20436 27226
rect 20436 27174 20482 27226
rect 20186 27172 20242 27174
rect 20266 27172 20322 27174
rect 20346 27172 20402 27174
rect 20426 27172 20482 27174
rect 19526 26682 19582 26684
rect 19606 26682 19662 26684
rect 19686 26682 19742 26684
rect 19766 26682 19822 26684
rect 19526 26630 19572 26682
rect 19572 26630 19582 26682
rect 19606 26630 19636 26682
rect 19636 26630 19648 26682
rect 19648 26630 19662 26682
rect 19686 26630 19700 26682
rect 19700 26630 19712 26682
rect 19712 26630 19742 26682
rect 19766 26630 19776 26682
rect 19776 26630 19822 26682
rect 19526 26628 19582 26630
rect 19606 26628 19662 26630
rect 19686 26628 19742 26630
rect 19766 26628 19822 26630
rect 20186 26138 20242 26140
rect 20266 26138 20322 26140
rect 20346 26138 20402 26140
rect 20426 26138 20482 26140
rect 20186 26086 20232 26138
rect 20232 26086 20242 26138
rect 20266 26086 20296 26138
rect 20296 26086 20308 26138
rect 20308 26086 20322 26138
rect 20346 26086 20360 26138
rect 20360 26086 20372 26138
rect 20372 26086 20402 26138
rect 20426 26086 20436 26138
rect 20436 26086 20482 26138
rect 20186 26084 20242 26086
rect 20266 26084 20322 26086
rect 20346 26084 20402 26086
rect 20426 26084 20482 26086
rect 19526 25594 19582 25596
rect 19606 25594 19662 25596
rect 19686 25594 19742 25596
rect 19766 25594 19822 25596
rect 19526 25542 19572 25594
rect 19572 25542 19582 25594
rect 19606 25542 19636 25594
rect 19636 25542 19648 25594
rect 19648 25542 19662 25594
rect 19686 25542 19700 25594
rect 19700 25542 19712 25594
rect 19712 25542 19742 25594
rect 19766 25542 19776 25594
rect 19776 25542 19822 25594
rect 19526 25540 19582 25542
rect 19606 25540 19662 25542
rect 19686 25540 19742 25542
rect 19766 25540 19822 25542
rect 20186 25050 20242 25052
rect 20266 25050 20322 25052
rect 20346 25050 20402 25052
rect 20426 25050 20482 25052
rect 20186 24998 20232 25050
rect 20232 24998 20242 25050
rect 20266 24998 20296 25050
rect 20296 24998 20308 25050
rect 20308 24998 20322 25050
rect 20346 24998 20360 25050
rect 20360 24998 20372 25050
rect 20372 24998 20402 25050
rect 20426 24998 20436 25050
rect 20436 24998 20482 25050
rect 20186 24996 20242 24998
rect 20266 24996 20322 24998
rect 20346 24996 20402 24998
rect 20426 24996 20482 24998
rect 19526 24506 19582 24508
rect 19606 24506 19662 24508
rect 19686 24506 19742 24508
rect 19766 24506 19822 24508
rect 19526 24454 19572 24506
rect 19572 24454 19582 24506
rect 19606 24454 19636 24506
rect 19636 24454 19648 24506
rect 19648 24454 19662 24506
rect 19686 24454 19700 24506
rect 19700 24454 19712 24506
rect 19712 24454 19742 24506
rect 19766 24454 19776 24506
rect 19776 24454 19822 24506
rect 19526 24452 19582 24454
rect 19606 24452 19662 24454
rect 19686 24452 19742 24454
rect 19766 24452 19822 24454
rect 20186 23962 20242 23964
rect 20266 23962 20322 23964
rect 20346 23962 20402 23964
rect 20426 23962 20482 23964
rect 20186 23910 20232 23962
rect 20232 23910 20242 23962
rect 20266 23910 20296 23962
rect 20296 23910 20308 23962
rect 20308 23910 20322 23962
rect 20346 23910 20360 23962
rect 20360 23910 20372 23962
rect 20372 23910 20402 23962
rect 20426 23910 20436 23962
rect 20436 23910 20482 23962
rect 20186 23908 20242 23910
rect 20266 23908 20322 23910
rect 20346 23908 20402 23910
rect 20426 23908 20482 23910
rect 19526 23418 19582 23420
rect 19606 23418 19662 23420
rect 19686 23418 19742 23420
rect 19766 23418 19822 23420
rect 19526 23366 19572 23418
rect 19572 23366 19582 23418
rect 19606 23366 19636 23418
rect 19636 23366 19648 23418
rect 19648 23366 19662 23418
rect 19686 23366 19700 23418
rect 19700 23366 19712 23418
rect 19712 23366 19742 23418
rect 19766 23366 19776 23418
rect 19776 23366 19822 23418
rect 19526 23364 19582 23366
rect 19606 23364 19662 23366
rect 19686 23364 19742 23366
rect 19766 23364 19822 23366
rect 12098 8186 12154 8188
rect 12178 8186 12234 8188
rect 12258 8186 12314 8188
rect 12338 8186 12394 8188
rect 12098 8134 12144 8186
rect 12144 8134 12154 8186
rect 12178 8134 12208 8186
rect 12208 8134 12220 8186
rect 12220 8134 12234 8186
rect 12258 8134 12272 8186
rect 12272 8134 12284 8186
rect 12284 8134 12314 8186
rect 12338 8134 12348 8186
rect 12348 8134 12394 8186
rect 12098 8132 12154 8134
rect 12178 8132 12234 8134
rect 12258 8132 12314 8134
rect 12338 8132 12394 8134
rect 12758 8730 12814 8732
rect 12838 8730 12894 8732
rect 12918 8730 12974 8732
rect 12998 8730 13054 8732
rect 12758 8678 12804 8730
rect 12804 8678 12814 8730
rect 12838 8678 12868 8730
rect 12868 8678 12880 8730
rect 12880 8678 12894 8730
rect 12918 8678 12932 8730
rect 12932 8678 12944 8730
rect 12944 8678 12974 8730
rect 12998 8678 13008 8730
rect 13008 8678 13054 8730
rect 12758 8676 12814 8678
rect 12838 8676 12894 8678
rect 12918 8676 12974 8678
rect 12998 8676 13054 8678
rect 15934 15408 15990 15464
rect 18326 21256 18382 21312
rect 19526 22330 19582 22332
rect 19606 22330 19662 22332
rect 19686 22330 19742 22332
rect 19766 22330 19822 22332
rect 19526 22278 19572 22330
rect 19572 22278 19582 22330
rect 19606 22278 19636 22330
rect 19636 22278 19648 22330
rect 19648 22278 19662 22330
rect 19686 22278 19700 22330
rect 19700 22278 19712 22330
rect 19712 22278 19742 22330
rect 19766 22278 19776 22330
rect 19776 22278 19822 22330
rect 19526 22276 19582 22278
rect 19606 22276 19662 22278
rect 19686 22276 19742 22278
rect 19766 22276 19822 22278
rect 20186 22874 20242 22876
rect 20266 22874 20322 22876
rect 20346 22874 20402 22876
rect 20426 22874 20482 22876
rect 20186 22822 20232 22874
rect 20232 22822 20242 22874
rect 20266 22822 20296 22874
rect 20296 22822 20308 22874
rect 20308 22822 20322 22874
rect 20346 22822 20360 22874
rect 20360 22822 20372 22874
rect 20372 22822 20402 22874
rect 20426 22822 20436 22874
rect 20436 22822 20482 22874
rect 20186 22820 20242 22822
rect 20266 22820 20322 22822
rect 20346 22820 20402 22822
rect 20426 22820 20482 22822
rect 20186 21786 20242 21788
rect 20266 21786 20322 21788
rect 20346 21786 20402 21788
rect 20426 21786 20482 21788
rect 20186 21734 20232 21786
rect 20232 21734 20242 21786
rect 20266 21734 20296 21786
rect 20296 21734 20308 21786
rect 20308 21734 20322 21786
rect 20346 21734 20360 21786
rect 20360 21734 20372 21786
rect 20372 21734 20402 21786
rect 20426 21734 20436 21786
rect 20436 21734 20482 21786
rect 20186 21732 20242 21734
rect 20266 21732 20322 21734
rect 20346 21732 20402 21734
rect 20426 21732 20482 21734
rect 19526 21242 19582 21244
rect 19606 21242 19662 21244
rect 19686 21242 19742 21244
rect 19766 21242 19822 21244
rect 19526 21190 19572 21242
rect 19572 21190 19582 21242
rect 19606 21190 19636 21242
rect 19636 21190 19648 21242
rect 19648 21190 19662 21242
rect 19686 21190 19700 21242
rect 19700 21190 19712 21242
rect 19712 21190 19742 21242
rect 19766 21190 19776 21242
rect 19776 21190 19822 21242
rect 19526 21188 19582 21190
rect 19606 21188 19662 21190
rect 19686 21188 19742 21190
rect 19766 21188 19822 21190
rect 27614 27226 27670 27228
rect 27694 27226 27750 27228
rect 27774 27226 27830 27228
rect 27854 27226 27910 27228
rect 27614 27174 27660 27226
rect 27660 27174 27670 27226
rect 27694 27174 27724 27226
rect 27724 27174 27736 27226
rect 27736 27174 27750 27226
rect 27774 27174 27788 27226
rect 27788 27174 27800 27226
rect 27800 27174 27830 27226
rect 27854 27174 27864 27226
rect 27864 27174 27910 27226
rect 27614 27172 27670 27174
rect 27694 27172 27750 27174
rect 27774 27172 27830 27174
rect 27854 27172 27910 27174
rect 26954 26682 27010 26684
rect 27034 26682 27090 26684
rect 27114 26682 27170 26684
rect 27194 26682 27250 26684
rect 26954 26630 27000 26682
rect 27000 26630 27010 26682
rect 27034 26630 27064 26682
rect 27064 26630 27076 26682
rect 27076 26630 27090 26682
rect 27114 26630 27128 26682
rect 27128 26630 27140 26682
rect 27140 26630 27170 26682
rect 27194 26630 27204 26682
rect 27204 26630 27250 26682
rect 26954 26628 27010 26630
rect 27034 26628 27090 26630
rect 27114 26628 27170 26630
rect 27194 26628 27250 26630
rect 27614 26138 27670 26140
rect 27694 26138 27750 26140
rect 27774 26138 27830 26140
rect 27854 26138 27910 26140
rect 27614 26086 27660 26138
rect 27660 26086 27670 26138
rect 27694 26086 27724 26138
rect 27724 26086 27736 26138
rect 27736 26086 27750 26138
rect 27774 26086 27788 26138
rect 27788 26086 27800 26138
rect 27800 26086 27830 26138
rect 27854 26086 27864 26138
rect 27864 26086 27910 26138
rect 27614 26084 27670 26086
rect 27694 26084 27750 26086
rect 27774 26084 27830 26086
rect 27854 26084 27910 26086
rect 26954 25594 27010 25596
rect 27034 25594 27090 25596
rect 27114 25594 27170 25596
rect 27194 25594 27250 25596
rect 26954 25542 27000 25594
rect 27000 25542 27010 25594
rect 27034 25542 27064 25594
rect 27064 25542 27076 25594
rect 27076 25542 27090 25594
rect 27114 25542 27128 25594
rect 27128 25542 27140 25594
rect 27140 25542 27170 25594
rect 27194 25542 27204 25594
rect 27204 25542 27250 25594
rect 26954 25540 27010 25542
rect 27034 25540 27090 25542
rect 27114 25540 27170 25542
rect 27194 25540 27250 25542
rect 27614 25050 27670 25052
rect 27694 25050 27750 25052
rect 27774 25050 27830 25052
rect 27854 25050 27910 25052
rect 27614 24998 27660 25050
rect 27660 24998 27670 25050
rect 27694 24998 27724 25050
rect 27724 24998 27736 25050
rect 27736 24998 27750 25050
rect 27774 24998 27788 25050
rect 27788 24998 27800 25050
rect 27800 24998 27830 25050
rect 27854 24998 27864 25050
rect 27864 24998 27910 25050
rect 27614 24996 27670 24998
rect 27694 24996 27750 24998
rect 27774 24996 27830 24998
rect 27854 24996 27910 24998
rect 26954 24506 27010 24508
rect 27034 24506 27090 24508
rect 27114 24506 27170 24508
rect 27194 24506 27250 24508
rect 26954 24454 27000 24506
rect 27000 24454 27010 24506
rect 27034 24454 27064 24506
rect 27064 24454 27076 24506
rect 27076 24454 27090 24506
rect 27114 24454 27128 24506
rect 27128 24454 27140 24506
rect 27140 24454 27170 24506
rect 27194 24454 27204 24506
rect 27204 24454 27250 24506
rect 26954 24452 27010 24454
rect 27034 24452 27090 24454
rect 27114 24452 27170 24454
rect 27194 24452 27250 24454
rect 27614 23962 27670 23964
rect 27694 23962 27750 23964
rect 27774 23962 27830 23964
rect 27854 23962 27910 23964
rect 27614 23910 27660 23962
rect 27660 23910 27670 23962
rect 27694 23910 27724 23962
rect 27724 23910 27736 23962
rect 27736 23910 27750 23962
rect 27774 23910 27788 23962
rect 27788 23910 27800 23962
rect 27800 23910 27830 23962
rect 27854 23910 27864 23962
rect 27864 23910 27910 23962
rect 27614 23908 27670 23910
rect 27694 23908 27750 23910
rect 27774 23908 27830 23910
rect 27854 23908 27910 23910
rect 21822 21956 21878 21992
rect 21822 21936 21824 21956
rect 21824 21936 21876 21956
rect 21876 21936 21878 21956
rect 19526 20154 19582 20156
rect 19606 20154 19662 20156
rect 19686 20154 19742 20156
rect 19766 20154 19822 20156
rect 19526 20102 19572 20154
rect 19572 20102 19582 20154
rect 19606 20102 19636 20154
rect 19636 20102 19648 20154
rect 19648 20102 19662 20154
rect 19686 20102 19700 20154
rect 19700 20102 19712 20154
rect 19712 20102 19742 20154
rect 19766 20102 19776 20154
rect 19776 20102 19822 20154
rect 19526 20100 19582 20102
rect 19606 20100 19662 20102
rect 19686 20100 19742 20102
rect 19766 20100 19822 20102
rect 12758 7642 12814 7644
rect 12838 7642 12894 7644
rect 12918 7642 12974 7644
rect 12998 7642 13054 7644
rect 12758 7590 12804 7642
rect 12804 7590 12814 7642
rect 12838 7590 12868 7642
rect 12868 7590 12880 7642
rect 12880 7590 12894 7642
rect 12918 7590 12932 7642
rect 12932 7590 12944 7642
rect 12944 7590 12974 7642
rect 12998 7590 13008 7642
rect 13008 7590 13054 7642
rect 12758 7588 12814 7590
rect 12838 7588 12894 7590
rect 12918 7588 12974 7590
rect 12998 7588 13054 7590
rect 12098 7098 12154 7100
rect 12178 7098 12234 7100
rect 12258 7098 12314 7100
rect 12338 7098 12394 7100
rect 12098 7046 12144 7098
rect 12144 7046 12154 7098
rect 12178 7046 12208 7098
rect 12208 7046 12220 7098
rect 12220 7046 12234 7098
rect 12258 7046 12272 7098
rect 12272 7046 12284 7098
rect 12284 7046 12314 7098
rect 12338 7046 12348 7098
rect 12348 7046 12394 7098
rect 12098 7044 12154 7046
rect 12178 7044 12234 7046
rect 12258 7044 12314 7046
rect 12338 7044 12394 7046
rect 12758 6554 12814 6556
rect 12838 6554 12894 6556
rect 12918 6554 12974 6556
rect 12998 6554 13054 6556
rect 12758 6502 12804 6554
rect 12804 6502 12814 6554
rect 12838 6502 12868 6554
rect 12868 6502 12880 6554
rect 12880 6502 12894 6554
rect 12918 6502 12932 6554
rect 12932 6502 12944 6554
rect 12944 6502 12974 6554
rect 12998 6502 13008 6554
rect 13008 6502 13054 6554
rect 12758 6500 12814 6502
rect 12838 6500 12894 6502
rect 12918 6500 12974 6502
rect 12998 6500 13054 6502
rect 12098 6010 12154 6012
rect 12178 6010 12234 6012
rect 12258 6010 12314 6012
rect 12338 6010 12394 6012
rect 12098 5958 12144 6010
rect 12144 5958 12154 6010
rect 12178 5958 12208 6010
rect 12208 5958 12220 6010
rect 12220 5958 12234 6010
rect 12258 5958 12272 6010
rect 12272 5958 12284 6010
rect 12284 5958 12314 6010
rect 12338 5958 12348 6010
rect 12348 5958 12394 6010
rect 12098 5956 12154 5958
rect 12178 5956 12234 5958
rect 12258 5956 12314 5958
rect 12338 5956 12394 5958
rect 12758 5466 12814 5468
rect 12838 5466 12894 5468
rect 12918 5466 12974 5468
rect 12998 5466 13054 5468
rect 12758 5414 12804 5466
rect 12804 5414 12814 5466
rect 12838 5414 12868 5466
rect 12868 5414 12880 5466
rect 12880 5414 12894 5466
rect 12918 5414 12932 5466
rect 12932 5414 12944 5466
rect 12944 5414 12974 5466
rect 12998 5414 13008 5466
rect 13008 5414 13054 5466
rect 12758 5412 12814 5414
rect 12838 5412 12894 5414
rect 12918 5412 12974 5414
rect 12998 5412 13054 5414
rect 12098 4922 12154 4924
rect 12178 4922 12234 4924
rect 12258 4922 12314 4924
rect 12338 4922 12394 4924
rect 12098 4870 12144 4922
rect 12144 4870 12154 4922
rect 12178 4870 12208 4922
rect 12208 4870 12220 4922
rect 12220 4870 12234 4922
rect 12258 4870 12272 4922
rect 12272 4870 12284 4922
rect 12284 4870 12314 4922
rect 12338 4870 12348 4922
rect 12348 4870 12394 4922
rect 12098 4868 12154 4870
rect 12178 4868 12234 4870
rect 12258 4868 12314 4870
rect 12338 4868 12394 4870
rect 12758 4378 12814 4380
rect 12838 4378 12894 4380
rect 12918 4378 12974 4380
rect 12998 4378 13054 4380
rect 12758 4326 12804 4378
rect 12804 4326 12814 4378
rect 12838 4326 12868 4378
rect 12868 4326 12880 4378
rect 12880 4326 12894 4378
rect 12918 4326 12932 4378
rect 12932 4326 12944 4378
rect 12944 4326 12974 4378
rect 12998 4326 13008 4378
rect 13008 4326 13054 4378
rect 12758 4324 12814 4326
rect 12838 4324 12894 4326
rect 12918 4324 12974 4326
rect 12998 4324 13054 4326
rect 12098 3834 12154 3836
rect 12178 3834 12234 3836
rect 12258 3834 12314 3836
rect 12338 3834 12394 3836
rect 12098 3782 12144 3834
rect 12144 3782 12154 3834
rect 12178 3782 12208 3834
rect 12208 3782 12220 3834
rect 12220 3782 12234 3834
rect 12258 3782 12272 3834
rect 12272 3782 12284 3834
rect 12284 3782 12314 3834
rect 12338 3782 12348 3834
rect 12348 3782 12394 3834
rect 12098 3780 12154 3782
rect 12178 3780 12234 3782
rect 12258 3780 12314 3782
rect 12338 3780 12394 3782
rect 12758 3290 12814 3292
rect 12838 3290 12894 3292
rect 12918 3290 12974 3292
rect 12998 3290 13054 3292
rect 12758 3238 12804 3290
rect 12804 3238 12814 3290
rect 12838 3238 12868 3290
rect 12868 3238 12880 3290
rect 12880 3238 12894 3290
rect 12918 3238 12932 3290
rect 12932 3238 12944 3290
rect 12944 3238 12974 3290
rect 12998 3238 13008 3290
rect 13008 3238 13054 3290
rect 12758 3236 12814 3238
rect 12838 3236 12894 3238
rect 12918 3236 12974 3238
rect 12998 3236 13054 3238
rect 12098 2746 12154 2748
rect 12178 2746 12234 2748
rect 12258 2746 12314 2748
rect 12338 2746 12394 2748
rect 12098 2694 12144 2746
rect 12144 2694 12154 2746
rect 12178 2694 12208 2746
rect 12208 2694 12220 2746
rect 12220 2694 12234 2746
rect 12258 2694 12272 2746
rect 12272 2694 12284 2746
rect 12284 2694 12314 2746
rect 12338 2694 12348 2746
rect 12348 2694 12394 2746
rect 12098 2692 12154 2694
rect 12178 2692 12234 2694
rect 12258 2692 12314 2694
rect 12338 2692 12394 2694
rect 12758 2202 12814 2204
rect 12838 2202 12894 2204
rect 12918 2202 12974 2204
rect 12998 2202 13054 2204
rect 12758 2150 12804 2202
rect 12804 2150 12814 2202
rect 12838 2150 12868 2202
rect 12868 2150 12880 2202
rect 12880 2150 12894 2202
rect 12918 2150 12932 2202
rect 12932 2150 12944 2202
rect 12944 2150 12974 2202
rect 12998 2150 13008 2202
rect 13008 2150 13054 2202
rect 12758 2148 12814 2150
rect 12838 2148 12894 2150
rect 12918 2148 12974 2150
rect 12998 2148 13054 2150
rect 19526 19066 19582 19068
rect 19606 19066 19662 19068
rect 19686 19066 19742 19068
rect 19766 19066 19822 19068
rect 19526 19014 19572 19066
rect 19572 19014 19582 19066
rect 19606 19014 19636 19066
rect 19636 19014 19648 19066
rect 19648 19014 19662 19066
rect 19686 19014 19700 19066
rect 19700 19014 19712 19066
rect 19712 19014 19742 19066
rect 19766 19014 19776 19066
rect 19776 19014 19822 19066
rect 19526 19012 19582 19014
rect 19606 19012 19662 19014
rect 19686 19012 19742 19014
rect 19766 19012 19822 19014
rect 19526 17978 19582 17980
rect 19606 17978 19662 17980
rect 19686 17978 19742 17980
rect 19766 17978 19822 17980
rect 19526 17926 19572 17978
rect 19572 17926 19582 17978
rect 19606 17926 19636 17978
rect 19636 17926 19648 17978
rect 19648 17926 19662 17978
rect 19686 17926 19700 17978
rect 19700 17926 19712 17978
rect 19712 17926 19742 17978
rect 19766 17926 19776 17978
rect 19776 17926 19822 17978
rect 19526 17924 19582 17926
rect 19606 17924 19662 17926
rect 19686 17924 19742 17926
rect 19766 17924 19822 17926
rect 19526 16890 19582 16892
rect 19606 16890 19662 16892
rect 19686 16890 19742 16892
rect 19766 16890 19822 16892
rect 19526 16838 19572 16890
rect 19572 16838 19582 16890
rect 19606 16838 19636 16890
rect 19636 16838 19648 16890
rect 19648 16838 19662 16890
rect 19686 16838 19700 16890
rect 19700 16838 19712 16890
rect 19712 16838 19742 16890
rect 19766 16838 19776 16890
rect 19776 16838 19822 16890
rect 19526 16836 19582 16838
rect 19606 16836 19662 16838
rect 19686 16836 19742 16838
rect 19766 16836 19822 16838
rect 20186 20698 20242 20700
rect 20266 20698 20322 20700
rect 20346 20698 20402 20700
rect 20426 20698 20482 20700
rect 20186 20646 20232 20698
rect 20232 20646 20242 20698
rect 20266 20646 20296 20698
rect 20296 20646 20308 20698
rect 20308 20646 20322 20698
rect 20346 20646 20360 20698
rect 20360 20646 20372 20698
rect 20372 20646 20402 20698
rect 20426 20646 20436 20698
rect 20436 20646 20482 20698
rect 20186 20644 20242 20646
rect 20266 20644 20322 20646
rect 20346 20644 20402 20646
rect 20426 20644 20482 20646
rect 20186 19610 20242 19612
rect 20266 19610 20322 19612
rect 20346 19610 20402 19612
rect 20426 19610 20482 19612
rect 20186 19558 20232 19610
rect 20232 19558 20242 19610
rect 20266 19558 20296 19610
rect 20296 19558 20308 19610
rect 20308 19558 20322 19610
rect 20346 19558 20360 19610
rect 20360 19558 20372 19610
rect 20372 19558 20402 19610
rect 20426 19558 20436 19610
rect 20436 19558 20482 19610
rect 20186 19556 20242 19558
rect 20266 19556 20322 19558
rect 20346 19556 20402 19558
rect 20426 19556 20482 19558
rect 20186 18522 20242 18524
rect 20266 18522 20322 18524
rect 20346 18522 20402 18524
rect 20426 18522 20482 18524
rect 20186 18470 20232 18522
rect 20232 18470 20242 18522
rect 20266 18470 20296 18522
rect 20296 18470 20308 18522
rect 20308 18470 20322 18522
rect 20346 18470 20360 18522
rect 20360 18470 20372 18522
rect 20372 18470 20402 18522
rect 20426 18470 20436 18522
rect 20436 18470 20482 18522
rect 20186 18468 20242 18470
rect 20266 18468 20322 18470
rect 20346 18468 20402 18470
rect 20426 18468 20482 18470
rect 20186 17434 20242 17436
rect 20266 17434 20322 17436
rect 20346 17434 20402 17436
rect 20426 17434 20482 17436
rect 20186 17382 20232 17434
rect 20232 17382 20242 17434
rect 20266 17382 20296 17434
rect 20296 17382 20308 17434
rect 20308 17382 20322 17434
rect 20346 17382 20360 17434
rect 20360 17382 20372 17434
rect 20372 17382 20402 17434
rect 20426 17382 20436 17434
rect 20436 17382 20482 17434
rect 20186 17380 20242 17382
rect 20266 17380 20322 17382
rect 20346 17380 20402 17382
rect 20426 17380 20482 17382
rect 19526 15802 19582 15804
rect 19606 15802 19662 15804
rect 19686 15802 19742 15804
rect 19766 15802 19822 15804
rect 19526 15750 19572 15802
rect 19572 15750 19582 15802
rect 19606 15750 19636 15802
rect 19636 15750 19648 15802
rect 19648 15750 19662 15802
rect 19686 15750 19700 15802
rect 19700 15750 19712 15802
rect 19712 15750 19742 15802
rect 19766 15750 19776 15802
rect 19776 15750 19822 15802
rect 19526 15748 19582 15750
rect 19606 15748 19662 15750
rect 19686 15748 19742 15750
rect 19766 15748 19822 15750
rect 19526 14714 19582 14716
rect 19606 14714 19662 14716
rect 19686 14714 19742 14716
rect 19766 14714 19822 14716
rect 19526 14662 19572 14714
rect 19572 14662 19582 14714
rect 19606 14662 19636 14714
rect 19636 14662 19648 14714
rect 19648 14662 19662 14714
rect 19686 14662 19700 14714
rect 19700 14662 19712 14714
rect 19712 14662 19742 14714
rect 19766 14662 19776 14714
rect 19776 14662 19822 14714
rect 19526 14660 19582 14662
rect 19606 14660 19662 14662
rect 19686 14660 19742 14662
rect 19766 14660 19822 14662
rect 19526 13626 19582 13628
rect 19606 13626 19662 13628
rect 19686 13626 19742 13628
rect 19766 13626 19822 13628
rect 19526 13574 19572 13626
rect 19572 13574 19582 13626
rect 19606 13574 19636 13626
rect 19636 13574 19648 13626
rect 19648 13574 19662 13626
rect 19686 13574 19700 13626
rect 19700 13574 19712 13626
rect 19712 13574 19742 13626
rect 19766 13574 19776 13626
rect 19776 13574 19822 13626
rect 19526 13572 19582 13574
rect 19606 13572 19662 13574
rect 19686 13572 19742 13574
rect 19766 13572 19822 13574
rect 20186 16346 20242 16348
rect 20266 16346 20322 16348
rect 20346 16346 20402 16348
rect 20426 16346 20482 16348
rect 20186 16294 20232 16346
rect 20232 16294 20242 16346
rect 20266 16294 20296 16346
rect 20296 16294 20308 16346
rect 20308 16294 20322 16346
rect 20346 16294 20360 16346
rect 20360 16294 20372 16346
rect 20372 16294 20402 16346
rect 20426 16294 20436 16346
rect 20436 16294 20482 16346
rect 20186 16292 20242 16294
rect 20266 16292 20322 16294
rect 20346 16292 20402 16294
rect 20426 16292 20482 16294
rect 20186 15258 20242 15260
rect 20266 15258 20322 15260
rect 20346 15258 20402 15260
rect 20426 15258 20482 15260
rect 20186 15206 20232 15258
rect 20232 15206 20242 15258
rect 20266 15206 20296 15258
rect 20296 15206 20308 15258
rect 20308 15206 20322 15258
rect 20346 15206 20360 15258
rect 20360 15206 20372 15258
rect 20372 15206 20402 15258
rect 20426 15206 20436 15258
rect 20436 15206 20482 15258
rect 20186 15204 20242 15206
rect 20266 15204 20322 15206
rect 20346 15204 20402 15206
rect 20426 15204 20482 15206
rect 20186 14170 20242 14172
rect 20266 14170 20322 14172
rect 20346 14170 20402 14172
rect 20426 14170 20482 14172
rect 20186 14118 20232 14170
rect 20232 14118 20242 14170
rect 20266 14118 20296 14170
rect 20296 14118 20308 14170
rect 20308 14118 20322 14170
rect 20346 14118 20360 14170
rect 20360 14118 20372 14170
rect 20372 14118 20402 14170
rect 20426 14118 20436 14170
rect 20436 14118 20482 14170
rect 20186 14116 20242 14118
rect 20266 14116 20322 14118
rect 20346 14116 20402 14118
rect 20426 14116 20482 14118
rect 26954 23418 27010 23420
rect 27034 23418 27090 23420
rect 27114 23418 27170 23420
rect 27194 23418 27250 23420
rect 26954 23366 27000 23418
rect 27000 23366 27010 23418
rect 27034 23366 27064 23418
rect 27064 23366 27076 23418
rect 27076 23366 27090 23418
rect 27114 23366 27128 23418
rect 27128 23366 27140 23418
rect 27140 23366 27170 23418
rect 27194 23366 27204 23418
rect 27204 23366 27250 23418
rect 26954 23364 27010 23366
rect 27034 23364 27090 23366
rect 27114 23364 27170 23366
rect 27194 23364 27250 23366
rect 20186 13082 20242 13084
rect 20266 13082 20322 13084
rect 20346 13082 20402 13084
rect 20426 13082 20482 13084
rect 20186 13030 20232 13082
rect 20232 13030 20242 13082
rect 20266 13030 20296 13082
rect 20296 13030 20308 13082
rect 20308 13030 20322 13082
rect 20346 13030 20360 13082
rect 20360 13030 20372 13082
rect 20372 13030 20402 13082
rect 20426 13030 20436 13082
rect 20436 13030 20482 13082
rect 20186 13028 20242 13030
rect 20266 13028 20322 13030
rect 20346 13028 20402 13030
rect 20426 13028 20482 13030
rect 19526 12538 19582 12540
rect 19606 12538 19662 12540
rect 19686 12538 19742 12540
rect 19766 12538 19822 12540
rect 19526 12486 19572 12538
rect 19572 12486 19582 12538
rect 19606 12486 19636 12538
rect 19636 12486 19648 12538
rect 19648 12486 19662 12538
rect 19686 12486 19700 12538
rect 19700 12486 19712 12538
rect 19712 12486 19742 12538
rect 19766 12486 19776 12538
rect 19776 12486 19822 12538
rect 19526 12484 19582 12486
rect 19606 12484 19662 12486
rect 19686 12484 19742 12486
rect 19766 12484 19822 12486
rect 20186 11994 20242 11996
rect 20266 11994 20322 11996
rect 20346 11994 20402 11996
rect 20426 11994 20482 11996
rect 20186 11942 20232 11994
rect 20232 11942 20242 11994
rect 20266 11942 20296 11994
rect 20296 11942 20308 11994
rect 20308 11942 20322 11994
rect 20346 11942 20360 11994
rect 20360 11942 20372 11994
rect 20372 11942 20402 11994
rect 20426 11942 20436 11994
rect 20436 11942 20482 11994
rect 20186 11940 20242 11942
rect 20266 11940 20322 11942
rect 20346 11940 20402 11942
rect 20426 11940 20482 11942
rect 19526 11450 19582 11452
rect 19606 11450 19662 11452
rect 19686 11450 19742 11452
rect 19766 11450 19822 11452
rect 19526 11398 19572 11450
rect 19572 11398 19582 11450
rect 19606 11398 19636 11450
rect 19636 11398 19648 11450
rect 19648 11398 19662 11450
rect 19686 11398 19700 11450
rect 19700 11398 19712 11450
rect 19712 11398 19742 11450
rect 19766 11398 19776 11450
rect 19776 11398 19822 11450
rect 19526 11396 19582 11398
rect 19606 11396 19662 11398
rect 19686 11396 19742 11398
rect 19766 11396 19822 11398
rect 19526 10362 19582 10364
rect 19606 10362 19662 10364
rect 19686 10362 19742 10364
rect 19766 10362 19822 10364
rect 19526 10310 19572 10362
rect 19572 10310 19582 10362
rect 19606 10310 19636 10362
rect 19636 10310 19648 10362
rect 19648 10310 19662 10362
rect 19686 10310 19700 10362
rect 19700 10310 19712 10362
rect 19712 10310 19742 10362
rect 19766 10310 19776 10362
rect 19776 10310 19822 10362
rect 19526 10308 19582 10310
rect 19606 10308 19662 10310
rect 19686 10308 19742 10310
rect 19766 10308 19822 10310
rect 19526 9274 19582 9276
rect 19606 9274 19662 9276
rect 19686 9274 19742 9276
rect 19766 9274 19822 9276
rect 19526 9222 19572 9274
rect 19572 9222 19582 9274
rect 19606 9222 19636 9274
rect 19636 9222 19648 9274
rect 19648 9222 19662 9274
rect 19686 9222 19700 9274
rect 19700 9222 19712 9274
rect 19712 9222 19742 9274
rect 19766 9222 19776 9274
rect 19776 9222 19822 9274
rect 19526 9220 19582 9222
rect 19606 9220 19662 9222
rect 19686 9220 19742 9222
rect 19766 9220 19822 9222
rect 19526 8186 19582 8188
rect 19606 8186 19662 8188
rect 19686 8186 19742 8188
rect 19766 8186 19822 8188
rect 19526 8134 19572 8186
rect 19572 8134 19582 8186
rect 19606 8134 19636 8186
rect 19636 8134 19648 8186
rect 19648 8134 19662 8186
rect 19686 8134 19700 8186
rect 19700 8134 19712 8186
rect 19712 8134 19742 8186
rect 19766 8134 19776 8186
rect 19776 8134 19822 8186
rect 19526 8132 19582 8134
rect 19606 8132 19662 8134
rect 19686 8132 19742 8134
rect 19766 8132 19822 8134
rect 20186 10906 20242 10908
rect 20266 10906 20322 10908
rect 20346 10906 20402 10908
rect 20426 10906 20482 10908
rect 20186 10854 20232 10906
rect 20232 10854 20242 10906
rect 20266 10854 20296 10906
rect 20296 10854 20308 10906
rect 20308 10854 20322 10906
rect 20346 10854 20360 10906
rect 20360 10854 20372 10906
rect 20372 10854 20402 10906
rect 20426 10854 20436 10906
rect 20436 10854 20482 10906
rect 20186 10852 20242 10854
rect 20266 10852 20322 10854
rect 20346 10852 20402 10854
rect 20426 10852 20482 10854
rect 21822 11076 21878 11112
rect 21822 11056 21824 11076
rect 21824 11056 21876 11076
rect 21876 11056 21878 11076
rect 20186 9818 20242 9820
rect 20266 9818 20322 9820
rect 20346 9818 20402 9820
rect 20426 9818 20482 9820
rect 20186 9766 20232 9818
rect 20232 9766 20242 9818
rect 20266 9766 20296 9818
rect 20296 9766 20308 9818
rect 20308 9766 20322 9818
rect 20346 9766 20360 9818
rect 20360 9766 20372 9818
rect 20372 9766 20402 9818
rect 20426 9766 20436 9818
rect 20436 9766 20482 9818
rect 20186 9764 20242 9766
rect 20266 9764 20322 9766
rect 20346 9764 20402 9766
rect 20426 9764 20482 9766
rect 20186 8730 20242 8732
rect 20266 8730 20322 8732
rect 20346 8730 20402 8732
rect 20426 8730 20482 8732
rect 20186 8678 20232 8730
rect 20232 8678 20242 8730
rect 20266 8678 20296 8730
rect 20296 8678 20308 8730
rect 20308 8678 20322 8730
rect 20346 8678 20360 8730
rect 20360 8678 20372 8730
rect 20372 8678 20402 8730
rect 20426 8678 20436 8730
rect 20436 8678 20482 8730
rect 20186 8676 20242 8678
rect 20266 8676 20322 8678
rect 20346 8676 20402 8678
rect 20426 8676 20482 8678
rect 19526 7098 19582 7100
rect 19606 7098 19662 7100
rect 19686 7098 19742 7100
rect 19766 7098 19822 7100
rect 19526 7046 19572 7098
rect 19572 7046 19582 7098
rect 19606 7046 19636 7098
rect 19636 7046 19648 7098
rect 19648 7046 19662 7098
rect 19686 7046 19700 7098
rect 19700 7046 19712 7098
rect 19712 7046 19742 7098
rect 19766 7046 19776 7098
rect 19776 7046 19822 7098
rect 19526 7044 19582 7046
rect 19606 7044 19662 7046
rect 19686 7044 19742 7046
rect 19766 7044 19822 7046
rect 19526 6010 19582 6012
rect 19606 6010 19662 6012
rect 19686 6010 19742 6012
rect 19766 6010 19822 6012
rect 19526 5958 19572 6010
rect 19572 5958 19582 6010
rect 19606 5958 19636 6010
rect 19636 5958 19648 6010
rect 19648 5958 19662 6010
rect 19686 5958 19700 6010
rect 19700 5958 19712 6010
rect 19712 5958 19742 6010
rect 19766 5958 19776 6010
rect 19776 5958 19822 6010
rect 19526 5956 19582 5958
rect 19606 5956 19662 5958
rect 19686 5956 19742 5958
rect 19766 5956 19822 5958
rect 19526 4922 19582 4924
rect 19606 4922 19662 4924
rect 19686 4922 19742 4924
rect 19766 4922 19822 4924
rect 19526 4870 19572 4922
rect 19572 4870 19582 4922
rect 19606 4870 19636 4922
rect 19636 4870 19648 4922
rect 19648 4870 19662 4922
rect 19686 4870 19700 4922
rect 19700 4870 19712 4922
rect 19712 4870 19742 4922
rect 19766 4870 19776 4922
rect 19776 4870 19822 4922
rect 19526 4868 19582 4870
rect 19606 4868 19662 4870
rect 19686 4868 19742 4870
rect 19766 4868 19822 4870
rect 19526 3834 19582 3836
rect 19606 3834 19662 3836
rect 19686 3834 19742 3836
rect 19766 3834 19822 3836
rect 19526 3782 19572 3834
rect 19572 3782 19582 3834
rect 19606 3782 19636 3834
rect 19636 3782 19648 3834
rect 19648 3782 19662 3834
rect 19686 3782 19700 3834
rect 19700 3782 19712 3834
rect 19712 3782 19742 3834
rect 19766 3782 19776 3834
rect 19776 3782 19822 3834
rect 19526 3780 19582 3782
rect 19606 3780 19662 3782
rect 19686 3780 19742 3782
rect 19766 3780 19822 3782
rect 19526 2746 19582 2748
rect 19606 2746 19662 2748
rect 19686 2746 19742 2748
rect 19766 2746 19822 2748
rect 19526 2694 19572 2746
rect 19572 2694 19582 2746
rect 19606 2694 19636 2746
rect 19636 2694 19648 2746
rect 19648 2694 19662 2746
rect 19686 2694 19700 2746
rect 19700 2694 19712 2746
rect 19712 2694 19742 2746
rect 19766 2694 19776 2746
rect 19776 2694 19822 2746
rect 19526 2692 19582 2694
rect 19606 2692 19662 2694
rect 19686 2692 19742 2694
rect 19766 2692 19822 2694
rect 20186 7642 20242 7644
rect 20266 7642 20322 7644
rect 20346 7642 20402 7644
rect 20426 7642 20482 7644
rect 20186 7590 20232 7642
rect 20232 7590 20242 7642
rect 20266 7590 20296 7642
rect 20296 7590 20308 7642
rect 20308 7590 20322 7642
rect 20346 7590 20360 7642
rect 20360 7590 20372 7642
rect 20372 7590 20402 7642
rect 20426 7590 20436 7642
rect 20436 7590 20482 7642
rect 20186 7588 20242 7590
rect 20266 7588 20322 7590
rect 20346 7588 20402 7590
rect 20426 7588 20482 7590
rect 26954 22330 27010 22332
rect 27034 22330 27090 22332
rect 27114 22330 27170 22332
rect 27194 22330 27250 22332
rect 26954 22278 27000 22330
rect 27000 22278 27010 22330
rect 27034 22278 27064 22330
rect 27064 22278 27076 22330
rect 27076 22278 27090 22330
rect 27114 22278 27128 22330
rect 27128 22278 27140 22330
rect 27140 22278 27170 22330
rect 27194 22278 27204 22330
rect 27204 22278 27250 22330
rect 26954 22276 27010 22278
rect 27034 22276 27090 22278
rect 27114 22276 27170 22278
rect 27194 22276 27250 22278
rect 27614 22874 27670 22876
rect 27694 22874 27750 22876
rect 27774 22874 27830 22876
rect 27854 22874 27910 22876
rect 27614 22822 27660 22874
rect 27660 22822 27670 22874
rect 27694 22822 27724 22874
rect 27724 22822 27736 22874
rect 27736 22822 27750 22874
rect 27774 22822 27788 22874
rect 27788 22822 27800 22874
rect 27800 22822 27830 22874
rect 27854 22822 27864 22874
rect 27864 22822 27910 22874
rect 27614 22820 27670 22822
rect 27694 22820 27750 22822
rect 27774 22820 27830 22822
rect 27854 22820 27910 22822
rect 26330 21972 26332 21992
rect 26332 21972 26384 21992
rect 26384 21972 26386 21992
rect 26330 21936 26386 21972
rect 25870 20984 25926 21040
rect 26954 21242 27010 21244
rect 27034 21242 27090 21244
rect 27114 21242 27170 21244
rect 27194 21242 27250 21244
rect 26954 21190 27000 21242
rect 27000 21190 27010 21242
rect 27034 21190 27064 21242
rect 27064 21190 27076 21242
rect 27076 21190 27090 21242
rect 27114 21190 27128 21242
rect 27128 21190 27140 21242
rect 27140 21190 27170 21242
rect 27194 21190 27204 21242
rect 27204 21190 27250 21242
rect 26954 21188 27010 21190
rect 27034 21188 27090 21190
rect 27114 21188 27170 21190
rect 27194 21188 27250 21190
rect 27158 21004 27214 21040
rect 27158 20984 27160 21004
rect 27160 20984 27212 21004
rect 27212 20984 27214 21004
rect 27614 21786 27670 21788
rect 27694 21786 27750 21788
rect 27774 21786 27830 21788
rect 27854 21786 27910 21788
rect 27614 21734 27660 21786
rect 27660 21734 27670 21786
rect 27694 21734 27724 21786
rect 27724 21734 27736 21786
rect 27736 21734 27750 21786
rect 27774 21734 27788 21786
rect 27788 21734 27800 21786
rect 27800 21734 27830 21786
rect 27854 21734 27864 21786
rect 27864 21734 27910 21786
rect 27614 21732 27670 21734
rect 27694 21732 27750 21734
rect 27774 21732 27830 21734
rect 27854 21732 27910 21734
rect 28078 21836 28080 21856
rect 28080 21836 28132 21856
rect 28132 21836 28134 21856
rect 28078 21800 28134 21836
rect 27614 20698 27670 20700
rect 27694 20698 27750 20700
rect 27774 20698 27830 20700
rect 27854 20698 27910 20700
rect 27614 20646 27660 20698
rect 27660 20646 27670 20698
rect 27694 20646 27724 20698
rect 27724 20646 27736 20698
rect 27736 20646 27750 20698
rect 27774 20646 27788 20698
rect 27788 20646 27800 20698
rect 27800 20646 27830 20698
rect 27854 20646 27864 20698
rect 27864 20646 27910 20698
rect 27614 20644 27670 20646
rect 27694 20644 27750 20646
rect 27774 20644 27830 20646
rect 27854 20644 27910 20646
rect 26954 20154 27010 20156
rect 27034 20154 27090 20156
rect 27114 20154 27170 20156
rect 27194 20154 27250 20156
rect 26954 20102 27000 20154
rect 27000 20102 27010 20154
rect 27034 20102 27064 20154
rect 27064 20102 27076 20154
rect 27076 20102 27090 20154
rect 27114 20102 27128 20154
rect 27128 20102 27140 20154
rect 27140 20102 27170 20154
rect 27194 20102 27204 20154
rect 27204 20102 27250 20154
rect 26954 20100 27010 20102
rect 27034 20100 27090 20102
rect 27114 20100 27170 20102
rect 27194 20100 27250 20102
rect 27618 20440 27674 20496
rect 27614 19610 27670 19612
rect 27694 19610 27750 19612
rect 27774 19610 27830 19612
rect 27854 19610 27910 19612
rect 27614 19558 27660 19610
rect 27660 19558 27670 19610
rect 27694 19558 27724 19610
rect 27724 19558 27736 19610
rect 27736 19558 27750 19610
rect 27774 19558 27788 19610
rect 27788 19558 27800 19610
rect 27800 19558 27830 19610
rect 27854 19558 27864 19610
rect 27864 19558 27910 19610
rect 27614 19556 27670 19558
rect 27694 19556 27750 19558
rect 27774 19556 27830 19558
rect 27854 19556 27910 19558
rect 26954 19066 27010 19068
rect 27034 19066 27090 19068
rect 27114 19066 27170 19068
rect 27194 19066 27250 19068
rect 26954 19014 27000 19066
rect 27000 19014 27010 19066
rect 27034 19014 27064 19066
rect 27064 19014 27076 19066
rect 27076 19014 27090 19066
rect 27114 19014 27128 19066
rect 27128 19014 27140 19066
rect 27140 19014 27170 19066
rect 27194 19014 27204 19066
rect 27204 19014 27250 19066
rect 26954 19012 27010 19014
rect 27034 19012 27090 19014
rect 27114 19012 27170 19014
rect 27194 19012 27250 19014
rect 26954 17978 27010 17980
rect 27034 17978 27090 17980
rect 27114 17978 27170 17980
rect 27194 17978 27250 17980
rect 26954 17926 27000 17978
rect 27000 17926 27010 17978
rect 27034 17926 27064 17978
rect 27064 17926 27076 17978
rect 27076 17926 27090 17978
rect 27114 17926 27128 17978
rect 27128 17926 27140 17978
rect 27140 17926 27170 17978
rect 27194 17926 27204 17978
rect 27204 17926 27250 17978
rect 26954 17924 27010 17926
rect 27034 17924 27090 17926
rect 27114 17924 27170 17926
rect 27194 17924 27250 17926
rect 27614 18522 27670 18524
rect 27694 18522 27750 18524
rect 27774 18522 27830 18524
rect 27854 18522 27910 18524
rect 27614 18470 27660 18522
rect 27660 18470 27670 18522
rect 27694 18470 27724 18522
rect 27724 18470 27736 18522
rect 27736 18470 27750 18522
rect 27774 18470 27788 18522
rect 27788 18470 27800 18522
rect 27800 18470 27830 18522
rect 27854 18470 27864 18522
rect 27864 18470 27910 18522
rect 27614 18468 27670 18470
rect 27694 18468 27750 18470
rect 27774 18468 27830 18470
rect 27854 18468 27910 18470
rect 28630 19780 28686 19816
rect 28630 19760 28632 19780
rect 28632 19760 28684 19780
rect 28684 19760 28686 19780
rect 28998 20324 29054 20360
rect 28998 20304 29000 20324
rect 29000 20304 29052 20324
rect 29052 20304 29054 20324
rect 29550 20340 29552 20360
rect 29552 20340 29604 20360
rect 29604 20340 29606 20360
rect 29550 20304 29606 20340
rect 27618 17720 27674 17776
rect 27614 17434 27670 17436
rect 27694 17434 27750 17436
rect 27774 17434 27830 17436
rect 27854 17434 27910 17436
rect 27614 17382 27660 17434
rect 27660 17382 27670 17434
rect 27694 17382 27724 17434
rect 27724 17382 27736 17434
rect 27736 17382 27750 17434
rect 27774 17382 27788 17434
rect 27788 17382 27800 17434
rect 27800 17382 27830 17434
rect 27854 17382 27864 17434
rect 27864 17382 27910 17434
rect 27614 17380 27670 17382
rect 27694 17380 27750 17382
rect 27774 17380 27830 17382
rect 27854 17380 27910 17382
rect 26954 16890 27010 16892
rect 27034 16890 27090 16892
rect 27114 16890 27170 16892
rect 27194 16890 27250 16892
rect 26954 16838 27000 16890
rect 27000 16838 27010 16890
rect 27034 16838 27064 16890
rect 27064 16838 27076 16890
rect 27076 16838 27090 16890
rect 27114 16838 27128 16890
rect 27128 16838 27140 16890
rect 27140 16838 27170 16890
rect 27194 16838 27204 16890
rect 27204 16838 27250 16890
rect 26954 16836 27010 16838
rect 27034 16836 27090 16838
rect 27114 16836 27170 16838
rect 27194 16836 27250 16838
rect 27802 17060 27858 17096
rect 27802 17040 27804 17060
rect 27804 17040 27856 17060
rect 27856 17040 27858 17060
rect 27614 16346 27670 16348
rect 27694 16346 27750 16348
rect 27774 16346 27830 16348
rect 27854 16346 27910 16348
rect 27614 16294 27660 16346
rect 27660 16294 27670 16346
rect 27694 16294 27724 16346
rect 27724 16294 27736 16346
rect 27736 16294 27750 16346
rect 27774 16294 27788 16346
rect 27788 16294 27800 16346
rect 27800 16294 27830 16346
rect 27854 16294 27864 16346
rect 27864 16294 27910 16346
rect 27614 16292 27670 16294
rect 27694 16292 27750 16294
rect 27774 16292 27830 16294
rect 27854 16292 27910 16294
rect 26954 15802 27010 15804
rect 27034 15802 27090 15804
rect 27114 15802 27170 15804
rect 27194 15802 27250 15804
rect 26954 15750 27000 15802
rect 27000 15750 27010 15802
rect 27034 15750 27064 15802
rect 27064 15750 27076 15802
rect 27076 15750 27090 15802
rect 27114 15750 27128 15802
rect 27128 15750 27140 15802
rect 27140 15750 27170 15802
rect 27194 15750 27204 15802
rect 27204 15750 27250 15802
rect 26954 15748 27010 15750
rect 27034 15748 27090 15750
rect 27114 15748 27170 15750
rect 27194 15748 27250 15750
rect 27618 15680 27674 15736
rect 27614 15258 27670 15260
rect 27694 15258 27750 15260
rect 27774 15258 27830 15260
rect 27854 15258 27910 15260
rect 27614 15206 27660 15258
rect 27660 15206 27670 15258
rect 27694 15206 27724 15258
rect 27724 15206 27736 15258
rect 27736 15206 27750 15258
rect 27774 15206 27788 15258
rect 27788 15206 27800 15258
rect 27800 15206 27830 15258
rect 27854 15206 27864 15258
rect 27864 15206 27910 15258
rect 27614 15204 27670 15206
rect 27694 15204 27750 15206
rect 27774 15204 27830 15206
rect 27854 15204 27910 15206
rect 26954 14714 27010 14716
rect 27034 14714 27090 14716
rect 27114 14714 27170 14716
rect 27194 14714 27250 14716
rect 26954 14662 27000 14714
rect 27000 14662 27010 14714
rect 27034 14662 27064 14714
rect 27064 14662 27076 14714
rect 27076 14662 27090 14714
rect 27114 14662 27128 14714
rect 27128 14662 27140 14714
rect 27140 14662 27170 14714
rect 27194 14662 27204 14714
rect 27204 14662 27250 14714
rect 26954 14660 27010 14662
rect 27034 14660 27090 14662
rect 27114 14660 27170 14662
rect 27194 14660 27250 14662
rect 27614 14170 27670 14172
rect 27694 14170 27750 14172
rect 27774 14170 27830 14172
rect 27854 14170 27910 14172
rect 27614 14118 27660 14170
rect 27660 14118 27670 14170
rect 27694 14118 27724 14170
rect 27724 14118 27736 14170
rect 27736 14118 27750 14170
rect 27774 14118 27788 14170
rect 27788 14118 27800 14170
rect 27800 14118 27830 14170
rect 27854 14118 27864 14170
rect 27864 14118 27910 14170
rect 27614 14116 27670 14118
rect 27694 14116 27750 14118
rect 27774 14116 27830 14118
rect 27854 14116 27910 14118
rect 27342 13640 27398 13696
rect 26954 13626 27010 13628
rect 27034 13626 27090 13628
rect 27114 13626 27170 13628
rect 27194 13626 27250 13628
rect 26954 13574 27000 13626
rect 27000 13574 27010 13626
rect 27034 13574 27064 13626
rect 27064 13574 27076 13626
rect 27076 13574 27090 13626
rect 27114 13574 27128 13626
rect 27128 13574 27140 13626
rect 27140 13574 27170 13626
rect 27194 13574 27204 13626
rect 27204 13574 27250 13626
rect 26954 13572 27010 13574
rect 27034 13572 27090 13574
rect 27114 13572 27170 13574
rect 27194 13572 27250 13574
rect 28630 18400 28686 18456
rect 30378 16360 30434 16416
rect 20186 6554 20242 6556
rect 20266 6554 20322 6556
rect 20346 6554 20402 6556
rect 20426 6554 20482 6556
rect 20186 6502 20232 6554
rect 20232 6502 20242 6554
rect 20266 6502 20296 6554
rect 20296 6502 20308 6554
rect 20308 6502 20322 6554
rect 20346 6502 20360 6554
rect 20360 6502 20372 6554
rect 20372 6502 20402 6554
rect 20426 6502 20436 6554
rect 20436 6502 20482 6554
rect 20186 6500 20242 6502
rect 20266 6500 20322 6502
rect 20346 6500 20402 6502
rect 20426 6500 20482 6502
rect 20186 5466 20242 5468
rect 20266 5466 20322 5468
rect 20346 5466 20402 5468
rect 20426 5466 20482 5468
rect 20186 5414 20232 5466
rect 20232 5414 20242 5466
rect 20266 5414 20296 5466
rect 20296 5414 20308 5466
rect 20308 5414 20322 5466
rect 20346 5414 20360 5466
rect 20360 5414 20372 5466
rect 20372 5414 20402 5466
rect 20426 5414 20436 5466
rect 20436 5414 20482 5466
rect 20186 5412 20242 5414
rect 20266 5412 20322 5414
rect 20346 5412 20402 5414
rect 20426 5412 20482 5414
rect 20186 4378 20242 4380
rect 20266 4378 20322 4380
rect 20346 4378 20402 4380
rect 20426 4378 20482 4380
rect 20186 4326 20232 4378
rect 20232 4326 20242 4378
rect 20266 4326 20296 4378
rect 20296 4326 20308 4378
rect 20308 4326 20322 4378
rect 20346 4326 20360 4378
rect 20360 4326 20372 4378
rect 20372 4326 20402 4378
rect 20426 4326 20436 4378
rect 20436 4326 20482 4378
rect 20186 4324 20242 4326
rect 20266 4324 20322 4326
rect 20346 4324 20402 4326
rect 20426 4324 20482 4326
rect 20186 3290 20242 3292
rect 20266 3290 20322 3292
rect 20346 3290 20402 3292
rect 20426 3290 20482 3292
rect 20186 3238 20232 3290
rect 20232 3238 20242 3290
rect 20266 3238 20296 3290
rect 20296 3238 20308 3290
rect 20308 3238 20322 3290
rect 20346 3238 20360 3290
rect 20360 3238 20372 3290
rect 20372 3238 20402 3290
rect 20426 3238 20436 3290
rect 20436 3238 20482 3290
rect 20186 3236 20242 3238
rect 20266 3236 20322 3238
rect 20346 3236 20402 3238
rect 20426 3236 20482 3238
rect 20186 2202 20242 2204
rect 20266 2202 20322 2204
rect 20346 2202 20402 2204
rect 20426 2202 20482 2204
rect 20186 2150 20232 2202
rect 20232 2150 20242 2202
rect 20266 2150 20296 2202
rect 20296 2150 20308 2202
rect 20308 2150 20322 2202
rect 20346 2150 20360 2202
rect 20360 2150 20372 2202
rect 20372 2150 20402 2202
rect 20426 2150 20436 2202
rect 20436 2150 20482 2202
rect 20186 2148 20242 2150
rect 20266 2148 20322 2150
rect 20346 2148 20402 2150
rect 20426 2148 20482 2150
rect 27614 13082 27670 13084
rect 27694 13082 27750 13084
rect 27774 13082 27830 13084
rect 27854 13082 27910 13084
rect 27614 13030 27660 13082
rect 27660 13030 27670 13082
rect 27694 13030 27724 13082
rect 27724 13030 27736 13082
rect 27736 13030 27750 13082
rect 27774 13030 27788 13082
rect 27788 13030 27800 13082
rect 27800 13030 27830 13082
rect 27854 13030 27864 13082
rect 27864 13030 27910 13082
rect 27614 13028 27670 13030
rect 27694 13028 27750 13030
rect 27774 13028 27830 13030
rect 27854 13028 27910 13030
rect 26954 12538 27010 12540
rect 27034 12538 27090 12540
rect 27114 12538 27170 12540
rect 27194 12538 27250 12540
rect 26954 12486 27000 12538
rect 27000 12486 27010 12538
rect 27034 12486 27064 12538
rect 27064 12486 27076 12538
rect 27076 12486 27090 12538
rect 27114 12486 27128 12538
rect 27128 12486 27140 12538
rect 27140 12486 27170 12538
rect 27194 12486 27204 12538
rect 27204 12486 27250 12538
rect 26954 12484 27010 12486
rect 27034 12484 27090 12486
rect 27114 12484 27170 12486
rect 27194 12484 27250 12486
rect 27614 11994 27670 11996
rect 27694 11994 27750 11996
rect 27774 11994 27830 11996
rect 27854 11994 27910 11996
rect 27614 11942 27660 11994
rect 27660 11942 27670 11994
rect 27694 11942 27724 11994
rect 27724 11942 27736 11994
rect 27736 11942 27750 11994
rect 27774 11942 27788 11994
rect 27788 11942 27800 11994
rect 27800 11942 27830 11994
rect 27854 11942 27864 11994
rect 27864 11942 27910 11994
rect 27614 11940 27670 11942
rect 27694 11940 27750 11942
rect 27774 11940 27830 11942
rect 27854 11940 27910 11942
rect 26954 11450 27010 11452
rect 27034 11450 27090 11452
rect 27114 11450 27170 11452
rect 27194 11450 27250 11452
rect 26954 11398 27000 11450
rect 27000 11398 27010 11450
rect 27034 11398 27064 11450
rect 27064 11398 27076 11450
rect 27076 11398 27090 11450
rect 27114 11398 27128 11450
rect 27128 11398 27140 11450
rect 27140 11398 27170 11450
rect 27194 11398 27204 11450
rect 27204 11398 27250 11450
rect 26954 11396 27010 11398
rect 27034 11396 27090 11398
rect 27114 11396 27170 11398
rect 27194 11396 27250 11398
rect 27614 10906 27670 10908
rect 27694 10906 27750 10908
rect 27774 10906 27830 10908
rect 27854 10906 27910 10908
rect 27614 10854 27660 10906
rect 27660 10854 27670 10906
rect 27694 10854 27724 10906
rect 27724 10854 27736 10906
rect 27736 10854 27750 10906
rect 27774 10854 27788 10906
rect 27788 10854 27800 10906
rect 27800 10854 27830 10906
rect 27854 10854 27864 10906
rect 27864 10854 27910 10906
rect 27614 10852 27670 10854
rect 27694 10852 27750 10854
rect 27774 10852 27830 10854
rect 27854 10852 27910 10854
rect 26954 10362 27010 10364
rect 27034 10362 27090 10364
rect 27114 10362 27170 10364
rect 27194 10362 27250 10364
rect 26954 10310 27000 10362
rect 27000 10310 27010 10362
rect 27034 10310 27064 10362
rect 27064 10310 27076 10362
rect 27076 10310 27090 10362
rect 27114 10310 27128 10362
rect 27128 10310 27140 10362
rect 27140 10310 27170 10362
rect 27194 10310 27204 10362
rect 27204 10310 27250 10362
rect 26954 10308 27010 10310
rect 27034 10308 27090 10310
rect 27114 10308 27170 10310
rect 27194 10308 27250 10310
rect 27614 9818 27670 9820
rect 27694 9818 27750 9820
rect 27774 9818 27830 9820
rect 27854 9818 27910 9820
rect 27614 9766 27660 9818
rect 27660 9766 27670 9818
rect 27694 9766 27724 9818
rect 27724 9766 27736 9818
rect 27736 9766 27750 9818
rect 27774 9766 27788 9818
rect 27788 9766 27800 9818
rect 27800 9766 27830 9818
rect 27854 9766 27864 9818
rect 27864 9766 27910 9818
rect 27614 9764 27670 9766
rect 27694 9764 27750 9766
rect 27774 9764 27830 9766
rect 27854 9764 27910 9766
rect 26954 9274 27010 9276
rect 27034 9274 27090 9276
rect 27114 9274 27170 9276
rect 27194 9274 27250 9276
rect 26954 9222 27000 9274
rect 27000 9222 27010 9274
rect 27034 9222 27064 9274
rect 27064 9222 27076 9274
rect 27076 9222 27090 9274
rect 27114 9222 27128 9274
rect 27128 9222 27140 9274
rect 27140 9222 27170 9274
rect 27194 9222 27204 9274
rect 27204 9222 27250 9274
rect 26954 9220 27010 9222
rect 27034 9220 27090 9222
rect 27114 9220 27170 9222
rect 27194 9220 27250 9222
rect 27614 8730 27670 8732
rect 27694 8730 27750 8732
rect 27774 8730 27830 8732
rect 27854 8730 27910 8732
rect 27614 8678 27660 8730
rect 27660 8678 27670 8730
rect 27694 8678 27724 8730
rect 27724 8678 27736 8730
rect 27736 8678 27750 8730
rect 27774 8678 27788 8730
rect 27788 8678 27800 8730
rect 27800 8678 27830 8730
rect 27854 8678 27864 8730
rect 27864 8678 27910 8730
rect 27614 8676 27670 8678
rect 27694 8676 27750 8678
rect 27774 8676 27830 8678
rect 27854 8676 27910 8678
rect 26954 8186 27010 8188
rect 27034 8186 27090 8188
rect 27114 8186 27170 8188
rect 27194 8186 27250 8188
rect 26954 8134 27000 8186
rect 27000 8134 27010 8186
rect 27034 8134 27064 8186
rect 27064 8134 27076 8186
rect 27076 8134 27090 8186
rect 27114 8134 27128 8186
rect 27128 8134 27140 8186
rect 27140 8134 27170 8186
rect 27194 8134 27204 8186
rect 27204 8134 27250 8186
rect 26954 8132 27010 8134
rect 27034 8132 27090 8134
rect 27114 8132 27170 8134
rect 27194 8132 27250 8134
rect 27614 7642 27670 7644
rect 27694 7642 27750 7644
rect 27774 7642 27830 7644
rect 27854 7642 27910 7644
rect 27614 7590 27660 7642
rect 27660 7590 27670 7642
rect 27694 7590 27724 7642
rect 27724 7590 27736 7642
rect 27736 7590 27750 7642
rect 27774 7590 27788 7642
rect 27788 7590 27800 7642
rect 27800 7590 27830 7642
rect 27854 7590 27864 7642
rect 27864 7590 27910 7642
rect 27614 7588 27670 7590
rect 27694 7588 27750 7590
rect 27774 7588 27830 7590
rect 27854 7588 27910 7590
rect 26954 7098 27010 7100
rect 27034 7098 27090 7100
rect 27114 7098 27170 7100
rect 27194 7098 27250 7100
rect 26954 7046 27000 7098
rect 27000 7046 27010 7098
rect 27034 7046 27064 7098
rect 27064 7046 27076 7098
rect 27076 7046 27090 7098
rect 27114 7046 27128 7098
rect 27128 7046 27140 7098
rect 27140 7046 27170 7098
rect 27194 7046 27204 7098
rect 27204 7046 27250 7098
rect 26954 7044 27010 7046
rect 27034 7044 27090 7046
rect 27114 7044 27170 7046
rect 27194 7044 27250 7046
rect 27614 6554 27670 6556
rect 27694 6554 27750 6556
rect 27774 6554 27830 6556
rect 27854 6554 27910 6556
rect 27614 6502 27660 6554
rect 27660 6502 27670 6554
rect 27694 6502 27724 6554
rect 27724 6502 27736 6554
rect 27736 6502 27750 6554
rect 27774 6502 27788 6554
rect 27788 6502 27800 6554
rect 27800 6502 27830 6554
rect 27854 6502 27864 6554
rect 27864 6502 27910 6554
rect 27614 6500 27670 6502
rect 27694 6500 27750 6502
rect 27774 6500 27830 6502
rect 27854 6500 27910 6502
rect 26954 6010 27010 6012
rect 27034 6010 27090 6012
rect 27114 6010 27170 6012
rect 27194 6010 27250 6012
rect 26954 5958 27000 6010
rect 27000 5958 27010 6010
rect 27034 5958 27064 6010
rect 27064 5958 27076 6010
rect 27076 5958 27090 6010
rect 27114 5958 27128 6010
rect 27128 5958 27140 6010
rect 27140 5958 27170 6010
rect 27194 5958 27204 6010
rect 27204 5958 27250 6010
rect 26954 5956 27010 5958
rect 27034 5956 27090 5958
rect 27114 5956 27170 5958
rect 27194 5956 27250 5958
rect 27614 5466 27670 5468
rect 27694 5466 27750 5468
rect 27774 5466 27830 5468
rect 27854 5466 27910 5468
rect 27614 5414 27660 5466
rect 27660 5414 27670 5466
rect 27694 5414 27724 5466
rect 27724 5414 27736 5466
rect 27736 5414 27750 5466
rect 27774 5414 27788 5466
rect 27788 5414 27800 5466
rect 27800 5414 27830 5466
rect 27854 5414 27864 5466
rect 27864 5414 27910 5466
rect 27614 5412 27670 5414
rect 27694 5412 27750 5414
rect 27774 5412 27830 5414
rect 27854 5412 27910 5414
rect 26954 4922 27010 4924
rect 27034 4922 27090 4924
rect 27114 4922 27170 4924
rect 27194 4922 27250 4924
rect 26954 4870 27000 4922
rect 27000 4870 27010 4922
rect 27034 4870 27064 4922
rect 27064 4870 27076 4922
rect 27076 4870 27090 4922
rect 27114 4870 27128 4922
rect 27128 4870 27140 4922
rect 27140 4870 27170 4922
rect 27194 4870 27204 4922
rect 27204 4870 27250 4922
rect 26954 4868 27010 4870
rect 27034 4868 27090 4870
rect 27114 4868 27170 4870
rect 27194 4868 27250 4870
rect 27614 4378 27670 4380
rect 27694 4378 27750 4380
rect 27774 4378 27830 4380
rect 27854 4378 27910 4380
rect 27614 4326 27660 4378
rect 27660 4326 27670 4378
rect 27694 4326 27724 4378
rect 27724 4326 27736 4378
rect 27736 4326 27750 4378
rect 27774 4326 27788 4378
rect 27788 4326 27800 4378
rect 27800 4326 27830 4378
rect 27854 4326 27864 4378
rect 27864 4326 27910 4378
rect 27614 4324 27670 4326
rect 27694 4324 27750 4326
rect 27774 4324 27830 4326
rect 27854 4324 27910 4326
rect 26954 3834 27010 3836
rect 27034 3834 27090 3836
rect 27114 3834 27170 3836
rect 27194 3834 27250 3836
rect 26954 3782 27000 3834
rect 27000 3782 27010 3834
rect 27034 3782 27064 3834
rect 27064 3782 27076 3834
rect 27076 3782 27090 3834
rect 27114 3782 27128 3834
rect 27128 3782 27140 3834
rect 27140 3782 27170 3834
rect 27194 3782 27204 3834
rect 27204 3782 27250 3834
rect 26954 3780 27010 3782
rect 27034 3780 27090 3782
rect 27114 3780 27170 3782
rect 27194 3780 27250 3782
rect 27614 3290 27670 3292
rect 27694 3290 27750 3292
rect 27774 3290 27830 3292
rect 27854 3290 27910 3292
rect 27614 3238 27660 3290
rect 27660 3238 27670 3290
rect 27694 3238 27724 3290
rect 27724 3238 27736 3290
rect 27736 3238 27750 3290
rect 27774 3238 27788 3290
rect 27788 3238 27800 3290
rect 27800 3238 27830 3290
rect 27854 3238 27864 3290
rect 27864 3238 27910 3290
rect 27614 3236 27670 3238
rect 27694 3236 27750 3238
rect 27774 3236 27830 3238
rect 27854 3236 27910 3238
rect 26954 2746 27010 2748
rect 27034 2746 27090 2748
rect 27114 2746 27170 2748
rect 27194 2746 27250 2748
rect 26954 2694 27000 2746
rect 27000 2694 27010 2746
rect 27034 2694 27064 2746
rect 27064 2694 27076 2746
rect 27076 2694 27090 2746
rect 27114 2694 27128 2746
rect 27128 2694 27140 2746
rect 27140 2694 27170 2746
rect 27194 2694 27204 2746
rect 27204 2694 27250 2746
rect 26954 2692 27010 2694
rect 27034 2692 27090 2694
rect 27114 2692 27170 2694
rect 27194 2692 27250 2694
rect 27614 2202 27670 2204
rect 27694 2202 27750 2204
rect 27774 2202 27830 2204
rect 27854 2202 27910 2204
rect 27614 2150 27660 2202
rect 27660 2150 27670 2202
rect 27694 2150 27724 2202
rect 27724 2150 27736 2202
rect 27736 2150 27750 2202
rect 27774 2150 27788 2202
rect 27788 2150 27800 2202
rect 27800 2150 27830 2202
rect 27854 2150 27864 2202
rect 27864 2150 27910 2202
rect 27614 2148 27670 2150
rect 27694 2148 27750 2150
rect 27774 2148 27830 2150
rect 27854 2148 27910 2150
<< metal3 >>
rect 5320 29408 5636 29409
rect 5320 29344 5326 29408
rect 5390 29344 5406 29408
rect 5470 29344 5486 29408
rect 5550 29344 5566 29408
rect 5630 29344 5636 29408
rect 5320 29343 5636 29344
rect 12748 29408 13064 29409
rect 12748 29344 12754 29408
rect 12818 29344 12834 29408
rect 12898 29344 12914 29408
rect 12978 29344 12994 29408
rect 13058 29344 13064 29408
rect 12748 29343 13064 29344
rect 20176 29408 20492 29409
rect 20176 29344 20182 29408
rect 20246 29344 20262 29408
rect 20326 29344 20342 29408
rect 20406 29344 20422 29408
rect 20486 29344 20492 29408
rect 20176 29343 20492 29344
rect 27604 29408 27920 29409
rect 27604 29344 27610 29408
rect 27674 29344 27690 29408
rect 27754 29344 27770 29408
rect 27834 29344 27850 29408
rect 27914 29344 27920 29408
rect 27604 29343 27920 29344
rect 4660 28864 4976 28865
rect 4660 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4976 28864
rect 4660 28799 4976 28800
rect 12088 28864 12404 28865
rect 12088 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12404 28864
rect 12088 28799 12404 28800
rect 19516 28864 19832 28865
rect 19516 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19832 28864
rect 19516 28799 19832 28800
rect 26944 28864 27260 28865
rect 26944 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27260 28864
rect 26944 28799 27260 28800
rect 5320 28320 5636 28321
rect 5320 28256 5326 28320
rect 5390 28256 5406 28320
rect 5470 28256 5486 28320
rect 5550 28256 5566 28320
rect 5630 28256 5636 28320
rect 5320 28255 5636 28256
rect 12748 28320 13064 28321
rect 12748 28256 12754 28320
rect 12818 28256 12834 28320
rect 12898 28256 12914 28320
rect 12978 28256 12994 28320
rect 13058 28256 13064 28320
rect 12748 28255 13064 28256
rect 20176 28320 20492 28321
rect 20176 28256 20182 28320
rect 20246 28256 20262 28320
rect 20326 28256 20342 28320
rect 20406 28256 20422 28320
rect 20486 28256 20492 28320
rect 20176 28255 20492 28256
rect 27604 28320 27920 28321
rect 27604 28256 27610 28320
rect 27674 28256 27690 28320
rect 27754 28256 27770 28320
rect 27834 28256 27850 28320
rect 27914 28256 27920 28320
rect 27604 28255 27920 28256
rect 4660 27776 4976 27777
rect 4660 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4976 27776
rect 4660 27711 4976 27712
rect 12088 27776 12404 27777
rect 12088 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12404 27776
rect 12088 27711 12404 27712
rect 19516 27776 19832 27777
rect 19516 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19832 27776
rect 19516 27711 19832 27712
rect 26944 27776 27260 27777
rect 26944 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27260 27776
rect 26944 27711 27260 27712
rect 5320 27232 5636 27233
rect 5320 27168 5326 27232
rect 5390 27168 5406 27232
rect 5470 27168 5486 27232
rect 5550 27168 5566 27232
rect 5630 27168 5636 27232
rect 5320 27167 5636 27168
rect 12748 27232 13064 27233
rect 12748 27168 12754 27232
rect 12818 27168 12834 27232
rect 12898 27168 12914 27232
rect 12978 27168 12994 27232
rect 13058 27168 13064 27232
rect 12748 27167 13064 27168
rect 20176 27232 20492 27233
rect 20176 27168 20182 27232
rect 20246 27168 20262 27232
rect 20326 27168 20342 27232
rect 20406 27168 20422 27232
rect 20486 27168 20492 27232
rect 20176 27167 20492 27168
rect 27604 27232 27920 27233
rect 27604 27168 27610 27232
rect 27674 27168 27690 27232
rect 27754 27168 27770 27232
rect 27834 27168 27850 27232
rect 27914 27168 27920 27232
rect 27604 27167 27920 27168
rect 4660 26688 4976 26689
rect 4660 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4976 26688
rect 4660 26623 4976 26624
rect 12088 26688 12404 26689
rect 12088 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12404 26688
rect 12088 26623 12404 26624
rect 19516 26688 19832 26689
rect 19516 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19832 26688
rect 19516 26623 19832 26624
rect 26944 26688 27260 26689
rect 26944 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27260 26688
rect 26944 26623 27260 26624
rect 5320 26144 5636 26145
rect 5320 26080 5326 26144
rect 5390 26080 5406 26144
rect 5470 26080 5486 26144
rect 5550 26080 5566 26144
rect 5630 26080 5636 26144
rect 5320 26079 5636 26080
rect 12748 26144 13064 26145
rect 12748 26080 12754 26144
rect 12818 26080 12834 26144
rect 12898 26080 12914 26144
rect 12978 26080 12994 26144
rect 13058 26080 13064 26144
rect 12748 26079 13064 26080
rect 20176 26144 20492 26145
rect 20176 26080 20182 26144
rect 20246 26080 20262 26144
rect 20326 26080 20342 26144
rect 20406 26080 20422 26144
rect 20486 26080 20492 26144
rect 20176 26079 20492 26080
rect 27604 26144 27920 26145
rect 27604 26080 27610 26144
rect 27674 26080 27690 26144
rect 27754 26080 27770 26144
rect 27834 26080 27850 26144
rect 27914 26080 27920 26144
rect 27604 26079 27920 26080
rect 0 25938 800 25968
rect 3969 25938 4035 25941
rect 0 25936 4035 25938
rect 0 25880 3974 25936
rect 4030 25880 4035 25936
rect 0 25878 4035 25880
rect 0 25848 800 25878
rect 3969 25875 4035 25878
rect 4660 25600 4976 25601
rect 4660 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4976 25600
rect 4660 25535 4976 25536
rect 12088 25600 12404 25601
rect 12088 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12404 25600
rect 12088 25535 12404 25536
rect 19516 25600 19832 25601
rect 19516 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19832 25600
rect 19516 25535 19832 25536
rect 26944 25600 27260 25601
rect 26944 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27260 25600
rect 26944 25535 27260 25536
rect 5320 25056 5636 25057
rect 5320 24992 5326 25056
rect 5390 24992 5406 25056
rect 5470 24992 5486 25056
rect 5550 24992 5566 25056
rect 5630 24992 5636 25056
rect 5320 24991 5636 24992
rect 12748 25056 13064 25057
rect 12748 24992 12754 25056
rect 12818 24992 12834 25056
rect 12898 24992 12914 25056
rect 12978 24992 12994 25056
rect 13058 24992 13064 25056
rect 12748 24991 13064 24992
rect 20176 25056 20492 25057
rect 20176 24992 20182 25056
rect 20246 24992 20262 25056
rect 20326 24992 20342 25056
rect 20406 24992 20422 25056
rect 20486 24992 20492 25056
rect 20176 24991 20492 24992
rect 27604 25056 27920 25057
rect 27604 24992 27610 25056
rect 27674 24992 27690 25056
rect 27754 24992 27770 25056
rect 27834 24992 27850 25056
rect 27914 24992 27920 25056
rect 27604 24991 27920 24992
rect 4660 24512 4976 24513
rect 4660 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4976 24512
rect 4660 24447 4976 24448
rect 12088 24512 12404 24513
rect 12088 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12404 24512
rect 12088 24447 12404 24448
rect 19516 24512 19832 24513
rect 19516 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19832 24512
rect 19516 24447 19832 24448
rect 26944 24512 27260 24513
rect 26944 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27260 24512
rect 26944 24447 27260 24448
rect 5320 23968 5636 23969
rect 5320 23904 5326 23968
rect 5390 23904 5406 23968
rect 5470 23904 5486 23968
rect 5550 23904 5566 23968
rect 5630 23904 5636 23968
rect 5320 23903 5636 23904
rect 12748 23968 13064 23969
rect 12748 23904 12754 23968
rect 12818 23904 12834 23968
rect 12898 23904 12914 23968
rect 12978 23904 12994 23968
rect 13058 23904 13064 23968
rect 12748 23903 13064 23904
rect 20176 23968 20492 23969
rect 20176 23904 20182 23968
rect 20246 23904 20262 23968
rect 20326 23904 20342 23968
rect 20406 23904 20422 23968
rect 20486 23904 20492 23968
rect 20176 23903 20492 23904
rect 27604 23968 27920 23969
rect 27604 23904 27610 23968
rect 27674 23904 27690 23968
rect 27754 23904 27770 23968
rect 27834 23904 27850 23968
rect 27914 23904 27920 23968
rect 27604 23903 27920 23904
rect 4660 23424 4976 23425
rect 4660 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4976 23424
rect 4660 23359 4976 23360
rect 12088 23424 12404 23425
rect 12088 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12404 23424
rect 12088 23359 12404 23360
rect 19516 23424 19832 23425
rect 19516 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19832 23424
rect 19516 23359 19832 23360
rect 26944 23424 27260 23425
rect 26944 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27260 23424
rect 26944 23359 27260 23360
rect 5320 22880 5636 22881
rect 5320 22816 5326 22880
rect 5390 22816 5406 22880
rect 5470 22816 5486 22880
rect 5550 22816 5566 22880
rect 5630 22816 5636 22880
rect 5320 22815 5636 22816
rect 12748 22880 13064 22881
rect 12748 22816 12754 22880
rect 12818 22816 12834 22880
rect 12898 22816 12914 22880
rect 12978 22816 12994 22880
rect 13058 22816 13064 22880
rect 12748 22815 13064 22816
rect 20176 22880 20492 22881
rect 20176 22816 20182 22880
rect 20246 22816 20262 22880
rect 20326 22816 20342 22880
rect 20406 22816 20422 22880
rect 20486 22816 20492 22880
rect 20176 22815 20492 22816
rect 27604 22880 27920 22881
rect 27604 22816 27610 22880
rect 27674 22816 27690 22880
rect 27754 22816 27770 22880
rect 27834 22816 27850 22880
rect 27914 22816 27920 22880
rect 27604 22815 27920 22816
rect 4660 22336 4976 22337
rect 4660 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4976 22336
rect 4660 22271 4976 22272
rect 12088 22336 12404 22337
rect 12088 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12404 22336
rect 12088 22271 12404 22272
rect 19516 22336 19832 22337
rect 19516 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19832 22336
rect 19516 22271 19832 22272
rect 26944 22336 27260 22337
rect 26944 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27260 22336
rect 26944 22271 27260 22272
rect 21817 21994 21883 21997
rect 26325 21994 26391 21997
rect 21817 21992 26391 21994
rect 21817 21936 21822 21992
rect 21878 21936 26330 21992
rect 26386 21936 26391 21992
rect 21817 21934 26391 21936
rect 21817 21931 21883 21934
rect 26325 21931 26391 21934
rect 28073 21858 28139 21861
rect 31200 21858 32000 21888
rect 28073 21856 32000 21858
rect 28073 21800 28078 21856
rect 28134 21800 32000 21856
rect 28073 21798 32000 21800
rect 28073 21795 28139 21798
rect 5320 21792 5636 21793
rect 5320 21728 5326 21792
rect 5390 21728 5406 21792
rect 5470 21728 5486 21792
rect 5550 21728 5566 21792
rect 5630 21728 5636 21792
rect 5320 21727 5636 21728
rect 12748 21792 13064 21793
rect 12748 21728 12754 21792
rect 12818 21728 12834 21792
rect 12898 21728 12914 21792
rect 12978 21728 12994 21792
rect 13058 21728 13064 21792
rect 12748 21727 13064 21728
rect 20176 21792 20492 21793
rect 20176 21728 20182 21792
rect 20246 21728 20262 21792
rect 20326 21728 20342 21792
rect 20406 21728 20422 21792
rect 20486 21728 20492 21792
rect 20176 21727 20492 21728
rect 27604 21792 27920 21793
rect 27604 21728 27610 21792
rect 27674 21728 27690 21792
rect 27754 21728 27770 21792
rect 27834 21728 27850 21792
rect 27914 21728 27920 21792
rect 31200 21768 32000 21798
rect 27604 21727 27920 21728
rect 14549 21314 14615 21317
rect 18321 21314 18387 21317
rect 14549 21312 18387 21314
rect 14549 21256 14554 21312
rect 14610 21256 18326 21312
rect 18382 21256 18387 21312
rect 14549 21254 18387 21256
rect 14549 21251 14615 21254
rect 18321 21251 18387 21254
rect 4660 21248 4976 21249
rect 0 21178 800 21208
rect 4660 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4976 21248
rect 4660 21183 4976 21184
rect 12088 21248 12404 21249
rect 12088 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12404 21248
rect 12088 21183 12404 21184
rect 19516 21248 19832 21249
rect 19516 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19832 21248
rect 19516 21183 19832 21184
rect 26944 21248 27260 21249
rect 26944 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27260 21248
rect 26944 21183 27260 21184
rect 933 21178 999 21181
rect 31200 21178 32000 21208
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 28950 21118 32000 21178
rect 25865 21042 25931 21045
rect 27153 21042 27219 21045
rect 28950 21042 29010 21118
rect 31200 21088 32000 21118
rect 25865 21040 29010 21042
rect 25865 20984 25870 21040
rect 25926 20984 27158 21040
rect 27214 20984 29010 21040
rect 25865 20982 29010 20984
rect 25865 20979 25931 20982
rect 27153 20979 27219 20982
rect 5320 20704 5636 20705
rect 5320 20640 5326 20704
rect 5390 20640 5406 20704
rect 5470 20640 5486 20704
rect 5550 20640 5566 20704
rect 5630 20640 5636 20704
rect 5320 20639 5636 20640
rect 12748 20704 13064 20705
rect 12748 20640 12754 20704
rect 12818 20640 12834 20704
rect 12898 20640 12914 20704
rect 12978 20640 12994 20704
rect 13058 20640 13064 20704
rect 12748 20639 13064 20640
rect 20176 20704 20492 20705
rect 20176 20640 20182 20704
rect 20246 20640 20262 20704
rect 20326 20640 20342 20704
rect 20406 20640 20422 20704
rect 20486 20640 20492 20704
rect 20176 20639 20492 20640
rect 27604 20704 27920 20705
rect 27604 20640 27610 20704
rect 27674 20640 27690 20704
rect 27754 20640 27770 20704
rect 27834 20640 27850 20704
rect 27914 20640 27920 20704
rect 27604 20639 27920 20640
rect 1485 20634 1551 20637
rect 798 20632 1551 20634
rect 798 20576 1490 20632
rect 1546 20576 1551 20632
rect 798 20574 1551 20576
rect 798 20528 858 20574
rect 1485 20571 1551 20574
rect 0 20438 858 20528
rect 27613 20498 27679 20501
rect 31200 20498 32000 20528
rect 27613 20496 32000 20498
rect 27613 20440 27618 20496
rect 27674 20440 32000 20496
rect 27613 20438 32000 20440
rect 0 20408 800 20438
rect 27613 20435 27679 20438
rect 31200 20408 32000 20438
rect 28993 20362 29059 20365
rect 29545 20362 29611 20365
rect 28993 20360 29611 20362
rect 28993 20304 28998 20360
rect 29054 20304 29550 20360
rect 29606 20304 29611 20360
rect 28993 20302 29611 20304
rect 28993 20299 29059 20302
rect 29545 20299 29611 20302
rect 4660 20160 4976 20161
rect 4660 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4976 20160
rect 4660 20095 4976 20096
rect 12088 20160 12404 20161
rect 12088 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12404 20160
rect 12088 20095 12404 20096
rect 19516 20160 19832 20161
rect 19516 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19832 20160
rect 19516 20095 19832 20096
rect 26944 20160 27260 20161
rect 26944 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27260 20160
rect 26944 20095 27260 20096
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 28625 19818 28691 19821
rect 31200 19818 32000 19848
rect 28625 19816 32000 19818
rect 28625 19760 28630 19816
rect 28686 19760 32000 19816
rect 28625 19758 32000 19760
rect 28625 19755 28691 19758
rect 31200 19728 32000 19758
rect 5320 19616 5636 19617
rect 5320 19552 5326 19616
rect 5390 19552 5406 19616
rect 5470 19552 5486 19616
rect 5550 19552 5566 19616
rect 5630 19552 5636 19616
rect 5320 19551 5636 19552
rect 12748 19616 13064 19617
rect 12748 19552 12754 19616
rect 12818 19552 12834 19616
rect 12898 19552 12914 19616
rect 12978 19552 12994 19616
rect 13058 19552 13064 19616
rect 12748 19551 13064 19552
rect 20176 19616 20492 19617
rect 20176 19552 20182 19616
rect 20246 19552 20262 19616
rect 20326 19552 20342 19616
rect 20406 19552 20422 19616
rect 20486 19552 20492 19616
rect 20176 19551 20492 19552
rect 27604 19616 27920 19617
rect 27604 19552 27610 19616
rect 27674 19552 27690 19616
rect 27754 19552 27770 19616
rect 27834 19552 27850 19616
rect 27914 19552 27920 19616
rect 27604 19551 27920 19552
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 4660 19072 4976 19073
rect 4660 19008 4666 19072
rect 4730 19008 4746 19072
rect 4810 19008 4826 19072
rect 4890 19008 4906 19072
rect 4970 19008 4976 19072
rect 4660 19007 4976 19008
rect 12088 19072 12404 19073
rect 12088 19008 12094 19072
rect 12158 19008 12174 19072
rect 12238 19008 12254 19072
rect 12318 19008 12334 19072
rect 12398 19008 12404 19072
rect 12088 19007 12404 19008
rect 19516 19072 19832 19073
rect 19516 19008 19522 19072
rect 19586 19008 19602 19072
rect 19666 19008 19682 19072
rect 19746 19008 19762 19072
rect 19826 19008 19832 19072
rect 19516 19007 19832 19008
rect 26944 19072 27260 19073
rect 26944 19008 26950 19072
rect 27014 19008 27030 19072
rect 27094 19008 27110 19072
rect 27174 19008 27190 19072
rect 27254 19008 27260 19072
rect 26944 19007 27260 19008
rect 5320 18528 5636 18529
rect 0 18458 800 18488
rect 5320 18464 5326 18528
rect 5390 18464 5406 18528
rect 5470 18464 5486 18528
rect 5550 18464 5566 18528
rect 5630 18464 5636 18528
rect 5320 18463 5636 18464
rect 12748 18528 13064 18529
rect 12748 18464 12754 18528
rect 12818 18464 12834 18528
rect 12898 18464 12914 18528
rect 12978 18464 12994 18528
rect 13058 18464 13064 18528
rect 12748 18463 13064 18464
rect 20176 18528 20492 18529
rect 20176 18464 20182 18528
rect 20246 18464 20262 18528
rect 20326 18464 20342 18528
rect 20406 18464 20422 18528
rect 20486 18464 20492 18528
rect 20176 18463 20492 18464
rect 27604 18528 27920 18529
rect 27604 18464 27610 18528
rect 27674 18464 27690 18528
rect 27754 18464 27770 18528
rect 27834 18464 27850 18528
rect 27914 18464 27920 18528
rect 27604 18463 27920 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 28625 18458 28691 18461
rect 31200 18458 32000 18488
rect 28625 18456 32000 18458
rect 28625 18400 28630 18456
rect 28686 18400 32000 18456
rect 28625 18398 32000 18400
rect 28625 18395 28691 18398
rect 31200 18368 32000 18398
rect 4660 17984 4976 17985
rect 4660 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4976 17984
rect 4660 17919 4976 17920
rect 12088 17984 12404 17985
rect 12088 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12404 17984
rect 12088 17919 12404 17920
rect 19516 17984 19832 17985
rect 19516 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19832 17984
rect 19516 17919 19832 17920
rect 26944 17984 27260 17985
rect 26944 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27260 17984
rect 26944 17919 27260 17920
rect 27613 17778 27679 17781
rect 31200 17778 32000 17808
rect 27613 17776 32000 17778
rect 27613 17720 27618 17776
rect 27674 17720 32000 17776
rect 27613 17718 32000 17720
rect 27613 17715 27679 17718
rect 31200 17688 32000 17718
rect 5320 17440 5636 17441
rect 5320 17376 5326 17440
rect 5390 17376 5406 17440
rect 5470 17376 5486 17440
rect 5550 17376 5566 17440
rect 5630 17376 5636 17440
rect 5320 17375 5636 17376
rect 12748 17440 13064 17441
rect 12748 17376 12754 17440
rect 12818 17376 12834 17440
rect 12898 17376 12914 17440
rect 12978 17376 12994 17440
rect 13058 17376 13064 17440
rect 12748 17375 13064 17376
rect 20176 17440 20492 17441
rect 20176 17376 20182 17440
rect 20246 17376 20262 17440
rect 20326 17376 20342 17440
rect 20406 17376 20422 17440
rect 20486 17376 20492 17440
rect 20176 17375 20492 17376
rect 27604 17440 27920 17441
rect 27604 17376 27610 17440
rect 27674 17376 27690 17440
rect 27754 17376 27770 17440
rect 27834 17376 27850 17440
rect 27914 17376 27920 17440
rect 27604 17375 27920 17376
rect 0 17098 800 17128
rect 7925 17098 7991 17101
rect 0 17096 7991 17098
rect 0 17040 7930 17096
rect 7986 17040 7991 17096
rect 0 17038 7991 17040
rect 0 17008 800 17038
rect 7925 17035 7991 17038
rect 27797 17098 27863 17101
rect 31200 17098 32000 17128
rect 27797 17096 32000 17098
rect 27797 17040 27802 17096
rect 27858 17040 32000 17096
rect 27797 17038 32000 17040
rect 27797 17035 27863 17038
rect 31200 17008 32000 17038
rect 4660 16896 4976 16897
rect 4660 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4976 16896
rect 4660 16831 4976 16832
rect 12088 16896 12404 16897
rect 12088 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12404 16896
rect 12088 16831 12404 16832
rect 19516 16896 19832 16897
rect 19516 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19832 16896
rect 19516 16831 19832 16832
rect 26944 16896 27260 16897
rect 26944 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27260 16896
rect 26944 16831 27260 16832
rect 0 16418 800 16448
rect 4429 16418 4495 16421
rect 0 16416 4495 16418
rect 0 16360 4434 16416
rect 4490 16360 4495 16416
rect 0 16358 4495 16360
rect 0 16328 800 16358
rect 4429 16355 4495 16358
rect 30373 16418 30439 16421
rect 31200 16418 32000 16448
rect 30373 16416 32000 16418
rect 30373 16360 30378 16416
rect 30434 16360 32000 16416
rect 30373 16358 32000 16360
rect 30373 16355 30439 16358
rect 5320 16352 5636 16353
rect 5320 16288 5326 16352
rect 5390 16288 5406 16352
rect 5470 16288 5486 16352
rect 5550 16288 5566 16352
rect 5630 16288 5636 16352
rect 5320 16287 5636 16288
rect 12748 16352 13064 16353
rect 12748 16288 12754 16352
rect 12818 16288 12834 16352
rect 12898 16288 12914 16352
rect 12978 16288 12994 16352
rect 13058 16288 13064 16352
rect 12748 16287 13064 16288
rect 20176 16352 20492 16353
rect 20176 16288 20182 16352
rect 20246 16288 20262 16352
rect 20326 16288 20342 16352
rect 20406 16288 20422 16352
rect 20486 16288 20492 16352
rect 20176 16287 20492 16288
rect 27604 16352 27920 16353
rect 27604 16288 27610 16352
rect 27674 16288 27690 16352
rect 27754 16288 27770 16352
rect 27834 16288 27850 16352
rect 27914 16288 27920 16352
rect 31200 16328 32000 16358
rect 27604 16287 27920 16288
rect 4660 15808 4976 15809
rect 0 15738 800 15768
rect 4660 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4976 15808
rect 4660 15743 4976 15744
rect 12088 15808 12404 15809
rect 12088 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12404 15808
rect 12088 15743 12404 15744
rect 19516 15808 19832 15809
rect 19516 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19832 15808
rect 19516 15743 19832 15744
rect 26944 15808 27260 15809
rect 26944 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27260 15808
rect 26944 15743 27260 15744
rect 4337 15738 4403 15741
rect 0 15736 4403 15738
rect 0 15680 4342 15736
rect 4398 15680 4403 15736
rect 0 15678 4403 15680
rect 0 15648 800 15678
rect 4337 15675 4403 15678
rect 27613 15738 27679 15741
rect 31200 15738 32000 15768
rect 27613 15736 32000 15738
rect 27613 15680 27618 15736
rect 27674 15680 32000 15736
rect 27613 15678 32000 15680
rect 27613 15675 27679 15678
rect 31200 15648 32000 15678
rect 12525 15466 12591 15469
rect 13721 15466 13787 15469
rect 15929 15466 15995 15469
rect 12525 15464 15995 15466
rect 12525 15408 12530 15464
rect 12586 15408 13726 15464
rect 13782 15408 15934 15464
rect 15990 15408 15995 15464
rect 12525 15406 15995 15408
rect 12525 15403 12591 15406
rect 13721 15403 13787 15406
rect 15929 15403 15995 15406
rect 5320 15264 5636 15265
rect 5320 15200 5326 15264
rect 5390 15200 5406 15264
rect 5470 15200 5486 15264
rect 5550 15200 5566 15264
rect 5630 15200 5636 15264
rect 5320 15199 5636 15200
rect 12748 15264 13064 15265
rect 12748 15200 12754 15264
rect 12818 15200 12834 15264
rect 12898 15200 12914 15264
rect 12978 15200 12994 15264
rect 13058 15200 13064 15264
rect 12748 15199 13064 15200
rect 20176 15264 20492 15265
rect 20176 15200 20182 15264
rect 20246 15200 20262 15264
rect 20326 15200 20342 15264
rect 20406 15200 20422 15264
rect 20486 15200 20492 15264
rect 20176 15199 20492 15200
rect 27604 15264 27920 15265
rect 27604 15200 27610 15264
rect 27674 15200 27690 15264
rect 27754 15200 27770 15264
rect 27834 15200 27850 15264
rect 27914 15200 27920 15264
rect 27604 15199 27920 15200
rect 0 15058 800 15088
rect 4061 15058 4127 15061
rect 0 15056 4127 15058
rect 0 15000 4066 15056
rect 4122 15000 4127 15056
rect 0 14998 4127 15000
rect 0 14968 800 14998
rect 4061 14995 4127 14998
rect 4660 14720 4976 14721
rect 4660 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4976 14720
rect 4660 14655 4976 14656
rect 12088 14720 12404 14721
rect 12088 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12404 14720
rect 12088 14655 12404 14656
rect 19516 14720 19832 14721
rect 19516 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19832 14720
rect 19516 14655 19832 14656
rect 26944 14720 27260 14721
rect 26944 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27260 14720
rect 26944 14655 27260 14656
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 5320 14176 5636 14177
rect 5320 14112 5326 14176
rect 5390 14112 5406 14176
rect 5470 14112 5486 14176
rect 5550 14112 5566 14176
rect 5630 14112 5636 14176
rect 5320 14111 5636 14112
rect 12748 14176 13064 14177
rect 12748 14112 12754 14176
rect 12818 14112 12834 14176
rect 12898 14112 12914 14176
rect 12978 14112 12994 14176
rect 13058 14112 13064 14176
rect 12748 14111 13064 14112
rect 20176 14176 20492 14177
rect 20176 14112 20182 14176
rect 20246 14112 20262 14176
rect 20326 14112 20342 14176
rect 20406 14112 20422 14176
rect 20486 14112 20492 14176
rect 20176 14111 20492 14112
rect 27604 14176 27920 14177
rect 27604 14112 27610 14176
rect 27674 14112 27690 14176
rect 27754 14112 27770 14176
rect 27834 14112 27850 14176
rect 27914 14112 27920 14176
rect 27604 14111 27920 14112
rect 8661 13834 8727 13837
rect 10777 13834 10843 13837
rect 8661 13832 10843 13834
rect 8661 13776 8666 13832
rect 8722 13776 10782 13832
rect 10838 13776 10843 13832
rect 8661 13774 10843 13776
rect 8661 13771 8727 13774
rect 10777 13771 10843 13774
rect 0 13698 800 13728
rect 4061 13698 4127 13701
rect 0 13696 4127 13698
rect 0 13640 4066 13696
rect 4122 13640 4127 13696
rect 0 13638 4127 13640
rect 0 13608 800 13638
rect 4061 13635 4127 13638
rect 27337 13698 27403 13701
rect 31200 13698 32000 13728
rect 27337 13696 32000 13698
rect 27337 13640 27342 13696
rect 27398 13640 32000 13696
rect 27337 13638 32000 13640
rect 27337 13635 27403 13638
rect 4660 13632 4976 13633
rect 4660 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4976 13632
rect 4660 13567 4976 13568
rect 12088 13632 12404 13633
rect 12088 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12404 13632
rect 12088 13567 12404 13568
rect 19516 13632 19832 13633
rect 19516 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19832 13632
rect 19516 13567 19832 13568
rect 26944 13632 27260 13633
rect 26944 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27260 13632
rect 31200 13608 32000 13638
rect 26944 13567 27260 13568
rect 5320 13088 5636 13089
rect 5320 13024 5326 13088
rect 5390 13024 5406 13088
rect 5470 13024 5486 13088
rect 5550 13024 5566 13088
rect 5630 13024 5636 13088
rect 5320 13023 5636 13024
rect 12748 13088 13064 13089
rect 12748 13024 12754 13088
rect 12818 13024 12834 13088
rect 12898 13024 12914 13088
rect 12978 13024 12994 13088
rect 13058 13024 13064 13088
rect 12748 13023 13064 13024
rect 20176 13088 20492 13089
rect 20176 13024 20182 13088
rect 20246 13024 20262 13088
rect 20326 13024 20342 13088
rect 20406 13024 20422 13088
rect 20486 13024 20492 13088
rect 20176 13023 20492 13024
rect 27604 13088 27920 13089
rect 27604 13024 27610 13088
rect 27674 13024 27690 13088
rect 27754 13024 27770 13088
rect 27834 13024 27850 13088
rect 27914 13024 27920 13088
rect 27604 13023 27920 13024
rect 4660 12544 4976 12545
rect 4660 12480 4666 12544
rect 4730 12480 4746 12544
rect 4810 12480 4826 12544
rect 4890 12480 4906 12544
rect 4970 12480 4976 12544
rect 4660 12479 4976 12480
rect 12088 12544 12404 12545
rect 12088 12480 12094 12544
rect 12158 12480 12174 12544
rect 12238 12480 12254 12544
rect 12318 12480 12334 12544
rect 12398 12480 12404 12544
rect 12088 12479 12404 12480
rect 19516 12544 19832 12545
rect 19516 12480 19522 12544
rect 19586 12480 19602 12544
rect 19666 12480 19682 12544
rect 19746 12480 19762 12544
rect 19826 12480 19832 12544
rect 19516 12479 19832 12480
rect 26944 12544 27260 12545
rect 26944 12480 26950 12544
rect 27014 12480 27030 12544
rect 27094 12480 27110 12544
rect 27174 12480 27190 12544
rect 27254 12480 27260 12544
rect 26944 12479 27260 12480
rect 11053 12474 11119 12477
rect 11605 12474 11671 12477
rect 11053 12472 11671 12474
rect 11053 12416 11058 12472
rect 11114 12416 11610 12472
rect 11666 12416 11671 12472
rect 11053 12414 11671 12416
rect 11053 12411 11119 12414
rect 11605 12411 11671 12414
rect 0 12338 800 12368
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12248 800 12278
rect 3969 12275 4035 12278
rect 5320 12000 5636 12001
rect 5320 11936 5326 12000
rect 5390 11936 5406 12000
rect 5470 11936 5486 12000
rect 5550 11936 5566 12000
rect 5630 11936 5636 12000
rect 5320 11935 5636 11936
rect 12748 12000 13064 12001
rect 12748 11936 12754 12000
rect 12818 11936 12834 12000
rect 12898 11936 12914 12000
rect 12978 11936 12994 12000
rect 13058 11936 13064 12000
rect 12748 11935 13064 11936
rect 20176 12000 20492 12001
rect 20176 11936 20182 12000
rect 20246 11936 20262 12000
rect 20326 11936 20342 12000
rect 20406 11936 20422 12000
rect 20486 11936 20492 12000
rect 20176 11935 20492 11936
rect 27604 12000 27920 12001
rect 27604 11936 27610 12000
rect 27674 11936 27690 12000
rect 27754 11936 27770 12000
rect 27834 11936 27850 12000
rect 27914 11936 27920 12000
rect 27604 11935 27920 11936
rect 4660 11456 4976 11457
rect 4660 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4976 11456
rect 4660 11391 4976 11392
rect 12088 11456 12404 11457
rect 12088 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12404 11456
rect 12088 11391 12404 11392
rect 19516 11456 19832 11457
rect 19516 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19832 11456
rect 19516 11391 19832 11392
rect 26944 11456 27260 11457
rect 26944 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27260 11456
rect 26944 11391 27260 11392
rect 21817 11114 21883 11117
rect 21817 11112 29010 11114
rect 21817 11056 21822 11112
rect 21878 11056 29010 11112
rect 21817 11054 29010 11056
rect 21817 11051 21883 11054
rect 0 10978 800 11008
rect 3969 10978 4035 10981
rect 0 10976 4035 10978
rect 0 10920 3974 10976
rect 4030 10920 4035 10976
rect 0 10918 4035 10920
rect 28950 10978 29010 11054
rect 31200 10978 32000 11008
rect 28950 10918 32000 10978
rect 0 10888 800 10918
rect 3969 10915 4035 10918
rect 5320 10912 5636 10913
rect 5320 10848 5326 10912
rect 5390 10848 5406 10912
rect 5470 10848 5486 10912
rect 5550 10848 5566 10912
rect 5630 10848 5636 10912
rect 5320 10847 5636 10848
rect 12748 10912 13064 10913
rect 12748 10848 12754 10912
rect 12818 10848 12834 10912
rect 12898 10848 12914 10912
rect 12978 10848 12994 10912
rect 13058 10848 13064 10912
rect 12748 10847 13064 10848
rect 20176 10912 20492 10913
rect 20176 10848 20182 10912
rect 20246 10848 20262 10912
rect 20326 10848 20342 10912
rect 20406 10848 20422 10912
rect 20486 10848 20492 10912
rect 20176 10847 20492 10848
rect 27604 10912 27920 10913
rect 27604 10848 27610 10912
rect 27674 10848 27690 10912
rect 27754 10848 27770 10912
rect 27834 10848 27850 10912
rect 27914 10848 27920 10912
rect 31200 10888 32000 10918
rect 27604 10847 27920 10848
rect 4660 10368 4976 10369
rect 4660 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4976 10368
rect 4660 10303 4976 10304
rect 12088 10368 12404 10369
rect 12088 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12404 10368
rect 12088 10303 12404 10304
rect 19516 10368 19832 10369
rect 19516 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19832 10368
rect 19516 10303 19832 10304
rect 26944 10368 27260 10369
rect 26944 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27260 10368
rect 26944 10303 27260 10304
rect 5320 9824 5636 9825
rect 5320 9760 5326 9824
rect 5390 9760 5406 9824
rect 5470 9760 5486 9824
rect 5550 9760 5566 9824
rect 5630 9760 5636 9824
rect 5320 9759 5636 9760
rect 12748 9824 13064 9825
rect 12748 9760 12754 9824
rect 12818 9760 12834 9824
rect 12898 9760 12914 9824
rect 12978 9760 12994 9824
rect 13058 9760 13064 9824
rect 12748 9759 13064 9760
rect 20176 9824 20492 9825
rect 20176 9760 20182 9824
rect 20246 9760 20262 9824
rect 20326 9760 20342 9824
rect 20406 9760 20422 9824
rect 20486 9760 20492 9824
rect 20176 9759 20492 9760
rect 27604 9824 27920 9825
rect 27604 9760 27610 9824
rect 27674 9760 27690 9824
rect 27754 9760 27770 9824
rect 27834 9760 27850 9824
rect 27914 9760 27920 9824
rect 27604 9759 27920 9760
rect 0 9618 800 9648
rect 4061 9618 4127 9621
rect 0 9616 4127 9618
rect 0 9560 4066 9616
rect 4122 9560 4127 9616
rect 0 9558 4127 9560
rect 0 9528 800 9558
rect 4061 9555 4127 9558
rect 4660 9280 4976 9281
rect 4660 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4976 9280
rect 4660 9215 4976 9216
rect 12088 9280 12404 9281
rect 12088 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12404 9280
rect 12088 9215 12404 9216
rect 19516 9280 19832 9281
rect 19516 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19832 9280
rect 19516 9215 19832 9216
rect 26944 9280 27260 9281
rect 26944 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27260 9280
rect 26944 9215 27260 9216
rect 5320 8736 5636 8737
rect 5320 8672 5326 8736
rect 5390 8672 5406 8736
rect 5470 8672 5486 8736
rect 5550 8672 5566 8736
rect 5630 8672 5636 8736
rect 5320 8671 5636 8672
rect 12748 8736 13064 8737
rect 12748 8672 12754 8736
rect 12818 8672 12834 8736
rect 12898 8672 12914 8736
rect 12978 8672 12994 8736
rect 13058 8672 13064 8736
rect 12748 8671 13064 8672
rect 20176 8736 20492 8737
rect 20176 8672 20182 8736
rect 20246 8672 20262 8736
rect 20326 8672 20342 8736
rect 20406 8672 20422 8736
rect 20486 8672 20492 8736
rect 20176 8671 20492 8672
rect 27604 8736 27920 8737
rect 27604 8672 27610 8736
rect 27674 8672 27690 8736
rect 27754 8672 27770 8736
rect 27834 8672 27850 8736
rect 27914 8672 27920 8736
rect 27604 8671 27920 8672
rect 0 8258 800 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 800 8198
rect 4061 8195 4127 8198
rect 4660 8192 4976 8193
rect 4660 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4976 8192
rect 4660 8127 4976 8128
rect 12088 8192 12404 8193
rect 12088 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12404 8192
rect 12088 8127 12404 8128
rect 19516 8192 19832 8193
rect 19516 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19832 8192
rect 19516 8127 19832 8128
rect 26944 8192 27260 8193
rect 26944 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27260 8192
rect 26944 8127 27260 8128
rect 8845 7986 8911 7989
rect 9581 7986 9647 7989
rect 8845 7984 9647 7986
rect 8845 7928 8850 7984
rect 8906 7928 9586 7984
rect 9642 7928 9647 7984
rect 8845 7926 9647 7928
rect 8845 7923 8911 7926
rect 9581 7923 9647 7926
rect 5320 7648 5636 7649
rect 5320 7584 5326 7648
rect 5390 7584 5406 7648
rect 5470 7584 5486 7648
rect 5550 7584 5566 7648
rect 5630 7584 5636 7648
rect 5320 7583 5636 7584
rect 12748 7648 13064 7649
rect 12748 7584 12754 7648
rect 12818 7584 12834 7648
rect 12898 7584 12914 7648
rect 12978 7584 12994 7648
rect 13058 7584 13064 7648
rect 12748 7583 13064 7584
rect 20176 7648 20492 7649
rect 20176 7584 20182 7648
rect 20246 7584 20262 7648
rect 20326 7584 20342 7648
rect 20406 7584 20422 7648
rect 20486 7584 20492 7648
rect 20176 7583 20492 7584
rect 27604 7648 27920 7649
rect 27604 7584 27610 7648
rect 27674 7584 27690 7648
rect 27754 7584 27770 7648
rect 27834 7584 27850 7648
rect 27914 7584 27920 7648
rect 27604 7583 27920 7584
rect 4660 7104 4976 7105
rect 4660 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4976 7104
rect 4660 7039 4976 7040
rect 12088 7104 12404 7105
rect 12088 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12404 7104
rect 12088 7039 12404 7040
rect 19516 7104 19832 7105
rect 19516 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19832 7104
rect 19516 7039 19832 7040
rect 26944 7104 27260 7105
rect 26944 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27260 7104
rect 26944 7039 27260 7040
rect 5320 6560 5636 6561
rect 5320 6496 5326 6560
rect 5390 6496 5406 6560
rect 5470 6496 5486 6560
rect 5550 6496 5566 6560
rect 5630 6496 5636 6560
rect 5320 6495 5636 6496
rect 12748 6560 13064 6561
rect 12748 6496 12754 6560
rect 12818 6496 12834 6560
rect 12898 6496 12914 6560
rect 12978 6496 12994 6560
rect 13058 6496 13064 6560
rect 12748 6495 13064 6496
rect 20176 6560 20492 6561
rect 20176 6496 20182 6560
rect 20246 6496 20262 6560
rect 20326 6496 20342 6560
rect 20406 6496 20422 6560
rect 20486 6496 20492 6560
rect 20176 6495 20492 6496
rect 27604 6560 27920 6561
rect 27604 6496 27610 6560
rect 27674 6496 27690 6560
rect 27754 6496 27770 6560
rect 27834 6496 27850 6560
rect 27914 6496 27920 6560
rect 27604 6495 27920 6496
rect 4660 6016 4976 6017
rect 4660 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4976 6016
rect 4660 5951 4976 5952
rect 12088 6016 12404 6017
rect 12088 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12404 6016
rect 12088 5951 12404 5952
rect 19516 6016 19832 6017
rect 19516 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19832 6016
rect 19516 5951 19832 5952
rect 26944 6016 27260 6017
rect 26944 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27260 6016
rect 26944 5951 27260 5952
rect 5320 5472 5636 5473
rect 5320 5408 5326 5472
rect 5390 5408 5406 5472
rect 5470 5408 5486 5472
rect 5550 5408 5566 5472
rect 5630 5408 5636 5472
rect 5320 5407 5636 5408
rect 12748 5472 13064 5473
rect 12748 5408 12754 5472
rect 12818 5408 12834 5472
rect 12898 5408 12914 5472
rect 12978 5408 12994 5472
rect 13058 5408 13064 5472
rect 12748 5407 13064 5408
rect 20176 5472 20492 5473
rect 20176 5408 20182 5472
rect 20246 5408 20262 5472
rect 20326 5408 20342 5472
rect 20406 5408 20422 5472
rect 20486 5408 20492 5472
rect 20176 5407 20492 5408
rect 27604 5472 27920 5473
rect 27604 5408 27610 5472
rect 27674 5408 27690 5472
rect 27754 5408 27770 5472
rect 27834 5408 27850 5472
rect 27914 5408 27920 5472
rect 27604 5407 27920 5408
rect 4660 4928 4976 4929
rect 4660 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4976 4928
rect 4660 4863 4976 4864
rect 12088 4928 12404 4929
rect 12088 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12404 4928
rect 12088 4863 12404 4864
rect 19516 4928 19832 4929
rect 19516 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19832 4928
rect 19516 4863 19832 4864
rect 26944 4928 27260 4929
rect 26944 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27260 4928
rect 26944 4863 27260 4864
rect 5320 4384 5636 4385
rect 5320 4320 5326 4384
rect 5390 4320 5406 4384
rect 5470 4320 5486 4384
rect 5550 4320 5566 4384
rect 5630 4320 5636 4384
rect 5320 4319 5636 4320
rect 12748 4384 13064 4385
rect 12748 4320 12754 4384
rect 12818 4320 12834 4384
rect 12898 4320 12914 4384
rect 12978 4320 12994 4384
rect 13058 4320 13064 4384
rect 12748 4319 13064 4320
rect 20176 4384 20492 4385
rect 20176 4320 20182 4384
rect 20246 4320 20262 4384
rect 20326 4320 20342 4384
rect 20406 4320 20422 4384
rect 20486 4320 20492 4384
rect 20176 4319 20492 4320
rect 27604 4384 27920 4385
rect 27604 4320 27610 4384
rect 27674 4320 27690 4384
rect 27754 4320 27770 4384
rect 27834 4320 27850 4384
rect 27914 4320 27920 4384
rect 27604 4319 27920 4320
rect 4660 3840 4976 3841
rect 4660 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4976 3840
rect 4660 3775 4976 3776
rect 12088 3840 12404 3841
rect 12088 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12404 3840
rect 12088 3775 12404 3776
rect 19516 3840 19832 3841
rect 19516 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19832 3840
rect 19516 3775 19832 3776
rect 26944 3840 27260 3841
rect 26944 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27260 3840
rect 26944 3775 27260 3776
rect 5320 3296 5636 3297
rect 5320 3232 5326 3296
rect 5390 3232 5406 3296
rect 5470 3232 5486 3296
rect 5550 3232 5566 3296
rect 5630 3232 5636 3296
rect 5320 3231 5636 3232
rect 12748 3296 13064 3297
rect 12748 3232 12754 3296
rect 12818 3232 12834 3296
rect 12898 3232 12914 3296
rect 12978 3232 12994 3296
rect 13058 3232 13064 3296
rect 12748 3231 13064 3232
rect 20176 3296 20492 3297
rect 20176 3232 20182 3296
rect 20246 3232 20262 3296
rect 20326 3232 20342 3296
rect 20406 3232 20422 3296
rect 20486 3232 20492 3296
rect 20176 3231 20492 3232
rect 27604 3296 27920 3297
rect 27604 3232 27610 3296
rect 27674 3232 27690 3296
rect 27754 3232 27770 3296
rect 27834 3232 27850 3296
rect 27914 3232 27920 3296
rect 27604 3231 27920 3232
rect 4660 2752 4976 2753
rect 4660 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4976 2752
rect 4660 2687 4976 2688
rect 12088 2752 12404 2753
rect 12088 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12404 2752
rect 12088 2687 12404 2688
rect 19516 2752 19832 2753
rect 19516 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19832 2752
rect 19516 2687 19832 2688
rect 26944 2752 27260 2753
rect 26944 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27260 2752
rect 26944 2687 27260 2688
rect 5320 2208 5636 2209
rect 5320 2144 5326 2208
rect 5390 2144 5406 2208
rect 5470 2144 5486 2208
rect 5550 2144 5566 2208
rect 5630 2144 5636 2208
rect 5320 2143 5636 2144
rect 12748 2208 13064 2209
rect 12748 2144 12754 2208
rect 12818 2144 12834 2208
rect 12898 2144 12914 2208
rect 12978 2144 12994 2208
rect 13058 2144 13064 2208
rect 12748 2143 13064 2144
rect 20176 2208 20492 2209
rect 20176 2144 20182 2208
rect 20246 2144 20262 2208
rect 20326 2144 20342 2208
rect 20406 2144 20422 2208
rect 20486 2144 20492 2208
rect 20176 2143 20492 2144
rect 27604 2208 27920 2209
rect 27604 2144 27610 2208
rect 27674 2144 27690 2208
rect 27754 2144 27770 2208
rect 27834 2144 27850 2208
rect 27914 2144 27920 2208
rect 27604 2143 27920 2144
<< via3 >>
rect 5326 29404 5390 29408
rect 5326 29348 5330 29404
rect 5330 29348 5386 29404
rect 5386 29348 5390 29404
rect 5326 29344 5390 29348
rect 5406 29404 5470 29408
rect 5406 29348 5410 29404
rect 5410 29348 5466 29404
rect 5466 29348 5470 29404
rect 5406 29344 5470 29348
rect 5486 29404 5550 29408
rect 5486 29348 5490 29404
rect 5490 29348 5546 29404
rect 5546 29348 5550 29404
rect 5486 29344 5550 29348
rect 5566 29404 5630 29408
rect 5566 29348 5570 29404
rect 5570 29348 5626 29404
rect 5626 29348 5630 29404
rect 5566 29344 5630 29348
rect 12754 29404 12818 29408
rect 12754 29348 12758 29404
rect 12758 29348 12814 29404
rect 12814 29348 12818 29404
rect 12754 29344 12818 29348
rect 12834 29404 12898 29408
rect 12834 29348 12838 29404
rect 12838 29348 12894 29404
rect 12894 29348 12898 29404
rect 12834 29344 12898 29348
rect 12914 29404 12978 29408
rect 12914 29348 12918 29404
rect 12918 29348 12974 29404
rect 12974 29348 12978 29404
rect 12914 29344 12978 29348
rect 12994 29404 13058 29408
rect 12994 29348 12998 29404
rect 12998 29348 13054 29404
rect 13054 29348 13058 29404
rect 12994 29344 13058 29348
rect 20182 29404 20246 29408
rect 20182 29348 20186 29404
rect 20186 29348 20242 29404
rect 20242 29348 20246 29404
rect 20182 29344 20246 29348
rect 20262 29404 20326 29408
rect 20262 29348 20266 29404
rect 20266 29348 20322 29404
rect 20322 29348 20326 29404
rect 20262 29344 20326 29348
rect 20342 29404 20406 29408
rect 20342 29348 20346 29404
rect 20346 29348 20402 29404
rect 20402 29348 20406 29404
rect 20342 29344 20406 29348
rect 20422 29404 20486 29408
rect 20422 29348 20426 29404
rect 20426 29348 20482 29404
rect 20482 29348 20486 29404
rect 20422 29344 20486 29348
rect 27610 29404 27674 29408
rect 27610 29348 27614 29404
rect 27614 29348 27670 29404
rect 27670 29348 27674 29404
rect 27610 29344 27674 29348
rect 27690 29404 27754 29408
rect 27690 29348 27694 29404
rect 27694 29348 27750 29404
rect 27750 29348 27754 29404
rect 27690 29344 27754 29348
rect 27770 29404 27834 29408
rect 27770 29348 27774 29404
rect 27774 29348 27830 29404
rect 27830 29348 27834 29404
rect 27770 29344 27834 29348
rect 27850 29404 27914 29408
rect 27850 29348 27854 29404
rect 27854 29348 27910 29404
rect 27910 29348 27914 29404
rect 27850 29344 27914 29348
rect 4666 28860 4730 28864
rect 4666 28804 4670 28860
rect 4670 28804 4726 28860
rect 4726 28804 4730 28860
rect 4666 28800 4730 28804
rect 4746 28860 4810 28864
rect 4746 28804 4750 28860
rect 4750 28804 4806 28860
rect 4806 28804 4810 28860
rect 4746 28800 4810 28804
rect 4826 28860 4890 28864
rect 4826 28804 4830 28860
rect 4830 28804 4886 28860
rect 4886 28804 4890 28860
rect 4826 28800 4890 28804
rect 4906 28860 4970 28864
rect 4906 28804 4910 28860
rect 4910 28804 4966 28860
rect 4966 28804 4970 28860
rect 4906 28800 4970 28804
rect 12094 28860 12158 28864
rect 12094 28804 12098 28860
rect 12098 28804 12154 28860
rect 12154 28804 12158 28860
rect 12094 28800 12158 28804
rect 12174 28860 12238 28864
rect 12174 28804 12178 28860
rect 12178 28804 12234 28860
rect 12234 28804 12238 28860
rect 12174 28800 12238 28804
rect 12254 28860 12318 28864
rect 12254 28804 12258 28860
rect 12258 28804 12314 28860
rect 12314 28804 12318 28860
rect 12254 28800 12318 28804
rect 12334 28860 12398 28864
rect 12334 28804 12338 28860
rect 12338 28804 12394 28860
rect 12394 28804 12398 28860
rect 12334 28800 12398 28804
rect 19522 28860 19586 28864
rect 19522 28804 19526 28860
rect 19526 28804 19582 28860
rect 19582 28804 19586 28860
rect 19522 28800 19586 28804
rect 19602 28860 19666 28864
rect 19602 28804 19606 28860
rect 19606 28804 19662 28860
rect 19662 28804 19666 28860
rect 19602 28800 19666 28804
rect 19682 28860 19746 28864
rect 19682 28804 19686 28860
rect 19686 28804 19742 28860
rect 19742 28804 19746 28860
rect 19682 28800 19746 28804
rect 19762 28860 19826 28864
rect 19762 28804 19766 28860
rect 19766 28804 19822 28860
rect 19822 28804 19826 28860
rect 19762 28800 19826 28804
rect 26950 28860 27014 28864
rect 26950 28804 26954 28860
rect 26954 28804 27010 28860
rect 27010 28804 27014 28860
rect 26950 28800 27014 28804
rect 27030 28860 27094 28864
rect 27030 28804 27034 28860
rect 27034 28804 27090 28860
rect 27090 28804 27094 28860
rect 27030 28800 27094 28804
rect 27110 28860 27174 28864
rect 27110 28804 27114 28860
rect 27114 28804 27170 28860
rect 27170 28804 27174 28860
rect 27110 28800 27174 28804
rect 27190 28860 27254 28864
rect 27190 28804 27194 28860
rect 27194 28804 27250 28860
rect 27250 28804 27254 28860
rect 27190 28800 27254 28804
rect 5326 28316 5390 28320
rect 5326 28260 5330 28316
rect 5330 28260 5386 28316
rect 5386 28260 5390 28316
rect 5326 28256 5390 28260
rect 5406 28316 5470 28320
rect 5406 28260 5410 28316
rect 5410 28260 5466 28316
rect 5466 28260 5470 28316
rect 5406 28256 5470 28260
rect 5486 28316 5550 28320
rect 5486 28260 5490 28316
rect 5490 28260 5546 28316
rect 5546 28260 5550 28316
rect 5486 28256 5550 28260
rect 5566 28316 5630 28320
rect 5566 28260 5570 28316
rect 5570 28260 5626 28316
rect 5626 28260 5630 28316
rect 5566 28256 5630 28260
rect 12754 28316 12818 28320
rect 12754 28260 12758 28316
rect 12758 28260 12814 28316
rect 12814 28260 12818 28316
rect 12754 28256 12818 28260
rect 12834 28316 12898 28320
rect 12834 28260 12838 28316
rect 12838 28260 12894 28316
rect 12894 28260 12898 28316
rect 12834 28256 12898 28260
rect 12914 28316 12978 28320
rect 12914 28260 12918 28316
rect 12918 28260 12974 28316
rect 12974 28260 12978 28316
rect 12914 28256 12978 28260
rect 12994 28316 13058 28320
rect 12994 28260 12998 28316
rect 12998 28260 13054 28316
rect 13054 28260 13058 28316
rect 12994 28256 13058 28260
rect 20182 28316 20246 28320
rect 20182 28260 20186 28316
rect 20186 28260 20242 28316
rect 20242 28260 20246 28316
rect 20182 28256 20246 28260
rect 20262 28316 20326 28320
rect 20262 28260 20266 28316
rect 20266 28260 20322 28316
rect 20322 28260 20326 28316
rect 20262 28256 20326 28260
rect 20342 28316 20406 28320
rect 20342 28260 20346 28316
rect 20346 28260 20402 28316
rect 20402 28260 20406 28316
rect 20342 28256 20406 28260
rect 20422 28316 20486 28320
rect 20422 28260 20426 28316
rect 20426 28260 20482 28316
rect 20482 28260 20486 28316
rect 20422 28256 20486 28260
rect 27610 28316 27674 28320
rect 27610 28260 27614 28316
rect 27614 28260 27670 28316
rect 27670 28260 27674 28316
rect 27610 28256 27674 28260
rect 27690 28316 27754 28320
rect 27690 28260 27694 28316
rect 27694 28260 27750 28316
rect 27750 28260 27754 28316
rect 27690 28256 27754 28260
rect 27770 28316 27834 28320
rect 27770 28260 27774 28316
rect 27774 28260 27830 28316
rect 27830 28260 27834 28316
rect 27770 28256 27834 28260
rect 27850 28316 27914 28320
rect 27850 28260 27854 28316
rect 27854 28260 27910 28316
rect 27910 28260 27914 28316
rect 27850 28256 27914 28260
rect 4666 27772 4730 27776
rect 4666 27716 4670 27772
rect 4670 27716 4726 27772
rect 4726 27716 4730 27772
rect 4666 27712 4730 27716
rect 4746 27772 4810 27776
rect 4746 27716 4750 27772
rect 4750 27716 4806 27772
rect 4806 27716 4810 27772
rect 4746 27712 4810 27716
rect 4826 27772 4890 27776
rect 4826 27716 4830 27772
rect 4830 27716 4886 27772
rect 4886 27716 4890 27772
rect 4826 27712 4890 27716
rect 4906 27772 4970 27776
rect 4906 27716 4910 27772
rect 4910 27716 4966 27772
rect 4966 27716 4970 27772
rect 4906 27712 4970 27716
rect 12094 27772 12158 27776
rect 12094 27716 12098 27772
rect 12098 27716 12154 27772
rect 12154 27716 12158 27772
rect 12094 27712 12158 27716
rect 12174 27772 12238 27776
rect 12174 27716 12178 27772
rect 12178 27716 12234 27772
rect 12234 27716 12238 27772
rect 12174 27712 12238 27716
rect 12254 27772 12318 27776
rect 12254 27716 12258 27772
rect 12258 27716 12314 27772
rect 12314 27716 12318 27772
rect 12254 27712 12318 27716
rect 12334 27772 12398 27776
rect 12334 27716 12338 27772
rect 12338 27716 12394 27772
rect 12394 27716 12398 27772
rect 12334 27712 12398 27716
rect 19522 27772 19586 27776
rect 19522 27716 19526 27772
rect 19526 27716 19582 27772
rect 19582 27716 19586 27772
rect 19522 27712 19586 27716
rect 19602 27772 19666 27776
rect 19602 27716 19606 27772
rect 19606 27716 19662 27772
rect 19662 27716 19666 27772
rect 19602 27712 19666 27716
rect 19682 27772 19746 27776
rect 19682 27716 19686 27772
rect 19686 27716 19742 27772
rect 19742 27716 19746 27772
rect 19682 27712 19746 27716
rect 19762 27772 19826 27776
rect 19762 27716 19766 27772
rect 19766 27716 19822 27772
rect 19822 27716 19826 27772
rect 19762 27712 19826 27716
rect 26950 27772 27014 27776
rect 26950 27716 26954 27772
rect 26954 27716 27010 27772
rect 27010 27716 27014 27772
rect 26950 27712 27014 27716
rect 27030 27772 27094 27776
rect 27030 27716 27034 27772
rect 27034 27716 27090 27772
rect 27090 27716 27094 27772
rect 27030 27712 27094 27716
rect 27110 27772 27174 27776
rect 27110 27716 27114 27772
rect 27114 27716 27170 27772
rect 27170 27716 27174 27772
rect 27110 27712 27174 27716
rect 27190 27772 27254 27776
rect 27190 27716 27194 27772
rect 27194 27716 27250 27772
rect 27250 27716 27254 27772
rect 27190 27712 27254 27716
rect 5326 27228 5390 27232
rect 5326 27172 5330 27228
rect 5330 27172 5386 27228
rect 5386 27172 5390 27228
rect 5326 27168 5390 27172
rect 5406 27228 5470 27232
rect 5406 27172 5410 27228
rect 5410 27172 5466 27228
rect 5466 27172 5470 27228
rect 5406 27168 5470 27172
rect 5486 27228 5550 27232
rect 5486 27172 5490 27228
rect 5490 27172 5546 27228
rect 5546 27172 5550 27228
rect 5486 27168 5550 27172
rect 5566 27228 5630 27232
rect 5566 27172 5570 27228
rect 5570 27172 5626 27228
rect 5626 27172 5630 27228
rect 5566 27168 5630 27172
rect 12754 27228 12818 27232
rect 12754 27172 12758 27228
rect 12758 27172 12814 27228
rect 12814 27172 12818 27228
rect 12754 27168 12818 27172
rect 12834 27228 12898 27232
rect 12834 27172 12838 27228
rect 12838 27172 12894 27228
rect 12894 27172 12898 27228
rect 12834 27168 12898 27172
rect 12914 27228 12978 27232
rect 12914 27172 12918 27228
rect 12918 27172 12974 27228
rect 12974 27172 12978 27228
rect 12914 27168 12978 27172
rect 12994 27228 13058 27232
rect 12994 27172 12998 27228
rect 12998 27172 13054 27228
rect 13054 27172 13058 27228
rect 12994 27168 13058 27172
rect 20182 27228 20246 27232
rect 20182 27172 20186 27228
rect 20186 27172 20242 27228
rect 20242 27172 20246 27228
rect 20182 27168 20246 27172
rect 20262 27228 20326 27232
rect 20262 27172 20266 27228
rect 20266 27172 20322 27228
rect 20322 27172 20326 27228
rect 20262 27168 20326 27172
rect 20342 27228 20406 27232
rect 20342 27172 20346 27228
rect 20346 27172 20402 27228
rect 20402 27172 20406 27228
rect 20342 27168 20406 27172
rect 20422 27228 20486 27232
rect 20422 27172 20426 27228
rect 20426 27172 20482 27228
rect 20482 27172 20486 27228
rect 20422 27168 20486 27172
rect 27610 27228 27674 27232
rect 27610 27172 27614 27228
rect 27614 27172 27670 27228
rect 27670 27172 27674 27228
rect 27610 27168 27674 27172
rect 27690 27228 27754 27232
rect 27690 27172 27694 27228
rect 27694 27172 27750 27228
rect 27750 27172 27754 27228
rect 27690 27168 27754 27172
rect 27770 27228 27834 27232
rect 27770 27172 27774 27228
rect 27774 27172 27830 27228
rect 27830 27172 27834 27228
rect 27770 27168 27834 27172
rect 27850 27228 27914 27232
rect 27850 27172 27854 27228
rect 27854 27172 27910 27228
rect 27910 27172 27914 27228
rect 27850 27168 27914 27172
rect 4666 26684 4730 26688
rect 4666 26628 4670 26684
rect 4670 26628 4726 26684
rect 4726 26628 4730 26684
rect 4666 26624 4730 26628
rect 4746 26684 4810 26688
rect 4746 26628 4750 26684
rect 4750 26628 4806 26684
rect 4806 26628 4810 26684
rect 4746 26624 4810 26628
rect 4826 26684 4890 26688
rect 4826 26628 4830 26684
rect 4830 26628 4886 26684
rect 4886 26628 4890 26684
rect 4826 26624 4890 26628
rect 4906 26684 4970 26688
rect 4906 26628 4910 26684
rect 4910 26628 4966 26684
rect 4966 26628 4970 26684
rect 4906 26624 4970 26628
rect 12094 26684 12158 26688
rect 12094 26628 12098 26684
rect 12098 26628 12154 26684
rect 12154 26628 12158 26684
rect 12094 26624 12158 26628
rect 12174 26684 12238 26688
rect 12174 26628 12178 26684
rect 12178 26628 12234 26684
rect 12234 26628 12238 26684
rect 12174 26624 12238 26628
rect 12254 26684 12318 26688
rect 12254 26628 12258 26684
rect 12258 26628 12314 26684
rect 12314 26628 12318 26684
rect 12254 26624 12318 26628
rect 12334 26684 12398 26688
rect 12334 26628 12338 26684
rect 12338 26628 12394 26684
rect 12394 26628 12398 26684
rect 12334 26624 12398 26628
rect 19522 26684 19586 26688
rect 19522 26628 19526 26684
rect 19526 26628 19582 26684
rect 19582 26628 19586 26684
rect 19522 26624 19586 26628
rect 19602 26684 19666 26688
rect 19602 26628 19606 26684
rect 19606 26628 19662 26684
rect 19662 26628 19666 26684
rect 19602 26624 19666 26628
rect 19682 26684 19746 26688
rect 19682 26628 19686 26684
rect 19686 26628 19742 26684
rect 19742 26628 19746 26684
rect 19682 26624 19746 26628
rect 19762 26684 19826 26688
rect 19762 26628 19766 26684
rect 19766 26628 19822 26684
rect 19822 26628 19826 26684
rect 19762 26624 19826 26628
rect 26950 26684 27014 26688
rect 26950 26628 26954 26684
rect 26954 26628 27010 26684
rect 27010 26628 27014 26684
rect 26950 26624 27014 26628
rect 27030 26684 27094 26688
rect 27030 26628 27034 26684
rect 27034 26628 27090 26684
rect 27090 26628 27094 26684
rect 27030 26624 27094 26628
rect 27110 26684 27174 26688
rect 27110 26628 27114 26684
rect 27114 26628 27170 26684
rect 27170 26628 27174 26684
rect 27110 26624 27174 26628
rect 27190 26684 27254 26688
rect 27190 26628 27194 26684
rect 27194 26628 27250 26684
rect 27250 26628 27254 26684
rect 27190 26624 27254 26628
rect 5326 26140 5390 26144
rect 5326 26084 5330 26140
rect 5330 26084 5386 26140
rect 5386 26084 5390 26140
rect 5326 26080 5390 26084
rect 5406 26140 5470 26144
rect 5406 26084 5410 26140
rect 5410 26084 5466 26140
rect 5466 26084 5470 26140
rect 5406 26080 5470 26084
rect 5486 26140 5550 26144
rect 5486 26084 5490 26140
rect 5490 26084 5546 26140
rect 5546 26084 5550 26140
rect 5486 26080 5550 26084
rect 5566 26140 5630 26144
rect 5566 26084 5570 26140
rect 5570 26084 5626 26140
rect 5626 26084 5630 26140
rect 5566 26080 5630 26084
rect 12754 26140 12818 26144
rect 12754 26084 12758 26140
rect 12758 26084 12814 26140
rect 12814 26084 12818 26140
rect 12754 26080 12818 26084
rect 12834 26140 12898 26144
rect 12834 26084 12838 26140
rect 12838 26084 12894 26140
rect 12894 26084 12898 26140
rect 12834 26080 12898 26084
rect 12914 26140 12978 26144
rect 12914 26084 12918 26140
rect 12918 26084 12974 26140
rect 12974 26084 12978 26140
rect 12914 26080 12978 26084
rect 12994 26140 13058 26144
rect 12994 26084 12998 26140
rect 12998 26084 13054 26140
rect 13054 26084 13058 26140
rect 12994 26080 13058 26084
rect 20182 26140 20246 26144
rect 20182 26084 20186 26140
rect 20186 26084 20242 26140
rect 20242 26084 20246 26140
rect 20182 26080 20246 26084
rect 20262 26140 20326 26144
rect 20262 26084 20266 26140
rect 20266 26084 20322 26140
rect 20322 26084 20326 26140
rect 20262 26080 20326 26084
rect 20342 26140 20406 26144
rect 20342 26084 20346 26140
rect 20346 26084 20402 26140
rect 20402 26084 20406 26140
rect 20342 26080 20406 26084
rect 20422 26140 20486 26144
rect 20422 26084 20426 26140
rect 20426 26084 20482 26140
rect 20482 26084 20486 26140
rect 20422 26080 20486 26084
rect 27610 26140 27674 26144
rect 27610 26084 27614 26140
rect 27614 26084 27670 26140
rect 27670 26084 27674 26140
rect 27610 26080 27674 26084
rect 27690 26140 27754 26144
rect 27690 26084 27694 26140
rect 27694 26084 27750 26140
rect 27750 26084 27754 26140
rect 27690 26080 27754 26084
rect 27770 26140 27834 26144
rect 27770 26084 27774 26140
rect 27774 26084 27830 26140
rect 27830 26084 27834 26140
rect 27770 26080 27834 26084
rect 27850 26140 27914 26144
rect 27850 26084 27854 26140
rect 27854 26084 27910 26140
rect 27910 26084 27914 26140
rect 27850 26080 27914 26084
rect 4666 25596 4730 25600
rect 4666 25540 4670 25596
rect 4670 25540 4726 25596
rect 4726 25540 4730 25596
rect 4666 25536 4730 25540
rect 4746 25596 4810 25600
rect 4746 25540 4750 25596
rect 4750 25540 4806 25596
rect 4806 25540 4810 25596
rect 4746 25536 4810 25540
rect 4826 25596 4890 25600
rect 4826 25540 4830 25596
rect 4830 25540 4886 25596
rect 4886 25540 4890 25596
rect 4826 25536 4890 25540
rect 4906 25596 4970 25600
rect 4906 25540 4910 25596
rect 4910 25540 4966 25596
rect 4966 25540 4970 25596
rect 4906 25536 4970 25540
rect 12094 25596 12158 25600
rect 12094 25540 12098 25596
rect 12098 25540 12154 25596
rect 12154 25540 12158 25596
rect 12094 25536 12158 25540
rect 12174 25596 12238 25600
rect 12174 25540 12178 25596
rect 12178 25540 12234 25596
rect 12234 25540 12238 25596
rect 12174 25536 12238 25540
rect 12254 25596 12318 25600
rect 12254 25540 12258 25596
rect 12258 25540 12314 25596
rect 12314 25540 12318 25596
rect 12254 25536 12318 25540
rect 12334 25596 12398 25600
rect 12334 25540 12338 25596
rect 12338 25540 12394 25596
rect 12394 25540 12398 25596
rect 12334 25536 12398 25540
rect 19522 25596 19586 25600
rect 19522 25540 19526 25596
rect 19526 25540 19582 25596
rect 19582 25540 19586 25596
rect 19522 25536 19586 25540
rect 19602 25596 19666 25600
rect 19602 25540 19606 25596
rect 19606 25540 19662 25596
rect 19662 25540 19666 25596
rect 19602 25536 19666 25540
rect 19682 25596 19746 25600
rect 19682 25540 19686 25596
rect 19686 25540 19742 25596
rect 19742 25540 19746 25596
rect 19682 25536 19746 25540
rect 19762 25596 19826 25600
rect 19762 25540 19766 25596
rect 19766 25540 19822 25596
rect 19822 25540 19826 25596
rect 19762 25536 19826 25540
rect 26950 25596 27014 25600
rect 26950 25540 26954 25596
rect 26954 25540 27010 25596
rect 27010 25540 27014 25596
rect 26950 25536 27014 25540
rect 27030 25596 27094 25600
rect 27030 25540 27034 25596
rect 27034 25540 27090 25596
rect 27090 25540 27094 25596
rect 27030 25536 27094 25540
rect 27110 25596 27174 25600
rect 27110 25540 27114 25596
rect 27114 25540 27170 25596
rect 27170 25540 27174 25596
rect 27110 25536 27174 25540
rect 27190 25596 27254 25600
rect 27190 25540 27194 25596
rect 27194 25540 27250 25596
rect 27250 25540 27254 25596
rect 27190 25536 27254 25540
rect 5326 25052 5390 25056
rect 5326 24996 5330 25052
rect 5330 24996 5386 25052
rect 5386 24996 5390 25052
rect 5326 24992 5390 24996
rect 5406 25052 5470 25056
rect 5406 24996 5410 25052
rect 5410 24996 5466 25052
rect 5466 24996 5470 25052
rect 5406 24992 5470 24996
rect 5486 25052 5550 25056
rect 5486 24996 5490 25052
rect 5490 24996 5546 25052
rect 5546 24996 5550 25052
rect 5486 24992 5550 24996
rect 5566 25052 5630 25056
rect 5566 24996 5570 25052
rect 5570 24996 5626 25052
rect 5626 24996 5630 25052
rect 5566 24992 5630 24996
rect 12754 25052 12818 25056
rect 12754 24996 12758 25052
rect 12758 24996 12814 25052
rect 12814 24996 12818 25052
rect 12754 24992 12818 24996
rect 12834 25052 12898 25056
rect 12834 24996 12838 25052
rect 12838 24996 12894 25052
rect 12894 24996 12898 25052
rect 12834 24992 12898 24996
rect 12914 25052 12978 25056
rect 12914 24996 12918 25052
rect 12918 24996 12974 25052
rect 12974 24996 12978 25052
rect 12914 24992 12978 24996
rect 12994 25052 13058 25056
rect 12994 24996 12998 25052
rect 12998 24996 13054 25052
rect 13054 24996 13058 25052
rect 12994 24992 13058 24996
rect 20182 25052 20246 25056
rect 20182 24996 20186 25052
rect 20186 24996 20242 25052
rect 20242 24996 20246 25052
rect 20182 24992 20246 24996
rect 20262 25052 20326 25056
rect 20262 24996 20266 25052
rect 20266 24996 20322 25052
rect 20322 24996 20326 25052
rect 20262 24992 20326 24996
rect 20342 25052 20406 25056
rect 20342 24996 20346 25052
rect 20346 24996 20402 25052
rect 20402 24996 20406 25052
rect 20342 24992 20406 24996
rect 20422 25052 20486 25056
rect 20422 24996 20426 25052
rect 20426 24996 20482 25052
rect 20482 24996 20486 25052
rect 20422 24992 20486 24996
rect 27610 25052 27674 25056
rect 27610 24996 27614 25052
rect 27614 24996 27670 25052
rect 27670 24996 27674 25052
rect 27610 24992 27674 24996
rect 27690 25052 27754 25056
rect 27690 24996 27694 25052
rect 27694 24996 27750 25052
rect 27750 24996 27754 25052
rect 27690 24992 27754 24996
rect 27770 25052 27834 25056
rect 27770 24996 27774 25052
rect 27774 24996 27830 25052
rect 27830 24996 27834 25052
rect 27770 24992 27834 24996
rect 27850 25052 27914 25056
rect 27850 24996 27854 25052
rect 27854 24996 27910 25052
rect 27910 24996 27914 25052
rect 27850 24992 27914 24996
rect 4666 24508 4730 24512
rect 4666 24452 4670 24508
rect 4670 24452 4726 24508
rect 4726 24452 4730 24508
rect 4666 24448 4730 24452
rect 4746 24508 4810 24512
rect 4746 24452 4750 24508
rect 4750 24452 4806 24508
rect 4806 24452 4810 24508
rect 4746 24448 4810 24452
rect 4826 24508 4890 24512
rect 4826 24452 4830 24508
rect 4830 24452 4886 24508
rect 4886 24452 4890 24508
rect 4826 24448 4890 24452
rect 4906 24508 4970 24512
rect 4906 24452 4910 24508
rect 4910 24452 4966 24508
rect 4966 24452 4970 24508
rect 4906 24448 4970 24452
rect 12094 24508 12158 24512
rect 12094 24452 12098 24508
rect 12098 24452 12154 24508
rect 12154 24452 12158 24508
rect 12094 24448 12158 24452
rect 12174 24508 12238 24512
rect 12174 24452 12178 24508
rect 12178 24452 12234 24508
rect 12234 24452 12238 24508
rect 12174 24448 12238 24452
rect 12254 24508 12318 24512
rect 12254 24452 12258 24508
rect 12258 24452 12314 24508
rect 12314 24452 12318 24508
rect 12254 24448 12318 24452
rect 12334 24508 12398 24512
rect 12334 24452 12338 24508
rect 12338 24452 12394 24508
rect 12394 24452 12398 24508
rect 12334 24448 12398 24452
rect 19522 24508 19586 24512
rect 19522 24452 19526 24508
rect 19526 24452 19582 24508
rect 19582 24452 19586 24508
rect 19522 24448 19586 24452
rect 19602 24508 19666 24512
rect 19602 24452 19606 24508
rect 19606 24452 19662 24508
rect 19662 24452 19666 24508
rect 19602 24448 19666 24452
rect 19682 24508 19746 24512
rect 19682 24452 19686 24508
rect 19686 24452 19742 24508
rect 19742 24452 19746 24508
rect 19682 24448 19746 24452
rect 19762 24508 19826 24512
rect 19762 24452 19766 24508
rect 19766 24452 19822 24508
rect 19822 24452 19826 24508
rect 19762 24448 19826 24452
rect 26950 24508 27014 24512
rect 26950 24452 26954 24508
rect 26954 24452 27010 24508
rect 27010 24452 27014 24508
rect 26950 24448 27014 24452
rect 27030 24508 27094 24512
rect 27030 24452 27034 24508
rect 27034 24452 27090 24508
rect 27090 24452 27094 24508
rect 27030 24448 27094 24452
rect 27110 24508 27174 24512
rect 27110 24452 27114 24508
rect 27114 24452 27170 24508
rect 27170 24452 27174 24508
rect 27110 24448 27174 24452
rect 27190 24508 27254 24512
rect 27190 24452 27194 24508
rect 27194 24452 27250 24508
rect 27250 24452 27254 24508
rect 27190 24448 27254 24452
rect 5326 23964 5390 23968
rect 5326 23908 5330 23964
rect 5330 23908 5386 23964
rect 5386 23908 5390 23964
rect 5326 23904 5390 23908
rect 5406 23964 5470 23968
rect 5406 23908 5410 23964
rect 5410 23908 5466 23964
rect 5466 23908 5470 23964
rect 5406 23904 5470 23908
rect 5486 23964 5550 23968
rect 5486 23908 5490 23964
rect 5490 23908 5546 23964
rect 5546 23908 5550 23964
rect 5486 23904 5550 23908
rect 5566 23964 5630 23968
rect 5566 23908 5570 23964
rect 5570 23908 5626 23964
rect 5626 23908 5630 23964
rect 5566 23904 5630 23908
rect 12754 23964 12818 23968
rect 12754 23908 12758 23964
rect 12758 23908 12814 23964
rect 12814 23908 12818 23964
rect 12754 23904 12818 23908
rect 12834 23964 12898 23968
rect 12834 23908 12838 23964
rect 12838 23908 12894 23964
rect 12894 23908 12898 23964
rect 12834 23904 12898 23908
rect 12914 23964 12978 23968
rect 12914 23908 12918 23964
rect 12918 23908 12974 23964
rect 12974 23908 12978 23964
rect 12914 23904 12978 23908
rect 12994 23964 13058 23968
rect 12994 23908 12998 23964
rect 12998 23908 13054 23964
rect 13054 23908 13058 23964
rect 12994 23904 13058 23908
rect 20182 23964 20246 23968
rect 20182 23908 20186 23964
rect 20186 23908 20242 23964
rect 20242 23908 20246 23964
rect 20182 23904 20246 23908
rect 20262 23964 20326 23968
rect 20262 23908 20266 23964
rect 20266 23908 20322 23964
rect 20322 23908 20326 23964
rect 20262 23904 20326 23908
rect 20342 23964 20406 23968
rect 20342 23908 20346 23964
rect 20346 23908 20402 23964
rect 20402 23908 20406 23964
rect 20342 23904 20406 23908
rect 20422 23964 20486 23968
rect 20422 23908 20426 23964
rect 20426 23908 20482 23964
rect 20482 23908 20486 23964
rect 20422 23904 20486 23908
rect 27610 23964 27674 23968
rect 27610 23908 27614 23964
rect 27614 23908 27670 23964
rect 27670 23908 27674 23964
rect 27610 23904 27674 23908
rect 27690 23964 27754 23968
rect 27690 23908 27694 23964
rect 27694 23908 27750 23964
rect 27750 23908 27754 23964
rect 27690 23904 27754 23908
rect 27770 23964 27834 23968
rect 27770 23908 27774 23964
rect 27774 23908 27830 23964
rect 27830 23908 27834 23964
rect 27770 23904 27834 23908
rect 27850 23964 27914 23968
rect 27850 23908 27854 23964
rect 27854 23908 27910 23964
rect 27910 23908 27914 23964
rect 27850 23904 27914 23908
rect 4666 23420 4730 23424
rect 4666 23364 4670 23420
rect 4670 23364 4726 23420
rect 4726 23364 4730 23420
rect 4666 23360 4730 23364
rect 4746 23420 4810 23424
rect 4746 23364 4750 23420
rect 4750 23364 4806 23420
rect 4806 23364 4810 23420
rect 4746 23360 4810 23364
rect 4826 23420 4890 23424
rect 4826 23364 4830 23420
rect 4830 23364 4886 23420
rect 4886 23364 4890 23420
rect 4826 23360 4890 23364
rect 4906 23420 4970 23424
rect 4906 23364 4910 23420
rect 4910 23364 4966 23420
rect 4966 23364 4970 23420
rect 4906 23360 4970 23364
rect 12094 23420 12158 23424
rect 12094 23364 12098 23420
rect 12098 23364 12154 23420
rect 12154 23364 12158 23420
rect 12094 23360 12158 23364
rect 12174 23420 12238 23424
rect 12174 23364 12178 23420
rect 12178 23364 12234 23420
rect 12234 23364 12238 23420
rect 12174 23360 12238 23364
rect 12254 23420 12318 23424
rect 12254 23364 12258 23420
rect 12258 23364 12314 23420
rect 12314 23364 12318 23420
rect 12254 23360 12318 23364
rect 12334 23420 12398 23424
rect 12334 23364 12338 23420
rect 12338 23364 12394 23420
rect 12394 23364 12398 23420
rect 12334 23360 12398 23364
rect 19522 23420 19586 23424
rect 19522 23364 19526 23420
rect 19526 23364 19582 23420
rect 19582 23364 19586 23420
rect 19522 23360 19586 23364
rect 19602 23420 19666 23424
rect 19602 23364 19606 23420
rect 19606 23364 19662 23420
rect 19662 23364 19666 23420
rect 19602 23360 19666 23364
rect 19682 23420 19746 23424
rect 19682 23364 19686 23420
rect 19686 23364 19742 23420
rect 19742 23364 19746 23420
rect 19682 23360 19746 23364
rect 19762 23420 19826 23424
rect 19762 23364 19766 23420
rect 19766 23364 19822 23420
rect 19822 23364 19826 23420
rect 19762 23360 19826 23364
rect 26950 23420 27014 23424
rect 26950 23364 26954 23420
rect 26954 23364 27010 23420
rect 27010 23364 27014 23420
rect 26950 23360 27014 23364
rect 27030 23420 27094 23424
rect 27030 23364 27034 23420
rect 27034 23364 27090 23420
rect 27090 23364 27094 23420
rect 27030 23360 27094 23364
rect 27110 23420 27174 23424
rect 27110 23364 27114 23420
rect 27114 23364 27170 23420
rect 27170 23364 27174 23420
rect 27110 23360 27174 23364
rect 27190 23420 27254 23424
rect 27190 23364 27194 23420
rect 27194 23364 27250 23420
rect 27250 23364 27254 23420
rect 27190 23360 27254 23364
rect 5326 22876 5390 22880
rect 5326 22820 5330 22876
rect 5330 22820 5386 22876
rect 5386 22820 5390 22876
rect 5326 22816 5390 22820
rect 5406 22876 5470 22880
rect 5406 22820 5410 22876
rect 5410 22820 5466 22876
rect 5466 22820 5470 22876
rect 5406 22816 5470 22820
rect 5486 22876 5550 22880
rect 5486 22820 5490 22876
rect 5490 22820 5546 22876
rect 5546 22820 5550 22876
rect 5486 22816 5550 22820
rect 5566 22876 5630 22880
rect 5566 22820 5570 22876
rect 5570 22820 5626 22876
rect 5626 22820 5630 22876
rect 5566 22816 5630 22820
rect 12754 22876 12818 22880
rect 12754 22820 12758 22876
rect 12758 22820 12814 22876
rect 12814 22820 12818 22876
rect 12754 22816 12818 22820
rect 12834 22876 12898 22880
rect 12834 22820 12838 22876
rect 12838 22820 12894 22876
rect 12894 22820 12898 22876
rect 12834 22816 12898 22820
rect 12914 22876 12978 22880
rect 12914 22820 12918 22876
rect 12918 22820 12974 22876
rect 12974 22820 12978 22876
rect 12914 22816 12978 22820
rect 12994 22876 13058 22880
rect 12994 22820 12998 22876
rect 12998 22820 13054 22876
rect 13054 22820 13058 22876
rect 12994 22816 13058 22820
rect 20182 22876 20246 22880
rect 20182 22820 20186 22876
rect 20186 22820 20242 22876
rect 20242 22820 20246 22876
rect 20182 22816 20246 22820
rect 20262 22876 20326 22880
rect 20262 22820 20266 22876
rect 20266 22820 20322 22876
rect 20322 22820 20326 22876
rect 20262 22816 20326 22820
rect 20342 22876 20406 22880
rect 20342 22820 20346 22876
rect 20346 22820 20402 22876
rect 20402 22820 20406 22876
rect 20342 22816 20406 22820
rect 20422 22876 20486 22880
rect 20422 22820 20426 22876
rect 20426 22820 20482 22876
rect 20482 22820 20486 22876
rect 20422 22816 20486 22820
rect 27610 22876 27674 22880
rect 27610 22820 27614 22876
rect 27614 22820 27670 22876
rect 27670 22820 27674 22876
rect 27610 22816 27674 22820
rect 27690 22876 27754 22880
rect 27690 22820 27694 22876
rect 27694 22820 27750 22876
rect 27750 22820 27754 22876
rect 27690 22816 27754 22820
rect 27770 22876 27834 22880
rect 27770 22820 27774 22876
rect 27774 22820 27830 22876
rect 27830 22820 27834 22876
rect 27770 22816 27834 22820
rect 27850 22876 27914 22880
rect 27850 22820 27854 22876
rect 27854 22820 27910 22876
rect 27910 22820 27914 22876
rect 27850 22816 27914 22820
rect 4666 22332 4730 22336
rect 4666 22276 4670 22332
rect 4670 22276 4726 22332
rect 4726 22276 4730 22332
rect 4666 22272 4730 22276
rect 4746 22332 4810 22336
rect 4746 22276 4750 22332
rect 4750 22276 4806 22332
rect 4806 22276 4810 22332
rect 4746 22272 4810 22276
rect 4826 22332 4890 22336
rect 4826 22276 4830 22332
rect 4830 22276 4886 22332
rect 4886 22276 4890 22332
rect 4826 22272 4890 22276
rect 4906 22332 4970 22336
rect 4906 22276 4910 22332
rect 4910 22276 4966 22332
rect 4966 22276 4970 22332
rect 4906 22272 4970 22276
rect 12094 22332 12158 22336
rect 12094 22276 12098 22332
rect 12098 22276 12154 22332
rect 12154 22276 12158 22332
rect 12094 22272 12158 22276
rect 12174 22332 12238 22336
rect 12174 22276 12178 22332
rect 12178 22276 12234 22332
rect 12234 22276 12238 22332
rect 12174 22272 12238 22276
rect 12254 22332 12318 22336
rect 12254 22276 12258 22332
rect 12258 22276 12314 22332
rect 12314 22276 12318 22332
rect 12254 22272 12318 22276
rect 12334 22332 12398 22336
rect 12334 22276 12338 22332
rect 12338 22276 12394 22332
rect 12394 22276 12398 22332
rect 12334 22272 12398 22276
rect 19522 22332 19586 22336
rect 19522 22276 19526 22332
rect 19526 22276 19582 22332
rect 19582 22276 19586 22332
rect 19522 22272 19586 22276
rect 19602 22332 19666 22336
rect 19602 22276 19606 22332
rect 19606 22276 19662 22332
rect 19662 22276 19666 22332
rect 19602 22272 19666 22276
rect 19682 22332 19746 22336
rect 19682 22276 19686 22332
rect 19686 22276 19742 22332
rect 19742 22276 19746 22332
rect 19682 22272 19746 22276
rect 19762 22332 19826 22336
rect 19762 22276 19766 22332
rect 19766 22276 19822 22332
rect 19822 22276 19826 22332
rect 19762 22272 19826 22276
rect 26950 22332 27014 22336
rect 26950 22276 26954 22332
rect 26954 22276 27010 22332
rect 27010 22276 27014 22332
rect 26950 22272 27014 22276
rect 27030 22332 27094 22336
rect 27030 22276 27034 22332
rect 27034 22276 27090 22332
rect 27090 22276 27094 22332
rect 27030 22272 27094 22276
rect 27110 22332 27174 22336
rect 27110 22276 27114 22332
rect 27114 22276 27170 22332
rect 27170 22276 27174 22332
rect 27110 22272 27174 22276
rect 27190 22332 27254 22336
rect 27190 22276 27194 22332
rect 27194 22276 27250 22332
rect 27250 22276 27254 22332
rect 27190 22272 27254 22276
rect 5326 21788 5390 21792
rect 5326 21732 5330 21788
rect 5330 21732 5386 21788
rect 5386 21732 5390 21788
rect 5326 21728 5390 21732
rect 5406 21788 5470 21792
rect 5406 21732 5410 21788
rect 5410 21732 5466 21788
rect 5466 21732 5470 21788
rect 5406 21728 5470 21732
rect 5486 21788 5550 21792
rect 5486 21732 5490 21788
rect 5490 21732 5546 21788
rect 5546 21732 5550 21788
rect 5486 21728 5550 21732
rect 5566 21788 5630 21792
rect 5566 21732 5570 21788
rect 5570 21732 5626 21788
rect 5626 21732 5630 21788
rect 5566 21728 5630 21732
rect 12754 21788 12818 21792
rect 12754 21732 12758 21788
rect 12758 21732 12814 21788
rect 12814 21732 12818 21788
rect 12754 21728 12818 21732
rect 12834 21788 12898 21792
rect 12834 21732 12838 21788
rect 12838 21732 12894 21788
rect 12894 21732 12898 21788
rect 12834 21728 12898 21732
rect 12914 21788 12978 21792
rect 12914 21732 12918 21788
rect 12918 21732 12974 21788
rect 12974 21732 12978 21788
rect 12914 21728 12978 21732
rect 12994 21788 13058 21792
rect 12994 21732 12998 21788
rect 12998 21732 13054 21788
rect 13054 21732 13058 21788
rect 12994 21728 13058 21732
rect 20182 21788 20246 21792
rect 20182 21732 20186 21788
rect 20186 21732 20242 21788
rect 20242 21732 20246 21788
rect 20182 21728 20246 21732
rect 20262 21788 20326 21792
rect 20262 21732 20266 21788
rect 20266 21732 20322 21788
rect 20322 21732 20326 21788
rect 20262 21728 20326 21732
rect 20342 21788 20406 21792
rect 20342 21732 20346 21788
rect 20346 21732 20402 21788
rect 20402 21732 20406 21788
rect 20342 21728 20406 21732
rect 20422 21788 20486 21792
rect 20422 21732 20426 21788
rect 20426 21732 20482 21788
rect 20482 21732 20486 21788
rect 20422 21728 20486 21732
rect 27610 21788 27674 21792
rect 27610 21732 27614 21788
rect 27614 21732 27670 21788
rect 27670 21732 27674 21788
rect 27610 21728 27674 21732
rect 27690 21788 27754 21792
rect 27690 21732 27694 21788
rect 27694 21732 27750 21788
rect 27750 21732 27754 21788
rect 27690 21728 27754 21732
rect 27770 21788 27834 21792
rect 27770 21732 27774 21788
rect 27774 21732 27830 21788
rect 27830 21732 27834 21788
rect 27770 21728 27834 21732
rect 27850 21788 27914 21792
rect 27850 21732 27854 21788
rect 27854 21732 27910 21788
rect 27910 21732 27914 21788
rect 27850 21728 27914 21732
rect 4666 21244 4730 21248
rect 4666 21188 4670 21244
rect 4670 21188 4726 21244
rect 4726 21188 4730 21244
rect 4666 21184 4730 21188
rect 4746 21244 4810 21248
rect 4746 21188 4750 21244
rect 4750 21188 4806 21244
rect 4806 21188 4810 21244
rect 4746 21184 4810 21188
rect 4826 21244 4890 21248
rect 4826 21188 4830 21244
rect 4830 21188 4886 21244
rect 4886 21188 4890 21244
rect 4826 21184 4890 21188
rect 4906 21244 4970 21248
rect 4906 21188 4910 21244
rect 4910 21188 4966 21244
rect 4966 21188 4970 21244
rect 4906 21184 4970 21188
rect 12094 21244 12158 21248
rect 12094 21188 12098 21244
rect 12098 21188 12154 21244
rect 12154 21188 12158 21244
rect 12094 21184 12158 21188
rect 12174 21244 12238 21248
rect 12174 21188 12178 21244
rect 12178 21188 12234 21244
rect 12234 21188 12238 21244
rect 12174 21184 12238 21188
rect 12254 21244 12318 21248
rect 12254 21188 12258 21244
rect 12258 21188 12314 21244
rect 12314 21188 12318 21244
rect 12254 21184 12318 21188
rect 12334 21244 12398 21248
rect 12334 21188 12338 21244
rect 12338 21188 12394 21244
rect 12394 21188 12398 21244
rect 12334 21184 12398 21188
rect 19522 21244 19586 21248
rect 19522 21188 19526 21244
rect 19526 21188 19582 21244
rect 19582 21188 19586 21244
rect 19522 21184 19586 21188
rect 19602 21244 19666 21248
rect 19602 21188 19606 21244
rect 19606 21188 19662 21244
rect 19662 21188 19666 21244
rect 19602 21184 19666 21188
rect 19682 21244 19746 21248
rect 19682 21188 19686 21244
rect 19686 21188 19742 21244
rect 19742 21188 19746 21244
rect 19682 21184 19746 21188
rect 19762 21244 19826 21248
rect 19762 21188 19766 21244
rect 19766 21188 19822 21244
rect 19822 21188 19826 21244
rect 19762 21184 19826 21188
rect 26950 21244 27014 21248
rect 26950 21188 26954 21244
rect 26954 21188 27010 21244
rect 27010 21188 27014 21244
rect 26950 21184 27014 21188
rect 27030 21244 27094 21248
rect 27030 21188 27034 21244
rect 27034 21188 27090 21244
rect 27090 21188 27094 21244
rect 27030 21184 27094 21188
rect 27110 21244 27174 21248
rect 27110 21188 27114 21244
rect 27114 21188 27170 21244
rect 27170 21188 27174 21244
rect 27110 21184 27174 21188
rect 27190 21244 27254 21248
rect 27190 21188 27194 21244
rect 27194 21188 27250 21244
rect 27250 21188 27254 21244
rect 27190 21184 27254 21188
rect 5326 20700 5390 20704
rect 5326 20644 5330 20700
rect 5330 20644 5386 20700
rect 5386 20644 5390 20700
rect 5326 20640 5390 20644
rect 5406 20700 5470 20704
rect 5406 20644 5410 20700
rect 5410 20644 5466 20700
rect 5466 20644 5470 20700
rect 5406 20640 5470 20644
rect 5486 20700 5550 20704
rect 5486 20644 5490 20700
rect 5490 20644 5546 20700
rect 5546 20644 5550 20700
rect 5486 20640 5550 20644
rect 5566 20700 5630 20704
rect 5566 20644 5570 20700
rect 5570 20644 5626 20700
rect 5626 20644 5630 20700
rect 5566 20640 5630 20644
rect 12754 20700 12818 20704
rect 12754 20644 12758 20700
rect 12758 20644 12814 20700
rect 12814 20644 12818 20700
rect 12754 20640 12818 20644
rect 12834 20700 12898 20704
rect 12834 20644 12838 20700
rect 12838 20644 12894 20700
rect 12894 20644 12898 20700
rect 12834 20640 12898 20644
rect 12914 20700 12978 20704
rect 12914 20644 12918 20700
rect 12918 20644 12974 20700
rect 12974 20644 12978 20700
rect 12914 20640 12978 20644
rect 12994 20700 13058 20704
rect 12994 20644 12998 20700
rect 12998 20644 13054 20700
rect 13054 20644 13058 20700
rect 12994 20640 13058 20644
rect 20182 20700 20246 20704
rect 20182 20644 20186 20700
rect 20186 20644 20242 20700
rect 20242 20644 20246 20700
rect 20182 20640 20246 20644
rect 20262 20700 20326 20704
rect 20262 20644 20266 20700
rect 20266 20644 20322 20700
rect 20322 20644 20326 20700
rect 20262 20640 20326 20644
rect 20342 20700 20406 20704
rect 20342 20644 20346 20700
rect 20346 20644 20402 20700
rect 20402 20644 20406 20700
rect 20342 20640 20406 20644
rect 20422 20700 20486 20704
rect 20422 20644 20426 20700
rect 20426 20644 20482 20700
rect 20482 20644 20486 20700
rect 20422 20640 20486 20644
rect 27610 20700 27674 20704
rect 27610 20644 27614 20700
rect 27614 20644 27670 20700
rect 27670 20644 27674 20700
rect 27610 20640 27674 20644
rect 27690 20700 27754 20704
rect 27690 20644 27694 20700
rect 27694 20644 27750 20700
rect 27750 20644 27754 20700
rect 27690 20640 27754 20644
rect 27770 20700 27834 20704
rect 27770 20644 27774 20700
rect 27774 20644 27830 20700
rect 27830 20644 27834 20700
rect 27770 20640 27834 20644
rect 27850 20700 27914 20704
rect 27850 20644 27854 20700
rect 27854 20644 27910 20700
rect 27910 20644 27914 20700
rect 27850 20640 27914 20644
rect 4666 20156 4730 20160
rect 4666 20100 4670 20156
rect 4670 20100 4726 20156
rect 4726 20100 4730 20156
rect 4666 20096 4730 20100
rect 4746 20156 4810 20160
rect 4746 20100 4750 20156
rect 4750 20100 4806 20156
rect 4806 20100 4810 20156
rect 4746 20096 4810 20100
rect 4826 20156 4890 20160
rect 4826 20100 4830 20156
rect 4830 20100 4886 20156
rect 4886 20100 4890 20156
rect 4826 20096 4890 20100
rect 4906 20156 4970 20160
rect 4906 20100 4910 20156
rect 4910 20100 4966 20156
rect 4966 20100 4970 20156
rect 4906 20096 4970 20100
rect 12094 20156 12158 20160
rect 12094 20100 12098 20156
rect 12098 20100 12154 20156
rect 12154 20100 12158 20156
rect 12094 20096 12158 20100
rect 12174 20156 12238 20160
rect 12174 20100 12178 20156
rect 12178 20100 12234 20156
rect 12234 20100 12238 20156
rect 12174 20096 12238 20100
rect 12254 20156 12318 20160
rect 12254 20100 12258 20156
rect 12258 20100 12314 20156
rect 12314 20100 12318 20156
rect 12254 20096 12318 20100
rect 12334 20156 12398 20160
rect 12334 20100 12338 20156
rect 12338 20100 12394 20156
rect 12394 20100 12398 20156
rect 12334 20096 12398 20100
rect 19522 20156 19586 20160
rect 19522 20100 19526 20156
rect 19526 20100 19582 20156
rect 19582 20100 19586 20156
rect 19522 20096 19586 20100
rect 19602 20156 19666 20160
rect 19602 20100 19606 20156
rect 19606 20100 19662 20156
rect 19662 20100 19666 20156
rect 19602 20096 19666 20100
rect 19682 20156 19746 20160
rect 19682 20100 19686 20156
rect 19686 20100 19742 20156
rect 19742 20100 19746 20156
rect 19682 20096 19746 20100
rect 19762 20156 19826 20160
rect 19762 20100 19766 20156
rect 19766 20100 19822 20156
rect 19822 20100 19826 20156
rect 19762 20096 19826 20100
rect 26950 20156 27014 20160
rect 26950 20100 26954 20156
rect 26954 20100 27010 20156
rect 27010 20100 27014 20156
rect 26950 20096 27014 20100
rect 27030 20156 27094 20160
rect 27030 20100 27034 20156
rect 27034 20100 27090 20156
rect 27090 20100 27094 20156
rect 27030 20096 27094 20100
rect 27110 20156 27174 20160
rect 27110 20100 27114 20156
rect 27114 20100 27170 20156
rect 27170 20100 27174 20156
rect 27110 20096 27174 20100
rect 27190 20156 27254 20160
rect 27190 20100 27194 20156
rect 27194 20100 27250 20156
rect 27250 20100 27254 20156
rect 27190 20096 27254 20100
rect 5326 19612 5390 19616
rect 5326 19556 5330 19612
rect 5330 19556 5386 19612
rect 5386 19556 5390 19612
rect 5326 19552 5390 19556
rect 5406 19612 5470 19616
rect 5406 19556 5410 19612
rect 5410 19556 5466 19612
rect 5466 19556 5470 19612
rect 5406 19552 5470 19556
rect 5486 19612 5550 19616
rect 5486 19556 5490 19612
rect 5490 19556 5546 19612
rect 5546 19556 5550 19612
rect 5486 19552 5550 19556
rect 5566 19612 5630 19616
rect 5566 19556 5570 19612
rect 5570 19556 5626 19612
rect 5626 19556 5630 19612
rect 5566 19552 5630 19556
rect 12754 19612 12818 19616
rect 12754 19556 12758 19612
rect 12758 19556 12814 19612
rect 12814 19556 12818 19612
rect 12754 19552 12818 19556
rect 12834 19612 12898 19616
rect 12834 19556 12838 19612
rect 12838 19556 12894 19612
rect 12894 19556 12898 19612
rect 12834 19552 12898 19556
rect 12914 19612 12978 19616
rect 12914 19556 12918 19612
rect 12918 19556 12974 19612
rect 12974 19556 12978 19612
rect 12914 19552 12978 19556
rect 12994 19612 13058 19616
rect 12994 19556 12998 19612
rect 12998 19556 13054 19612
rect 13054 19556 13058 19612
rect 12994 19552 13058 19556
rect 20182 19612 20246 19616
rect 20182 19556 20186 19612
rect 20186 19556 20242 19612
rect 20242 19556 20246 19612
rect 20182 19552 20246 19556
rect 20262 19612 20326 19616
rect 20262 19556 20266 19612
rect 20266 19556 20322 19612
rect 20322 19556 20326 19612
rect 20262 19552 20326 19556
rect 20342 19612 20406 19616
rect 20342 19556 20346 19612
rect 20346 19556 20402 19612
rect 20402 19556 20406 19612
rect 20342 19552 20406 19556
rect 20422 19612 20486 19616
rect 20422 19556 20426 19612
rect 20426 19556 20482 19612
rect 20482 19556 20486 19612
rect 20422 19552 20486 19556
rect 27610 19612 27674 19616
rect 27610 19556 27614 19612
rect 27614 19556 27670 19612
rect 27670 19556 27674 19612
rect 27610 19552 27674 19556
rect 27690 19612 27754 19616
rect 27690 19556 27694 19612
rect 27694 19556 27750 19612
rect 27750 19556 27754 19612
rect 27690 19552 27754 19556
rect 27770 19612 27834 19616
rect 27770 19556 27774 19612
rect 27774 19556 27830 19612
rect 27830 19556 27834 19612
rect 27770 19552 27834 19556
rect 27850 19612 27914 19616
rect 27850 19556 27854 19612
rect 27854 19556 27910 19612
rect 27910 19556 27914 19612
rect 27850 19552 27914 19556
rect 4666 19068 4730 19072
rect 4666 19012 4670 19068
rect 4670 19012 4726 19068
rect 4726 19012 4730 19068
rect 4666 19008 4730 19012
rect 4746 19068 4810 19072
rect 4746 19012 4750 19068
rect 4750 19012 4806 19068
rect 4806 19012 4810 19068
rect 4746 19008 4810 19012
rect 4826 19068 4890 19072
rect 4826 19012 4830 19068
rect 4830 19012 4886 19068
rect 4886 19012 4890 19068
rect 4826 19008 4890 19012
rect 4906 19068 4970 19072
rect 4906 19012 4910 19068
rect 4910 19012 4966 19068
rect 4966 19012 4970 19068
rect 4906 19008 4970 19012
rect 12094 19068 12158 19072
rect 12094 19012 12098 19068
rect 12098 19012 12154 19068
rect 12154 19012 12158 19068
rect 12094 19008 12158 19012
rect 12174 19068 12238 19072
rect 12174 19012 12178 19068
rect 12178 19012 12234 19068
rect 12234 19012 12238 19068
rect 12174 19008 12238 19012
rect 12254 19068 12318 19072
rect 12254 19012 12258 19068
rect 12258 19012 12314 19068
rect 12314 19012 12318 19068
rect 12254 19008 12318 19012
rect 12334 19068 12398 19072
rect 12334 19012 12338 19068
rect 12338 19012 12394 19068
rect 12394 19012 12398 19068
rect 12334 19008 12398 19012
rect 19522 19068 19586 19072
rect 19522 19012 19526 19068
rect 19526 19012 19582 19068
rect 19582 19012 19586 19068
rect 19522 19008 19586 19012
rect 19602 19068 19666 19072
rect 19602 19012 19606 19068
rect 19606 19012 19662 19068
rect 19662 19012 19666 19068
rect 19602 19008 19666 19012
rect 19682 19068 19746 19072
rect 19682 19012 19686 19068
rect 19686 19012 19742 19068
rect 19742 19012 19746 19068
rect 19682 19008 19746 19012
rect 19762 19068 19826 19072
rect 19762 19012 19766 19068
rect 19766 19012 19822 19068
rect 19822 19012 19826 19068
rect 19762 19008 19826 19012
rect 26950 19068 27014 19072
rect 26950 19012 26954 19068
rect 26954 19012 27010 19068
rect 27010 19012 27014 19068
rect 26950 19008 27014 19012
rect 27030 19068 27094 19072
rect 27030 19012 27034 19068
rect 27034 19012 27090 19068
rect 27090 19012 27094 19068
rect 27030 19008 27094 19012
rect 27110 19068 27174 19072
rect 27110 19012 27114 19068
rect 27114 19012 27170 19068
rect 27170 19012 27174 19068
rect 27110 19008 27174 19012
rect 27190 19068 27254 19072
rect 27190 19012 27194 19068
rect 27194 19012 27250 19068
rect 27250 19012 27254 19068
rect 27190 19008 27254 19012
rect 5326 18524 5390 18528
rect 5326 18468 5330 18524
rect 5330 18468 5386 18524
rect 5386 18468 5390 18524
rect 5326 18464 5390 18468
rect 5406 18524 5470 18528
rect 5406 18468 5410 18524
rect 5410 18468 5466 18524
rect 5466 18468 5470 18524
rect 5406 18464 5470 18468
rect 5486 18524 5550 18528
rect 5486 18468 5490 18524
rect 5490 18468 5546 18524
rect 5546 18468 5550 18524
rect 5486 18464 5550 18468
rect 5566 18524 5630 18528
rect 5566 18468 5570 18524
rect 5570 18468 5626 18524
rect 5626 18468 5630 18524
rect 5566 18464 5630 18468
rect 12754 18524 12818 18528
rect 12754 18468 12758 18524
rect 12758 18468 12814 18524
rect 12814 18468 12818 18524
rect 12754 18464 12818 18468
rect 12834 18524 12898 18528
rect 12834 18468 12838 18524
rect 12838 18468 12894 18524
rect 12894 18468 12898 18524
rect 12834 18464 12898 18468
rect 12914 18524 12978 18528
rect 12914 18468 12918 18524
rect 12918 18468 12974 18524
rect 12974 18468 12978 18524
rect 12914 18464 12978 18468
rect 12994 18524 13058 18528
rect 12994 18468 12998 18524
rect 12998 18468 13054 18524
rect 13054 18468 13058 18524
rect 12994 18464 13058 18468
rect 20182 18524 20246 18528
rect 20182 18468 20186 18524
rect 20186 18468 20242 18524
rect 20242 18468 20246 18524
rect 20182 18464 20246 18468
rect 20262 18524 20326 18528
rect 20262 18468 20266 18524
rect 20266 18468 20322 18524
rect 20322 18468 20326 18524
rect 20262 18464 20326 18468
rect 20342 18524 20406 18528
rect 20342 18468 20346 18524
rect 20346 18468 20402 18524
rect 20402 18468 20406 18524
rect 20342 18464 20406 18468
rect 20422 18524 20486 18528
rect 20422 18468 20426 18524
rect 20426 18468 20482 18524
rect 20482 18468 20486 18524
rect 20422 18464 20486 18468
rect 27610 18524 27674 18528
rect 27610 18468 27614 18524
rect 27614 18468 27670 18524
rect 27670 18468 27674 18524
rect 27610 18464 27674 18468
rect 27690 18524 27754 18528
rect 27690 18468 27694 18524
rect 27694 18468 27750 18524
rect 27750 18468 27754 18524
rect 27690 18464 27754 18468
rect 27770 18524 27834 18528
rect 27770 18468 27774 18524
rect 27774 18468 27830 18524
rect 27830 18468 27834 18524
rect 27770 18464 27834 18468
rect 27850 18524 27914 18528
rect 27850 18468 27854 18524
rect 27854 18468 27910 18524
rect 27910 18468 27914 18524
rect 27850 18464 27914 18468
rect 4666 17980 4730 17984
rect 4666 17924 4670 17980
rect 4670 17924 4726 17980
rect 4726 17924 4730 17980
rect 4666 17920 4730 17924
rect 4746 17980 4810 17984
rect 4746 17924 4750 17980
rect 4750 17924 4806 17980
rect 4806 17924 4810 17980
rect 4746 17920 4810 17924
rect 4826 17980 4890 17984
rect 4826 17924 4830 17980
rect 4830 17924 4886 17980
rect 4886 17924 4890 17980
rect 4826 17920 4890 17924
rect 4906 17980 4970 17984
rect 4906 17924 4910 17980
rect 4910 17924 4966 17980
rect 4966 17924 4970 17980
rect 4906 17920 4970 17924
rect 12094 17980 12158 17984
rect 12094 17924 12098 17980
rect 12098 17924 12154 17980
rect 12154 17924 12158 17980
rect 12094 17920 12158 17924
rect 12174 17980 12238 17984
rect 12174 17924 12178 17980
rect 12178 17924 12234 17980
rect 12234 17924 12238 17980
rect 12174 17920 12238 17924
rect 12254 17980 12318 17984
rect 12254 17924 12258 17980
rect 12258 17924 12314 17980
rect 12314 17924 12318 17980
rect 12254 17920 12318 17924
rect 12334 17980 12398 17984
rect 12334 17924 12338 17980
rect 12338 17924 12394 17980
rect 12394 17924 12398 17980
rect 12334 17920 12398 17924
rect 19522 17980 19586 17984
rect 19522 17924 19526 17980
rect 19526 17924 19582 17980
rect 19582 17924 19586 17980
rect 19522 17920 19586 17924
rect 19602 17980 19666 17984
rect 19602 17924 19606 17980
rect 19606 17924 19662 17980
rect 19662 17924 19666 17980
rect 19602 17920 19666 17924
rect 19682 17980 19746 17984
rect 19682 17924 19686 17980
rect 19686 17924 19742 17980
rect 19742 17924 19746 17980
rect 19682 17920 19746 17924
rect 19762 17980 19826 17984
rect 19762 17924 19766 17980
rect 19766 17924 19822 17980
rect 19822 17924 19826 17980
rect 19762 17920 19826 17924
rect 26950 17980 27014 17984
rect 26950 17924 26954 17980
rect 26954 17924 27010 17980
rect 27010 17924 27014 17980
rect 26950 17920 27014 17924
rect 27030 17980 27094 17984
rect 27030 17924 27034 17980
rect 27034 17924 27090 17980
rect 27090 17924 27094 17980
rect 27030 17920 27094 17924
rect 27110 17980 27174 17984
rect 27110 17924 27114 17980
rect 27114 17924 27170 17980
rect 27170 17924 27174 17980
rect 27110 17920 27174 17924
rect 27190 17980 27254 17984
rect 27190 17924 27194 17980
rect 27194 17924 27250 17980
rect 27250 17924 27254 17980
rect 27190 17920 27254 17924
rect 5326 17436 5390 17440
rect 5326 17380 5330 17436
rect 5330 17380 5386 17436
rect 5386 17380 5390 17436
rect 5326 17376 5390 17380
rect 5406 17436 5470 17440
rect 5406 17380 5410 17436
rect 5410 17380 5466 17436
rect 5466 17380 5470 17436
rect 5406 17376 5470 17380
rect 5486 17436 5550 17440
rect 5486 17380 5490 17436
rect 5490 17380 5546 17436
rect 5546 17380 5550 17436
rect 5486 17376 5550 17380
rect 5566 17436 5630 17440
rect 5566 17380 5570 17436
rect 5570 17380 5626 17436
rect 5626 17380 5630 17436
rect 5566 17376 5630 17380
rect 12754 17436 12818 17440
rect 12754 17380 12758 17436
rect 12758 17380 12814 17436
rect 12814 17380 12818 17436
rect 12754 17376 12818 17380
rect 12834 17436 12898 17440
rect 12834 17380 12838 17436
rect 12838 17380 12894 17436
rect 12894 17380 12898 17436
rect 12834 17376 12898 17380
rect 12914 17436 12978 17440
rect 12914 17380 12918 17436
rect 12918 17380 12974 17436
rect 12974 17380 12978 17436
rect 12914 17376 12978 17380
rect 12994 17436 13058 17440
rect 12994 17380 12998 17436
rect 12998 17380 13054 17436
rect 13054 17380 13058 17436
rect 12994 17376 13058 17380
rect 20182 17436 20246 17440
rect 20182 17380 20186 17436
rect 20186 17380 20242 17436
rect 20242 17380 20246 17436
rect 20182 17376 20246 17380
rect 20262 17436 20326 17440
rect 20262 17380 20266 17436
rect 20266 17380 20322 17436
rect 20322 17380 20326 17436
rect 20262 17376 20326 17380
rect 20342 17436 20406 17440
rect 20342 17380 20346 17436
rect 20346 17380 20402 17436
rect 20402 17380 20406 17436
rect 20342 17376 20406 17380
rect 20422 17436 20486 17440
rect 20422 17380 20426 17436
rect 20426 17380 20482 17436
rect 20482 17380 20486 17436
rect 20422 17376 20486 17380
rect 27610 17436 27674 17440
rect 27610 17380 27614 17436
rect 27614 17380 27670 17436
rect 27670 17380 27674 17436
rect 27610 17376 27674 17380
rect 27690 17436 27754 17440
rect 27690 17380 27694 17436
rect 27694 17380 27750 17436
rect 27750 17380 27754 17436
rect 27690 17376 27754 17380
rect 27770 17436 27834 17440
rect 27770 17380 27774 17436
rect 27774 17380 27830 17436
rect 27830 17380 27834 17436
rect 27770 17376 27834 17380
rect 27850 17436 27914 17440
rect 27850 17380 27854 17436
rect 27854 17380 27910 17436
rect 27910 17380 27914 17436
rect 27850 17376 27914 17380
rect 4666 16892 4730 16896
rect 4666 16836 4670 16892
rect 4670 16836 4726 16892
rect 4726 16836 4730 16892
rect 4666 16832 4730 16836
rect 4746 16892 4810 16896
rect 4746 16836 4750 16892
rect 4750 16836 4806 16892
rect 4806 16836 4810 16892
rect 4746 16832 4810 16836
rect 4826 16892 4890 16896
rect 4826 16836 4830 16892
rect 4830 16836 4886 16892
rect 4886 16836 4890 16892
rect 4826 16832 4890 16836
rect 4906 16892 4970 16896
rect 4906 16836 4910 16892
rect 4910 16836 4966 16892
rect 4966 16836 4970 16892
rect 4906 16832 4970 16836
rect 12094 16892 12158 16896
rect 12094 16836 12098 16892
rect 12098 16836 12154 16892
rect 12154 16836 12158 16892
rect 12094 16832 12158 16836
rect 12174 16892 12238 16896
rect 12174 16836 12178 16892
rect 12178 16836 12234 16892
rect 12234 16836 12238 16892
rect 12174 16832 12238 16836
rect 12254 16892 12318 16896
rect 12254 16836 12258 16892
rect 12258 16836 12314 16892
rect 12314 16836 12318 16892
rect 12254 16832 12318 16836
rect 12334 16892 12398 16896
rect 12334 16836 12338 16892
rect 12338 16836 12394 16892
rect 12394 16836 12398 16892
rect 12334 16832 12398 16836
rect 19522 16892 19586 16896
rect 19522 16836 19526 16892
rect 19526 16836 19582 16892
rect 19582 16836 19586 16892
rect 19522 16832 19586 16836
rect 19602 16892 19666 16896
rect 19602 16836 19606 16892
rect 19606 16836 19662 16892
rect 19662 16836 19666 16892
rect 19602 16832 19666 16836
rect 19682 16892 19746 16896
rect 19682 16836 19686 16892
rect 19686 16836 19742 16892
rect 19742 16836 19746 16892
rect 19682 16832 19746 16836
rect 19762 16892 19826 16896
rect 19762 16836 19766 16892
rect 19766 16836 19822 16892
rect 19822 16836 19826 16892
rect 19762 16832 19826 16836
rect 26950 16892 27014 16896
rect 26950 16836 26954 16892
rect 26954 16836 27010 16892
rect 27010 16836 27014 16892
rect 26950 16832 27014 16836
rect 27030 16892 27094 16896
rect 27030 16836 27034 16892
rect 27034 16836 27090 16892
rect 27090 16836 27094 16892
rect 27030 16832 27094 16836
rect 27110 16892 27174 16896
rect 27110 16836 27114 16892
rect 27114 16836 27170 16892
rect 27170 16836 27174 16892
rect 27110 16832 27174 16836
rect 27190 16892 27254 16896
rect 27190 16836 27194 16892
rect 27194 16836 27250 16892
rect 27250 16836 27254 16892
rect 27190 16832 27254 16836
rect 5326 16348 5390 16352
rect 5326 16292 5330 16348
rect 5330 16292 5386 16348
rect 5386 16292 5390 16348
rect 5326 16288 5390 16292
rect 5406 16348 5470 16352
rect 5406 16292 5410 16348
rect 5410 16292 5466 16348
rect 5466 16292 5470 16348
rect 5406 16288 5470 16292
rect 5486 16348 5550 16352
rect 5486 16292 5490 16348
rect 5490 16292 5546 16348
rect 5546 16292 5550 16348
rect 5486 16288 5550 16292
rect 5566 16348 5630 16352
rect 5566 16292 5570 16348
rect 5570 16292 5626 16348
rect 5626 16292 5630 16348
rect 5566 16288 5630 16292
rect 12754 16348 12818 16352
rect 12754 16292 12758 16348
rect 12758 16292 12814 16348
rect 12814 16292 12818 16348
rect 12754 16288 12818 16292
rect 12834 16348 12898 16352
rect 12834 16292 12838 16348
rect 12838 16292 12894 16348
rect 12894 16292 12898 16348
rect 12834 16288 12898 16292
rect 12914 16348 12978 16352
rect 12914 16292 12918 16348
rect 12918 16292 12974 16348
rect 12974 16292 12978 16348
rect 12914 16288 12978 16292
rect 12994 16348 13058 16352
rect 12994 16292 12998 16348
rect 12998 16292 13054 16348
rect 13054 16292 13058 16348
rect 12994 16288 13058 16292
rect 20182 16348 20246 16352
rect 20182 16292 20186 16348
rect 20186 16292 20242 16348
rect 20242 16292 20246 16348
rect 20182 16288 20246 16292
rect 20262 16348 20326 16352
rect 20262 16292 20266 16348
rect 20266 16292 20322 16348
rect 20322 16292 20326 16348
rect 20262 16288 20326 16292
rect 20342 16348 20406 16352
rect 20342 16292 20346 16348
rect 20346 16292 20402 16348
rect 20402 16292 20406 16348
rect 20342 16288 20406 16292
rect 20422 16348 20486 16352
rect 20422 16292 20426 16348
rect 20426 16292 20482 16348
rect 20482 16292 20486 16348
rect 20422 16288 20486 16292
rect 27610 16348 27674 16352
rect 27610 16292 27614 16348
rect 27614 16292 27670 16348
rect 27670 16292 27674 16348
rect 27610 16288 27674 16292
rect 27690 16348 27754 16352
rect 27690 16292 27694 16348
rect 27694 16292 27750 16348
rect 27750 16292 27754 16348
rect 27690 16288 27754 16292
rect 27770 16348 27834 16352
rect 27770 16292 27774 16348
rect 27774 16292 27830 16348
rect 27830 16292 27834 16348
rect 27770 16288 27834 16292
rect 27850 16348 27914 16352
rect 27850 16292 27854 16348
rect 27854 16292 27910 16348
rect 27910 16292 27914 16348
rect 27850 16288 27914 16292
rect 4666 15804 4730 15808
rect 4666 15748 4670 15804
rect 4670 15748 4726 15804
rect 4726 15748 4730 15804
rect 4666 15744 4730 15748
rect 4746 15804 4810 15808
rect 4746 15748 4750 15804
rect 4750 15748 4806 15804
rect 4806 15748 4810 15804
rect 4746 15744 4810 15748
rect 4826 15804 4890 15808
rect 4826 15748 4830 15804
rect 4830 15748 4886 15804
rect 4886 15748 4890 15804
rect 4826 15744 4890 15748
rect 4906 15804 4970 15808
rect 4906 15748 4910 15804
rect 4910 15748 4966 15804
rect 4966 15748 4970 15804
rect 4906 15744 4970 15748
rect 12094 15804 12158 15808
rect 12094 15748 12098 15804
rect 12098 15748 12154 15804
rect 12154 15748 12158 15804
rect 12094 15744 12158 15748
rect 12174 15804 12238 15808
rect 12174 15748 12178 15804
rect 12178 15748 12234 15804
rect 12234 15748 12238 15804
rect 12174 15744 12238 15748
rect 12254 15804 12318 15808
rect 12254 15748 12258 15804
rect 12258 15748 12314 15804
rect 12314 15748 12318 15804
rect 12254 15744 12318 15748
rect 12334 15804 12398 15808
rect 12334 15748 12338 15804
rect 12338 15748 12394 15804
rect 12394 15748 12398 15804
rect 12334 15744 12398 15748
rect 19522 15804 19586 15808
rect 19522 15748 19526 15804
rect 19526 15748 19582 15804
rect 19582 15748 19586 15804
rect 19522 15744 19586 15748
rect 19602 15804 19666 15808
rect 19602 15748 19606 15804
rect 19606 15748 19662 15804
rect 19662 15748 19666 15804
rect 19602 15744 19666 15748
rect 19682 15804 19746 15808
rect 19682 15748 19686 15804
rect 19686 15748 19742 15804
rect 19742 15748 19746 15804
rect 19682 15744 19746 15748
rect 19762 15804 19826 15808
rect 19762 15748 19766 15804
rect 19766 15748 19822 15804
rect 19822 15748 19826 15804
rect 19762 15744 19826 15748
rect 26950 15804 27014 15808
rect 26950 15748 26954 15804
rect 26954 15748 27010 15804
rect 27010 15748 27014 15804
rect 26950 15744 27014 15748
rect 27030 15804 27094 15808
rect 27030 15748 27034 15804
rect 27034 15748 27090 15804
rect 27090 15748 27094 15804
rect 27030 15744 27094 15748
rect 27110 15804 27174 15808
rect 27110 15748 27114 15804
rect 27114 15748 27170 15804
rect 27170 15748 27174 15804
rect 27110 15744 27174 15748
rect 27190 15804 27254 15808
rect 27190 15748 27194 15804
rect 27194 15748 27250 15804
rect 27250 15748 27254 15804
rect 27190 15744 27254 15748
rect 5326 15260 5390 15264
rect 5326 15204 5330 15260
rect 5330 15204 5386 15260
rect 5386 15204 5390 15260
rect 5326 15200 5390 15204
rect 5406 15260 5470 15264
rect 5406 15204 5410 15260
rect 5410 15204 5466 15260
rect 5466 15204 5470 15260
rect 5406 15200 5470 15204
rect 5486 15260 5550 15264
rect 5486 15204 5490 15260
rect 5490 15204 5546 15260
rect 5546 15204 5550 15260
rect 5486 15200 5550 15204
rect 5566 15260 5630 15264
rect 5566 15204 5570 15260
rect 5570 15204 5626 15260
rect 5626 15204 5630 15260
rect 5566 15200 5630 15204
rect 12754 15260 12818 15264
rect 12754 15204 12758 15260
rect 12758 15204 12814 15260
rect 12814 15204 12818 15260
rect 12754 15200 12818 15204
rect 12834 15260 12898 15264
rect 12834 15204 12838 15260
rect 12838 15204 12894 15260
rect 12894 15204 12898 15260
rect 12834 15200 12898 15204
rect 12914 15260 12978 15264
rect 12914 15204 12918 15260
rect 12918 15204 12974 15260
rect 12974 15204 12978 15260
rect 12914 15200 12978 15204
rect 12994 15260 13058 15264
rect 12994 15204 12998 15260
rect 12998 15204 13054 15260
rect 13054 15204 13058 15260
rect 12994 15200 13058 15204
rect 20182 15260 20246 15264
rect 20182 15204 20186 15260
rect 20186 15204 20242 15260
rect 20242 15204 20246 15260
rect 20182 15200 20246 15204
rect 20262 15260 20326 15264
rect 20262 15204 20266 15260
rect 20266 15204 20322 15260
rect 20322 15204 20326 15260
rect 20262 15200 20326 15204
rect 20342 15260 20406 15264
rect 20342 15204 20346 15260
rect 20346 15204 20402 15260
rect 20402 15204 20406 15260
rect 20342 15200 20406 15204
rect 20422 15260 20486 15264
rect 20422 15204 20426 15260
rect 20426 15204 20482 15260
rect 20482 15204 20486 15260
rect 20422 15200 20486 15204
rect 27610 15260 27674 15264
rect 27610 15204 27614 15260
rect 27614 15204 27670 15260
rect 27670 15204 27674 15260
rect 27610 15200 27674 15204
rect 27690 15260 27754 15264
rect 27690 15204 27694 15260
rect 27694 15204 27750 15260
rect 27750 15204 27754 15260
rect 27690 15200 27754 15204
rect 27770 15260 27834 15264
rect 27770 15204 27774 15260
rect 27774 15204 27830 15260
rect 27830 15204 27834 15260
rect 27770 15200 27834 15204
rect 27850 15260 27914 15264
rect 27850 15204 27854 15260
rect 27854 15204 27910 15260
rect 27910 15204 27914 15260
rect 27850 15200 27914 15204
rect 4666 14716 4730 14720
rect 4666 14660 4670 14716
rect 4670 14660 4726 14716
rect 4726 14660 4730 14716
rect 4666 14656 4730 14660
rect 4746 14716 4810 14720
rect 4746 14660 4750 14716
rect 4750 14660 4806 14716
rect 4806 14660 4810 14716
rect 4746 14656 4810 14660
rect 4826 14716 4890 14720
rect 4826 14660 4830 14716
rect 4830 14660 4886 14716
rect 4886 14660 4890 14716
rect 4826 14656 4890 14660
rect 4906 14716 4970 14720
rect 4906 14660 4910 14716
rect 4910 14660 4966 14716
rect 4966 14660 4970 14716
rect 4906 14656 4970 14660
rect 12094 14716 12158 14720
rect 12094 14660 12098 14716
rect 12098 14660 12154 14716
rect 12154 14660 12158 14716
rect 12094 14656 12158 14660
rect 12174 14716 12238 14720
rect 12174 14660 12178 14716
rect 12178 14660 12234 14716
rect 12234 14660 12238 14716
rect 12174 14656 12238 14660
rect 12254 14716 12318 14720
rect 12254 14660 12258 14716
rect 12258 14660 12314 14716
rect 12314 14660 12318 14716
rect 12254 14656 12318 14660
rect 12334 14716 12398 14720
rect 12334 14660 12338 14716
rect 12338 14660 12394 14716
rect 12394 14660 12398 14716
rect 12334 14656 12398 14660
rect 19522 14716 19586 14720
rect 19522 14660 19526 14716
rect 19526 14660 19582 14716
rect 19582 14660 19586 14716
rect 19522 14656 19586 14660
rect 19602 14716 19666 14720
rect 19602 14660 19606 14716
rect 19606 14660 19662 14716
rect 19662 14660 19666 14716
rect 19602 14656 19666 14660
rect 19682 14716 19746 14720
rect 19682 14660 19686 14716
rect 19686 14660 19742 14716
rect 19742 14660 19746 14716
rect 19682 14656 19746 14660
rect 19762 14716 19826 14720
rect 19762 14660 19766 14716
rect 19766 14660 19822 14716
rect 19822 14660 19826 14716
rect 19762 14656 19826 14660
rect 26950 14716 27014 14720
rect 26950 14660 26954 14716
rect 26954 14660 27010 14716
rect 27010 14660 27014 14716
rect 26950 14656 27014 14660
rect 27030 14716 27094 14720
rect 27030 14660 27034 14716
rect 27034 14660 27090 14716
rect 27090 14660 27094 14716
rect 27030 14656 27094 14660
rect 27110 14716 27174 14720
rect 27110 14660 27114 14716
rect 27114 14660 27170 14716
rect 27170 14660 27174 14716
rect 27110 14656 27174 14660
rect 27190 14716 27254 14720
rect 27190 14660 27194 14716
rect 27194 14660 27250 14716
rect 27250 14660 27254 14716
rect 27190 14656 27254 14660
rect 5326 14172 5390 14176
rect 5326 14116 5330 14172
rect 5330 14116 5386 14172
rect 5386 14116 5390 14172
rect 5326 14112 5390 14116
rect 5406 14172 5470 14176
rect 5406 14116 5410 14172
rect 5410 14116 5466 14172
rect 5466 14116 5470 14172
rect 5406 14112 5470 14116
rect 5486 14172 5550 14176
rect 5486 14116 5490 14172
rect 5490 14116 5546 14172
rect 5546 14116 5550 14172
rect 5486 14112 5550 14116
rect 5566 14172 5630 14176
rect 5566 14116 5570 14172
rect 5570 14116 5626 14172
rect 5626 14116 5630 14172
rect 5566 14112 5630 14116
rect 12754 14172 12818 14176
rect 12754 14116 12758 14172
rect 12758 14116 12814 14172
rect 12814 14116 12818 14172
rect 12754 14112 12818 14116
rect 12834 14172 12898 14176
rect 12834 14116 12838 14172
rect 12838 14116 12894 14172
rect 12894 14116 12898 14172
rect 12834 14112 12898 14116
rect 12914 14172 12978 14176
rect 12914 14116 12918 14172
rect 12918 14116 12974 14172
rect 12974 14116 12978 14172
rect 12914 14112 12978 14116
rect 12994 14172 13058 14176
rect 12994 14116 12998 14172
rect 12998 14116 13054 14172
rect 13054 14116 13058 14172
rect 12994 14112 13058 14116
rect 20182 14172 20246 14176
rect 20182 14116 20186 14172
rect 20186 14116 20242 14172
rect 20242 14116 20246 14172
rect 20182 14112 20246 14116
rect 20262 14172 20326 14176
rect 20262 14116 20266 14172
rect 20266 14116 20322 14172
rect 20322 14116 20326 14172
rect 20262 14112 20326 14116
rect 20342 14172 20406 14176
rect 20342 14116 20346 14172
rect 20346 14116 20402 14172
rect 20402 14116 20406 14172
rect 20342 14112 20406 14116
rect 20422 14172 20486 14176
rect 20422 14116 20426 14172
rect 20426 14116 20482 14172
rect 20482 14116 20486 14172
rect 20422 14112 20486 14116
rect 27610 14172 27674 14176
rect 27610 14116 27614 14172
rect 27614 14116 27670 14172
rect 27670 14116 27674 14172
rect 27610 14112 27674 14116
rect 27690 14172 27754 14176
rect 27690 14116 27694 14172
rect 27694 14116 27750 14172
rect 27750 14116 27754 14172
rect 27690 14112 27754 14116
rect 27770 14172 27834 14176
rect 27770 14116 27774 14172
rect 27774 14116 27830 14172
rect 27830 14116 27834 14172
rect 27770 14112 27834 14116
rect 27850 14172 27914 14176
rect 27850 14116 27854 14172
rect 27854 14116 27910 14172
rect 27910 14116 27914 14172
rect 27850 14112 27914 14116
rect 4666 13628 4730 13632
rect 4666 13572 4670 13628
rect 4670 13572 4726 13628
rect 4726 13572 4730 13628
rect 4666 13568 4730 13572
rect 4746 13628 4810 13632
rect 4746 13572 4750 13628
rect 4750 13572 4806 13628
rect 4806 13572 4810 13628
rect 4746 13568 4810 13572
rect 4826 13628 4890 13632
rect 4826 13572 4830 13628
rect 4830 13572 4886 13628
rect 4886 13572 4890 13628
rect 4826 13568 4890 13572
rect 4906 13628 4970 13632
rect 4906 13572 4910 13628
rect 4910 13572 4966 13628
rect 4966 13572 4970 13628
rect 4906 13568 4970 13572
rect 12094 13628 12158 13632
rect 12094 13572 12098 13628
rect 12098 13572 12154 13628
rect 12154 13572 12158 13628
rect 12094 13568 12158 13572
rect 12174 13628 12238 13632
rect 12174 13572 12178 13628
rect 12178 13572 12234 13628
rect 12234 13572 12238 13628
rect 12174 13568 12238 13572
rect 12254 13628 12318 13632
rect 12254 13572 12258 13628
rect 12258 13572 12314 13628
rect 12314 13572 12318 13628
rect 12254 13568 12318 13572
rect 12334 13628 12398 13632
rect 12334 13572 12338 13628
rect 12338 13572 12394 13628
rect 12394 13572 12398 13628
rect 12334 13568 12398 13572
rect 19522 13628 19586 13632
rect 19522 13572 19526 13628
rect 19526 13572 19582 13628
rect 19582 13572 19586 13628
rect 19522 13568 19586 13572
rect 19602 13628 19666 13632
rect 19602 13572 19606 13628
rect 19606 13572 19662 13628
rect 19662 13572 19666 13628
rect 19602 13568 19666 13572
rect 19682 13628 19746 13632
rect 19682 13572 19686 13628
rect 19686 13572 19742 13628
rect 19742 13572 19746 13628
rect 19682 13568 19746 13572
rect 19762 13628 19826 13632
rect 19762 13572 19766 13628
rect 19766 13572 19822 13628
rect 19822 13572 19826 13628
rect 19762 13568 19826 13572
rect 26950 13628 27014 13632
rect 26950 13572 26954 13628
rect 26954 13572 27010 13628
rect 27010 13572 27014 13628
rect 26950 13568 27014 13572
rect 27030 13628 27094 13632
rect 27030 13572 27034 13628
rect 27034 13572 27090 13628
rect 27090 13572 27094 13628
rect 27030 13568 27094 13572
rect 27110 13628 27174 13632
rect 27110 13572 27114 13628
rect 27114 13572 27170 13628
rect 27170 13572 27174 13628
rect 27110 13568 27174 13572
rect 27190 13628 27254 13632
rect 27190 13572 27194 13628
rect 27194 13572 27250 13628
rect 27250 13572 27254 13628
rect 27190 13568 27254 13572
rect 5326 13084 5390 13088
rect 5326 13028 5330 13084
rect 5330 13028 5386 13084
rect 5386 13028 5390 13084
rect 5326 13024 5390 13028
rect 5406 13084 5470 13088
rect 5406 13028 5410 13084
rect 5410 13028 5466 13084
rect 5466 13028 5470 13084
rect 5406 13024 5470 13028
rect 5486 13084 5550 13088
rect 5486 13028 5490 13084
rect 5490 13028 5546 13084
rect 5546 13028 5550 13084
rect 5486 13024 5550 13028
rect 5566 13084 5630 13088
rect 5566 13028 5570 13084
rect 5570 13028 5626 13084
rect 5626 13028 5630 13084
rect 5566 13024 5630 13028
rect 12754 13084 12818 13088
rect 12754 13028 12758 13084
rect 12758 13028 12814 13084
rect 12814 13028 12818 13084
rect 12754 13024 12818 13028
rect 12834 13084 12898 13088
rect 12834 13028 12838 13084
rect 12838 13028 12894 13084
rect 12894 13028 12898 13084
rect 12834 13024 12898 13028
rect 12914 13084 12978 13088
rect 12914 13028 12918 13084
rect 12918 13028 12974 13084
rect 12974 13028 12978 13084
rect 12914 13024 12978 13028
rect 12994 13084 13058 13088
rect 12994 13028 12998 13084
rect 12998 13028 13054 13084
rect 13054 13028 13058 13084
rect 12994 13024 13058 13028
rect 20182 13084 20246 13088
rect 20182 13028 20186 13084
rect 20186 13028 20242 13084
rect 20242 13028 20246 13084
rect 20182 13024 20246 13028
rect 20262 13084 20326 13088
rect 20262 13028 20266 13084
rect 20266 13028 20322 13084
rect 20322 13028 20326 13084
rect 20262 13024 20326 13028
rect 20342 13084 20406 13088
rect 20342 13028 20346 13084
rect 20346 13028 20402 13084
rect 20402 13028 20406 13084
rect 20342 13024 20406 13028
rect 20422 13084 20486 13088
rect 20422 13028 20426 13084
rect 20426 13028 20482 13084
rect 20482 13028 20486 13084
rect 20422 13024 20486 13028
rect 27610 13084 27674 13088
rect 27610 13028 27614 13084
rect 27614 13028 27670 13084
rect 27670 13028 27674 13084
rect 27610 13024 27674 13028
rect 27690 13084 27754 13088
rect 27690 13028 27694 13084
rect 27694 13028 27750 13084
rect 27750 13028 27754 13084
rect 27690 13024 27754 13028
rect 27770 13084 27834 13088
rect 27770 13028 27774 13084
rect 27774 13028 27830 13084
rect 27830 13028 27834 13084
rect 27770 13024 27834 13028
rect 27850 13084 27914 13088
rect 27850 13028 27854 13084
rect 27854 13028 27910 13084
rect 27910 13028 27914 13084
rect 27850 13024 27914 13028
rect 4666 12540 4730 12544
rect 4666 12484 4670 12540
rect 4670 12484 4726 12540
rect 4726 12484 4730 12540
rect 4666 12480 4730 12484
rect 4746 12540 4810 12544
rect 4746 12484 4750 12540
rect 4750 12484 4806 12540
rect 4806 12484 4810 12540
rect 4746 12480 4810 12484
rect 4826 12540 4890 12544
rect 4826 12484 4830 12540
rect 4830 12484 4886 12540
rect 4886 12484 4890 12540
rect 4826 12480 4890 12484
rect 4906 12540 4970 12544
rect 4906 12484 4910 12540
rect 4910 12484 4966 12540
rect 4966 12484 4970 12540
rect 4906 12480 4970 12484
rect 12094 12540 12158 12544
rect 12094 12484 12098 12540
rect 12098 12484 12154 12540
rect 12154 12484 12158 12540
rect 12094 12480 12158 12484
rect 12174 12540 12238 12544
rect 12174 12484 12178 12540
rect 12178 12484 12234 12540
rect 12234 12484 12238 12540
rect 12174 12480 12238 12484
rect 12254 12540 12318 12544
rect 12254 12484 12258 12540
rect 12258 12484 12314 12540
rect 12314 12484 12318 12540
rect 12254 12480 12318 12484
rect 12334 12540 12398 12544
rect 12334 12484 12338 12540
rect 12338 12484 12394 12540
rect 12394 12484 12398 12540
rect 12334 12480 12398 12484
rect 19522 12540 19586 12544
rect 19522 12484 19526 12540
rect 19526 12484 19582 12540
rect 19582 12484 19586 12540
rect 19522 12480 19586 12484
rect 19602 12540 19666 12544
rect 19602 12484 19606 12540
rect 19606 12484 19662 12540
rect 19662 12484 19666 12540
rect 19602 12480 19666 12484
rect 19682 12540 19746 12544
rect 19682 12484 19686 12540
rect 19686 12484 19742 12540
rect 19742 12484 19746 12540
rect 19682 12480 19746 12484
rect 19762 12540 19826 12544
rect 19762 12484 19766 12540
rect 19766 12484 19822 12540
rect 19822 12484 19826 12540
rect 19762 12480 19826 12484
rect 26950 12540 27014 12544
rect 26950 12484 26954 12540
rect 26954 12484 27010 12540
rect 27010 12484 27014 12540
rect 26950 12480 27014 12484
rect 27030 12540 27094 12544
rect 27030 12484 27034 12540
rect 27034 12484 27090 12540
rect 27090 12484 27094 12540
rect 27030 12480 27094 12484
rect 27110 12540 27174 12544
rect 27110 12484 27114 12540
rect 27114 12484 27170 12540
rect 27170 12484 27174 12540
rect 27110 12480 27174 12484
rect 27190 12540 27254 12544
rect 27190 12484 27194 12540
rect 27194 12484 27250 12540
rect 27250 12484 27254 12540
rect 27190 12480 27254 12484
rect 5326 11996 5390 12000
rect 5326 11940 5330 11996
rect 5330 11940 5386 11996
rect 5386 11940 5390 11996
rect 5326 11936 5390 11940
rect 5406 11996 5470 12000
rect 5406 11940 5410 11996
rect 5410 11940 5466 11996
rect 5466 11940 5470 11996
rect 5406 11936 5470 11940
rect 5486 11996 5550 12000
rect 5486 11940 5490 11996
rect 5490 11940 5546 11996
rect 5546 11940 5550 11996
rect 5486 11936 5550 11940
rect 5566 11996 5630 12000
rect 5566 11940 5570 11996
rect 5570 11940 5626 11996
rect 5626 11940 5630 11996
rect 5566 11936 5630 11940
rect 12754 11996 12818 12000
rect 12754 11940 12758 11996
rect 12758 11940 12814 11996
rect 12814 11940 12818 11996
rect 12754 11936 12818 11940
rect 12834 11996 12898 12000
rect 12834 11940 12838 11996
rect 12838 11940 12894 11996
rect 12894 11940 12898 11996
rect 12834 11936 12898 11940
rect 12914 11996 12978 12000
rect 12914 11940 12918 11996
rect 12918 11940 12974 11996
rect 12974 11940 12978 11996
rect 12914 11936 12978 11940
rect 12994 11996 13058 12000
rect 12994 11940 12998 11996
rect 12998 11940 13054 11996
rect 13054 11940 13058 11996
rect 12994 11936 13058 11940
rect 20182 11996 20246 12000
rect 20182 11940 20186 11996
rect 20186 11940 20242 11996
rect 20242 11940 20246 11996
rect 20182 11936 20246 11940
rect 20262 11996 20326 12000
rect 20262 11940 20266 11996
rect 20266 11940 20322 11996
rect 20322 11940 20326 11996
rect 20262 11936 20326 11940
rect 20342 11996 20406 12000
rect 20342 11940 20346 11996
rect 20346 11940 20402 11996
rect 20402 11940 20406 11996
rect 20342 11936 20406 11940
rect 20422 11996 20486 12000
rect 20422 11940 20426 11996
rect 20426 11940 20482 11996
rect 20482 11940 20486 11996
rect 20422 11936 20486 11940
rect 27610 11996 27674 12000
rect 27610 11940 27614 11996
rect 27614 11940 27670 11996
rect 27670 11940 27674 11996
rect 27610 11936 27674 11940
rect 27690 11996 27754 12000
rect 27690 11940 27694 11996
rect 27694 11940 27750 11996
rect 27750 11940 27754 11996
rect 27690 11936 27754 11940
rect 27770 11996 27834 12000
rect 27770 11940 27774 11996
rect 27774 11940 27830 11996
rect 27830 11940 27834 11996
rect 27770 11936 27834 11940
rect 27850 11996 27914 12000
rect 27850 11940 27854 11996
rect 27854 11940 27910 11996
rect 27910 11940 27914 11996
rect 27850 11936 27914 11940
rect 4666 11452 4730 11456
rect 4666 11396 4670 11452
rect 4670 11396 4726 11452
rect 4726 11396 4730 11452
rect 4666 11392 4730 11396
rect 4746 11452 4810 11456
rect 4746 11396 4750 11452
rect 4750 11396 4806 11452
rect 4806 11396 4810 11452
rect 4746 11392 4810 11396
rect 4826 11452 4890 11456
rect 4826 11396 4830 11452
rect 4830 11396 4886 11452
rect 4886 11396 4890 11452
rect 4826 11392 4890 11396
rect 4906 11452 4970 11456
rect 4906 11396 4910 11452
rect 4910 11396 4966 11452
rect 4966 11396 4970 11452
rect 4906 11392 4970 11396
rect 12094 11452 12158 11456
rect 12094 11396 12098 11452
rect 12098 11396 12154 11452
rect 12154 11396 12158 11452
rect 12094 11392 12158 11396
rect 12174 11452 12238 11456
rect 12174 11396 12178 11452
rect 12178 11396 12234 11452
rect 12234 11396 12238 11452
rect 12174 11392 12238 11396
rect 12254 11452 12318 11456
rect 12254 11396 12258 11452
rect 12258 11396 12314 11452
rect 12314 11396 12318 11452
rect 12254 11392 12318 11396
rect 12334 11452 12398 11456
rect 12334 11396 12338 11452
rect 12338 11396 12394 11452
rect 12394 11396 12398 11452
rect 12334 11392 12398 11396
rect 19522 11452 19586 11456
rect 19522 11396 19526 11452
rect 19526 11396 19582 11452
rect 19582 11396 19586 11452
rect 19522 11392 19586 11396
rect 19602 11452 19666 11456
rect 19602 11396 19606 11452
rect 19606 11396 19662 11452
rect 19662 11396 19666 11452
rect 19602 11392 19666 11396
rect 19682 11452 19746 11456
rect 19682 11396 19686 11452
rect 19686 11396 19742 11452
rect 19742 11396 19746 11452
rect 19682 11392 19746 11396
rect 19762 11452 19826 11456
rect 19762 11396 19766 11452
rect 19766 11396 19822 11452
rect 19822 11396 19826 11452
rect 19762 11392 19826 11396
rect 26950 11452 27014 11456
rect 26950 11396 26954 11452
rect 26954 11396 27010 11452
rect 27010 11396 27014 11452
rect 26950 11392 27014 11396
rect 27030 11452 27094 11456
rect 27030 11396 27034 11452
rect 27034 11396 27090 11452
rect 27090 11396 27094 11452
rect 27030 11392 27094 11396
rect 27110 11452 27174 11456
rect 27110 11396 27114 11452
rect 27114 11396 27170 11452
rect 27170 11396 27174 11452
rect 27110 11392 27174 11396
rect 27190 11452 27254 11456
rect 27190 11396 27194 11452
rect 27194 11396 27250 11452
rect 27250 11396 27254 11452
rect 27190 11392 27254 11396
rect 5326 10908 5390 10912
rect 5326 10852 5330 10908
rect 5330 10852 5386 10908
rect 5386 10852 5390 10908
rect 5326 10848 5390 10852
rect 5406 10908 5470 10912
rect 5406 10852 5410 10908
rect 5410 10852 5466 10908
rect 5466 10852 5470 10908
rect 5406 10848 5470 10852
rect 5486 10908 5550 10912
rect 5486 10852 5490 10908
rect 5490 10852 5546 10908
rect 5546 10852 5550 10908
rect 5486 10848 5550 10852
rect 5566 10908 5630 10912
rect 5566 10852 5570 10908
rect 5570 10852 5626 10908
rect 5626 10852 5630 10908
rect 5566 10848 5630 10852
rect 12754 10908 12818 10912
rect 12754 10852 12758 10908
rect 12758 10852 12814 10908
rect 12814 10852 12818 10908
rect 12754 10848 12818 10852
rect 12834 10908 12898 10912
rect 12834 10852 12838 10908
rect 12838 10852 12894 10908
rect 12894 10852 12898 10908
rect 12834 10848 12898 10852
rect 12914 10908 12978 10912
rect 12914 10852 12918 10908
rect 12918 10852 12974 10908
rect 12974 10852 12978 10908
rect 12914 10848 12978 10852
rect 12994 10908 13058 10912
rect 12994 10852 12998 10908
rect 12998 10852 13054 10908
rect 13054 10852 13058 10908
rect 12994 10848 13058 10852
rect 20182 10908 20246 10912
rect 20182 10852 20186 10908
rect 20186 10852 20242 10908
rect 20242 10852 20246 10908
rect 20182 10848 20246 10852
rect 20262 10908 20326 10912
rect 20262 10852 20266 10908
rect 20266 10852 20322 10908
rect 20322 10852 20326 10908
rect 20262 10848 20326 10852
rect 20342 10908 20406 10912
rect 20342 10852 20346 10908
rect 20346 10852 20402 10908
rect 20402 10852 20406 10908
rect 20342 10848 20406 10852
rect 20422 10908 20486 10912
rect 20422 10852 20426 10908
rect 20426 10852 20482 10908
rect 20482 10852 20486 10908
rect 20422 10848 20486 10852
rect 27610 10908 27674 10912
rect 27610 10852 27614 10908
rect 27614 10852 27670 10908
rect 27670 10852 27674 10908
rect 27610 10848 27674 10852
rect 27690 10908 27754 10912
rect 27690 10852 27694 10908
rect 27694 10852 27750 10908
rect 27750 10852 27754 10908
rect 27690 10848 27754 10852
rect 27770 10908 27834 10912
rect 27770 10852 27774 10908
rect 27774 10852 27830 10908
rect 27830 10852 27834 10908
rect 27770 10848 27834 10852
rect 27850 10908 27914 10912
rect 27850 10852 27854 10908
rect 27854 10852 27910 10908
rect 27910 10852 27914 10908
rect 27850 10848 27914 10852
rect 4666 10364 4730 10368
rect 4666 10308 4670 10364
rect 4670 10308 4726 10364
rect 4726 10308 4730 10364
rect 4666 10304 4730 10308
rect 4746 10364 4810 10368
rect 4746 10308 4750 10364
rect 4750 10308 4806 10364
rect 4806 10308 4810 10364
rect 4746 10304 4810 10308
rect 4826 10364 4890 10368
rect 4826 10308 4830 10364
rect 4830 10308 4886 10364
rect 4886 10308 4890 10364
rect 4826 10304 4890 10308
rect 4906 10364 4970 10368
rect 4906 10308 4910 10364
rect 4910 10308 4966 10364
rect 4966 10308 4970 10364
rect 4906 10304 4970 10308
rect 12094 10364 12158 10368
rect 12094 10308 12098 10364
rect 12098 10308 12154 10364
rect 12154 10308 12158 10364
rect 12094 10304 12158 10308
rect 12174 10364 12238 10368
rect 12174 10308 12178 10364
rect 12178 10308 12234 10364
rect 12234 10308 12238 10364
rect 12174 10304 12238 10308
rect 12254 10364 12318 10368
rect 12254 10308 12258 10364
rect 12258 10308 12314 10364
rect 12314 10308 12318 10364
rect 12254 10304 12318 10308
rect 12334 10364 12398 10368
rect 12334 10308 12338 10364
rect 12338 10308 12394 10364
rect 12394 10308 12398 10364
rect 12334 10304 12398 10308
rect 19522 10364 19586 10368
rect 19522 10308 19526 10364
rect 19526 10308 19582 10364
rect 19582 10308 19586 10364
rect 19522 10304 19586 10308
rect 19602 10364 19666 10368
rect 19602 10308 19606 10364
rect 19606 10308 19662 10364
rect 19662 10308 19666 10364
rect 19602 10304 19666 10308
rect 19682 10364 19746 10368
rect 19682 10308 19686 10364
rect 19686 10308 19742 10364
rect 19742 10308 19746 10364
rect 19682 10304 19746 10308
rect 19762 10364 19826 10368
rect 19762 10308 19766 10364
rect 19766 10308 19822 10364
rect 19822 10308 19826 10364
rect 19762 10304 19826 10308
rect 26950 10364 27014 10368
rect 26950 10308 26954 10364
rect 26954 10308 27010 10364
rect 27010 10308 27014 10364
rect 26950 10304 27014 10308
rect 27030 10364 27094 10368
rect 27030 10308 27034 10364
rect 27034 10308 27090 10364
rect 27090 10308 27094 10364
rect 27030 10304 27094 10308
rect 27110 10364 27174 10368
rect 27110 10308 27114 10364
rect 27114 10308 27170 10364
rect 27170 10308 27174 10364
rect 27110 10304 27174 10308
rect 27190 10364 27254 10368
rect 27190 10308 27194 10364
rect 27194 10308 27250 10364
rect 27250 10308 27254 10364
rect 27190 10304 27254 10308
rect 5326 9820 5390 9824
rect 5326 9764 5330 9820
rect 5330 9764 5386 9820
rect 5386 9764 5390 9820
rect 5326 9760 5390 9764
rect 5406 9820 5470 9824
rect 5406 9764 5410 9820
rect 5410 9764 5466 9820
rect 5466 9764 5470 9820
rect 5406 9760 5470 9764
rect 5486 9820 5550 9824
rect 5486 9764 5490 9820
rect 5490 9764 5546 9820
rect 5546 9764 5550 9820
rect 5486 9760 5550 9764
rect 5566 9820 5630 9824
rect 5566 9764 5570 9820
rect 5570 9764 5626 9820
rect 5626 9764 5630 9820
rect 5566 9760 5630 9764
rect 12754 9820 12818 9824
rect 12754 9764 12758 9820
rect 12758 9764 12814 9820
rect 12814 9764 12818 9820
rect 12754 9760 12818 9764
rect 12834 9820 12898 9824
rect 12834 9764 12838 9820
rect 12838 9764 12894 9820
rect 12894 9764 12898 9820
rect 12834 9760 12898 9764
rect 12914 9820 12978 9824
rect 12914 9764 12918 9820
rect 12918 9764 12974 9820
rect 12974 9764 12978 9820
rect 12914 9760 12978 9764
rect 12994 9820 13058 9824
rect 12994 9764 12998 9820
rect 12998 9764 13054 9820
rect 13054 9764 13058 9820
rect 12994 9760 13058 9764
rect 20182 9820 20246 9824
rect 20182 9764 20186 9820
rect 20186 9764 20242 9820
rect 20242 9764 20246 9820
rect 20182 9760 20246 9764
rect 20262 9820 20326 9824
rect 20262 9764 20266 9820
rect 20266 9764 20322 9820
rect 20322 9764 20326 9820
rect 20262 9760 20326 9764
rect 20342 9820 20406 9824
rect 20342 9764 20346 9820
rect 20346 9764 20402 9820
rect 20402 9764 20406 9820
rect 20342 9760 20406 9764
rect 20422 9820 20486 9824
rect 20422 9764 20426 9820
rect 20426 9764 20482 9820
rect 20482 9764 20486 9820
rect 20422 9760 20486 9764
rect 27610 9820 27674 9824
rect 27610 9764 27614 9820
rect 27614 9764 27670 9820
rect 27670 9764 27674 9820
rect 27610 9760 27674 9764
rect 27690 9820 27754 9824
rect 27690 9764 27694 9820
rect 27694 9764 27750 9820
rect 27750 9764 27754 9820
rect 27690 9760 27754 9764
rect 27770 9820 27834 9824
rect 27770 9764 27774 9820
rect 27774 9764 27830 9820
rect 27830 9764 27834 9820
rect 27770 9760 27834 9764
rect 27850 9820 27914 9824
rect 27850 9764 27854 9820
rect 27854 9764 27910 9820
rect 27910 9764 27914 9820
rect 27850 9760 27914 9764
rect 4666 9276 4730 9280
rect 4666 9220 4670 9276
rect 4670 9220 4726 9276
rect 4726 9220 4730 9276
rect 4666 9216 4730 9220
rect 4746 9276 4810 9280
rect 4746 9220 4750 9276
rect 4750 9220 4806 9276
rect 4806 9220 4810 9276
rect 4746 9216 4810 9220
rect 4826 9276 4890 9280
rect 4826 9220 4830 9276
rect 4830 9220 4886 9276
rect 4886 9220 4890 9276
rect 4826 9216 4890 9220
rect 4906 9276 4970 9280
rect 4906 9220 4910 9276
rect 4910 9220 4966 9276
rect 4966 9220 4970 9276
rect 4906 9216 4970 9220
rect 12094 9276 12158 9280
rect 12094 9220 12098 9276
rect 12098 9220 12154 9276
rect 12154 9220 12158 9276
rect 12094 9216 12158 9220
rect 12174 9276 12238 9280
rect 12174 9220 12178 9276
rect 12178 9220 12234 9276
rect 12234 9220 12238 9276
rect 12174 9216 12238 9220
rect 12254 9276 12318 9280
rect 12254 9220 12258 9276
rect 12258 9220 12314 9276
rect 12314 9220 12318 9276
rect 12254 9216 12318 9220
rect 12334 9276 12398 9280
rect 12334 9220 12338 9276
rect 12338 9220 12394 9276
rect 12394 9220 12398 9276
rect 12334 9216 12398 9220
rect 19522 9276 19586 9280
rect 19522 9220 19526 9276
rect 19526 9220 19582 9276
rect 19582 9220 19586 9276
rect 19522 9216 19586 9220
rect 19602 9276 19666 9280
rect 19602 9220 19606 9276
rect 19606 9220 19662 9276
rect 19662 9220 19666 9276
rect 19602 9216 19666 9220
rect 19682 9276 19746 9280
rect 19682 9220 19686 9276
rect 19686 9220 19742 9276
rect 19742 9220 19746 9276
rect 19682 9216 19746 9220
rect 19762 9276 19826 9280
rect 19762 9220 19766 9276
rect 19766 9220 19822 9276
rect 19822 9220 19826 9276
rect 19762 9216 19826 9220
rect 26950 9276 27014 9280
rect 26950 9220 26954 9276
rect 26954 9220 27010 9276
rect 27010 9220 27014 9276
rect 26950 9216 27014 9220
rect 27030 9276 27094 9280
rect 27030 9220 27034 9276
rect 27034 9220 27090 9276
rect 27090 9220 27094 9276
rect 27030 9216 27094 9220
rect 27110 9276 27174 9280
rect 27110 9220 27114 9276
rect 27114 9220 27170 9276
rect 27170 9220 27174 9276
rect 27110 9216 27174 9220
rect 27190 9276 27254 9280
rect 27190 9220 27194 9276
rect 27194 9220 27250 9276
rect 27250 9220 27254 9276
rect 27190 9216 27254 9220
rect 5326 8732 5390 8736
rect 5326 8676 5330 8732
rect 5330 8676 5386 8732
rect 5386 8676 5390 8732
rect 5326 8672 5390 8676
rect 5406 8732 5470 8736
rect 5406 8676 5410 8732
rect 5410 8676 5466 8732
rect 5466 8676 5470 8732
rect 5406 8672 5470 8676
rect 5486 8732 5550 8736
rect 5486 8676 5490 8732
rect 5490 8676 5546 8732
rect 5546 8676 5550 8732
rect 5486 8672 5550 8676
rect 5566 8732 5630 8736
rect 5566 8676 5570 8732
rect 5570 8676 5626 8732
rect 5626 8676 5630 8732
rect 5566 8672 5630 8676
rect 12754 8732 12818 8736
rect 12754 8676 12758 8732
rect 12758 8676 12814 8732
rect 12814 8676 12818 8732
rect 12754 8672 12818 8676
rect 12834 8732 12898 8736
rect 12834 8676 12838 8732
rect 12838 8676 12894 8732
rect 12894 8676 12898 8732
rect 12834 8672 12898 8676
rect 12914 8732 12978 8736
rect 12914 8676 12918 8732
rect 12918 8676 12974 8732
rect 12974 8676 12978 8732
rect 12914 8672 12978 8676
rect 12994 8732 13058 8736
rect 12994 8676 12998 8732
rect 12998 8676 13054 8732
rect 13054 8676 13058 8732
rect 12994 8672 13058 8676
rect 20182 8732 20246 8736
rect 20182 8676 20186 8732
rect 20186 8676 20242 8732
rect 20242 8676 20246 8732
rect 20182 8672 20246 8676
rect 20262 8732 20326 8736
rect 20262 8676 20266 8732
rect 20266 8676 20322 8732
rect 20322 8676 20326 8732
rect 20262 8672 20326 8676
rect 20342 8732 20406 8736
rect 20342 8676 20346 8732
rect 20346 8676 20402 8732
rect 20402 8676 20406 8732
rect 20342 8672 20406 8676
rect 20422 8732 20486 8736
rect 20422 8676 20426 8732
rect 20426 8676 20482 8732
rect 20482 8676 20486 8732
rect 20422 8672 20486 8676
rect 27610 8732 27674 8736
rect 27610 8676 27614 8732
rect 27614 8676 27670 8732
rect 27670 8676 27674 8732
rect 27610 8672 27674 8676
rect 27690 8732 27754 8736
rect 27690 8676 27694 8732
rect 27694 8676 27750 8732
rect 27750 8676 27754 8732
rect 27690 8672 27754 8676
rect 27770 8732 27834 8736
rect 27770 8676 27774 8732
rect 27774 8676 27830 8732
rect 27830 8676 27834 8732
rect 27770 8672 27834 8676
rect 27850 8732 27914 8736
rect 27850 8676 27854 8732
rect 27854 8676 27910 8732
rect 27910 8676 27914 8732
rect 27850 8672 27914 8676
rect 4666 8188 4730 8192
rect 4666 8132 4670 8188
rect 4670 8132 4726 8188
rect 4726 8132 4730 8188
rect 4666 8128 4730 8132
rect 4746 8188 4810 8192
rect 4746 8132 4750 8188
rect 4750 8132 4806 8188
rect 4806 8132 4810 8188
rect 4746 8128 4810 8132
rect 4826 8188 4890 8192
rect 4826 8132 4830 8188
rect 4830 8132 4886 8188
rect 4886 8132 4890 8188
rect 4826 8128 4890 8132
rect 4906 8188 4970 8192
rect 4906 8132 4910 8188
rect 4910 8132 4966 8188
rect 4966 8132 4970 8188
rect 4906 8128 4970 8132
rect 12094 8188 12158 8192
rect 12094 8132 12098 8188
rect 12098 8132 12154 8188
rect 12154 8132 12158 8188
rect 12094 8128 12158 8132
rect 12174 8188 12238 8192
rect 12174 8132 12178 8188
rect 12178 8132 12234 8188
rect 12234 8132 12238 8188
rect 12174 8128 12238 8132
rect 12254 8188 12318 8192
rect 12254 8132 12258 8188
rect 12258 8132 12314 8188
rect 12314 8132 12318 8188
rect 12254 8128 12318 8132
rect 12334 8188 12398 8192
rect 12334 8132 12338 8188
rect 12338 8132 12394 8188
rect 12394 8132 12398 8188
rect 12334 8128 12398 8132
rect 19522 8188 19586 8192
rect 19522 8132 19526 8188
rect 19526 8132 19582 8188
rect 19582 8132 19586 8188
rect 19522 8128 19586 8132
rect 19602 8188 19666 8192
rect 19602 8132 19606 8188
rect 19606 8132 19662 8188
rect 19662 8132 19666 8188
rect 19602 8128 19666 8132
rect 19682 8188 19746 8192
rect 19682 8132 19686 8188
rect 19686 8132 19742 8188
rect 19742 8132 19746 8188
rect 19682 8128 19746 8132
rect 19762 8188 19826 8192
rect 19762 8132 19766 8188
rect 19766 8132 19822 8188
rect 19822 8132 19826 8188
rect 19762 8128 19826 8132
rect 26950 8188 27014 8192
rect 26950 8132 26954 8188
rect 26954 8132 27010 8188
rect 27010 8132 27014 8188
rect 26950 8128 27014 8132
rect 27030 8188 27094 8192
rect 27030 8132 27034 8188
rect 27034 8132 27090 8188
rect 27090 8132 27094 8188
rect 27030 8128 27094 8132
rect 27110 8188 27174 8192
rect 27110 8132 27114 8188
rect 27114 8132 27170 8188
rect 27170 8132 27174 8188
rect 27110 8128 27174 8132
rect 27190 8188 27254 8192
rect 27190 8132 27194 8188
rect 27194 8132 27250 8188
rect 27250 8132 27254 8188
rect 27190 8128 27254 8132
rect 5326 7644 5390 7648
rect 5326 7588 5330 7644
rect 5330 7588 5386 7644
rect 5386 7588 5390 7644
rect 5326 7584 5390 7588
rect 5406 7644 5470 7648
rect 5406 7588 5410 7644
rect 5410 7588 5466 7644
rect 5466 7588 5470 7644
rect 5406 7584 5470 7588
rect 5486 7644 5550 7648
rect 5486 7588 5490 7644
rect 5490 7588 5546 7644
rect 5546 7588 5550 7644
rect 5486 7584 5550 7588
rect 5566 7644 5630 7648
rect 5566 7588 5570 7644
rect 5570 7588 5626 7644
rect 5626 7588 5630 7644
rect 5566 7584 5630 7588
rect 12754 7644 12818 7648
rect 12754 7588 12758 7644
rect 12758 7588 12814 7644
rect 12814 7588 12818 7644
rect 12754 7584 12818 7588
rect 12834 7644 12898 7648
rect 12834 7588 12838 7644
rect 12838 7588 12894 7644
rect 12894 7588 12898 7644
rect 12834 7584 12898 7588
rect 12914 7644 12978 7648
rect 12914 7588 12918 7644
rect 12918 7588 12974 7644
rect 12974 7588 12978 7644
rect 12914 7584 12978 7588
rect 12994 7644 13058 7648
rect 12994 7588 12998 7644
rect 12998 7588 13054 7644
rect 13054 7588 13058 7644
rect 12994 7584 13058 7588
rect 20182 7644 20246 7648
rect 20182 7588 20186 7644
rect 20186 7588 20242 7644
rect 20242 7588 20246 7644
rect 20182 7584 20246 7588
rect 20262 7644 20326 7648
rect 20262 7588 20266 7644
rect 20266 7588 20322 7644
rect 20322 7588 20326 7644
rect 20262 7584 20326 7588
rect 20342 7644 20406 7648
rect 20342 7588 20346 7644
rect 20346 7588 20402 7644
rect 20402 7588 20406 7644
rect 20342 7584 20406 7588
rect 20422 7644 20486 7648
rect 20422 7588 20426 7644
rect 20426 7588 20482 7644
rect 20482 7588 20486 7644
rect 20422 7584 20486 7588
rect 27610 7644 27674 7648
rect 27610 7588 27614 7644
rect 27614 7588 27670 7644
rect 27670 7588 27674 7644
rect 27610 7584 27674 7588
rect 27690 7644 27754 7648
rect 27690 7588 27694 7644
rect 27694 7588 27750 7644
rect 27750 7588 27754 7644
rect 27690 7584 27754 7588
rect 27770 7644 27834 7648
rect 27770 7588 27774 7644
rect 27774 7588 27830 7644
rect 27830 7588 27834 7644
rect 27770 7584 27834 7588
rect 27850 7644 27914 7648
rect 27850 7588 27854 7644
rect 27854 7588 27910 7644
rect 27910 7588 27914 7644
rect 27850 7584 27914 7588
rect 4666 7100 4730 7104
rect 4666 7044 4670 7100
rect 4670 7044 4726 7100
rect 4726 7044 4730 7100
rect 4666 7040 4730 7044
rect 4746 7100 4810 7104
rect 4746 7044 4750 7100
rect 4750 7044 4806 7100
rect 4806 7044 4810 7100
rect 4746 7040 4810 7044
rect 4826 7100 4890 7104
rect 4826 7044 4830 7100
rect 4830 7044 4886 7100
rect 4886 7044 4890 7100
rect 4826 7040 4890 7044
rect 4906 7100 4970 7104
rect 4906 7044 4910 7100
rect 4910 7044 4966 7100
rect 4966 7044 4970 7100
rect 4906 7040 4970 7044
rect 12094 7100 12158 7104
rect 12094 7044 12098 7100
rect 12098 7044 12154 7100
rect 12154 7044 12158 7100
rect 12094 7040 12158 7044
rect 12174 7100 12238 7104
rect 12174 7044 12178 7100
rect 12178 7044 12234 7100
rect 12234 7044 12238 7100
rect 12174 7040 12238 7044
rect 12254 7100 12318 7104
rect 12254 7044 12258 7100
rect 12258 7044 12314 7100
rect 12314 7044 12318 7100
rect 12254 7040 12318 7044
rect 12334 7100 12398 7104
rect 12334 7044 12338 7100
rect 12338 7044 12394 7100
rect 12394 7044 12398 7100
rect 12334 7040 12398 7044
rect 19522 7100 19586 7104
rect 19522 7044 19526 7100
rect 19526 7044 19582 7100
rect 19582 7044 19586 7100
rect 19522 7040 19586 7044
rect 19602 7100 19666 7104
rect 19602 7044 19606 7100
rect 19606 7044 19662 7100
rect 19662 7044 19666 7100
rect 19602 7040 19666 7044
rect 19682 7100 19746 7104
rect 19682 7044 19686 7100
rect 19686 7044 19742 7100
rect 19742 7044 19746 7100
rect 19682 7040 19746 7044
rect 19762 7100 19826 7104
rect 19762 7044 19766 7100
rect 19766 7044 19822 7100
rect 19822 7044 19826 7100
rect 19762 7040 19826 7044
rect 26950 7100 27014 7104
rect 26950 7044 26954 7100
rect 26954 7044 27010 7100
rect 27010 7044 27014 7100
rect 26950 7040 27014 7044
rect 27030 7100 27094 7104
rect 27030 7044 27034 7100
rect 27034 7044 27090 7100
rect 27090 7044 27094 7100
rect 27030 7040 27094 7044
rect 27110 7100 27174 7104
rect 27110 7044 27114 7100
rect 27114 7044 27170 7100
rect 27170 7044 27174 7100
rect 27110 7040 27174 7044
rect 27190 7100 27254 7104
rect 27190 7044 27194 7100
rect 27194 7044 27250 7100
rect 27250 7044 27254 7100
rect 27190 7040 27254 7044
rect 5326 6556 5390 6560
rect 5326 6500 5330 6556
rect 5330 6500 5386 6556
rect 5386 6500 5390 6556
rect 5326 6496 5390 6500
rect 5406 6556 5470 6560
rect 5406 6500 5410 6556
rect 5410 6500 5466 6556
rect 5466 6500 5470 6556
rect 5406 6496 5470 6500
rect 5486 6556 5550 6560
rect 5486 6500 5490 6556
rect 5490 6500 5546 6556
rect 5546 6500 5550 6556
rect 5486 6496 5550 6500
rect 5566 6556 5630 6560
rect 5566 6500 5570 6556
rect 5570 6500 5626 6556
rect 5626 6500 5630 6556
rect 5566 6496 5630 6500
rect 12754 6556 12818 6560
rect 12754 6500 12758 6556
rect 12758 6500 12814 6556
rect 12814 6500 12818 6556
rect 12754 6496 12818 6500
rect 12834 6556 12898 6560
rect 12834 6500 12838 6556
rect 12838 6500 12894 6556
rect 12894 6500 12898 6556
rect 12834 6496 12898 6500
rect 12914 6556 12978 6560
rect 12914 6500 12918 6556
rect 12918 6500 12974 6556
rect 12974 6500 12978 6556
rect 12914 6496 12978 6500
rect 12994 6556 13058 6560
rect 12994 6500 12998 6556
rect 12998 6500 13054 6556
rect 13054 6500 13058 6556
rect 12994 6496 13058 6500
rect 20182 6556 20246 6560
rect 20182 6500 20186 6556
rect 20186 6500 20242 6556
rect 20242 6500 20246 6556
rect 20182 6496 20246 6500
rect 20262 6556 20326 6560
rect 20262 6500 20266 6556
rect 20266 6500 20322 6556
rect 20322 6500 20326 6556
rect 20262 6496 20326 6500
rect 20342 6556 20406 6560
rect 20342 6500 20346 6556
rect 20346 6500 20402 6556
rect 20402 6500 20406 6556
rect 20342 6496 20406 6500
rect 20422 6556 20486 6560
rect 20422 6500 20426 6556
rect 20426 6500 20482 6556
rect 20482 6500 20486 6556
rect 20422 6496 20486 6500
rect 27610 6556 27674 6560
rect 27610 6500 27614 6556
rect 27614 6500 27670 6556
rect 27670 6500 27674 6556
rect 27610 6496 27674 6500
rect 27690 6556 27754 6560
rect 27690 6500 27694 6556
rect 27694 6500 27750 6556
rect 27750 6500 27754 6556
rect 27690 6496 27754 6500
rect 27770 6556 27834 6560
rect 27770 6500 27774 6556
rect 27774 6500 27830 6556
rect 27830 6500 27834 6556
rect 27770 6496 27834 6500
rect 27850 6556 27914 6560
rect 27850 6500 27854 6556
rect 27854 6500 27910 6556
rect 27910 6500 27914 6556
rect 27850 6496 27914 6500
rect 4666 6012 4730 6016
rect 4666 5956 4670 6012
rect 4670 5956 4726 6012
rect 4726 5956 4730 6012
rect 4666 5952 4730 5956
rect 4746 6012 4810 6016
rect 4746 5956 4750 6012
rect 4750 5956 4806 6012
rect 4806 5956 4810 6012
rect 4746 5952 4810 5956
rect 4826 6012 4890 6016
rect 4826 5956 4830 6012
rect 4830 5956 4886 6012
rect 4886 5956 4890 6012
rect 4826 5952 4890 5956
rect 4906 6012 4970 6016
rect 4906 5956 4910 6012
rect 4910 5956 4966 6012
rect 4966 5956 4970 6012
rect 4906 5952 4970 5956
rect 12094 6012 12158 6016
rect 12094 5956 12098 6012
rect 12098 5956 12154 6012
rect 12154 5956 12158 6012
rect 12094 5952 12158 5956
rect 12174 6012 12238 6016
rect 12174 5956 12178 6012
rect 12178 5956 12234 6012
rect 12234 5956 12238 6012
rect 12174 5952 12238 5956
rect 12254 6012 12318 6016
rect 12254 5956 12258 6012
rect 12258 5956 12314 6012
rect 12314 5956 12318 6012
rect 12254 5952 12318 5956
rect 12334 6012 12398 6016
rect 12334 5956 12338 6012
rect 12338 5956 12394 6012
rect 12394 5956 12398 6012
rect 12334 5952 12398 5956
rect 19522 6012 19586 6016
rect 19522 5956 19526 6012
rect 19526 5956 19582 6012
rect 19582 5956 19586 6012
rect 19522 5952 19586 5956
rect 19602 6012 19666 6016
rect 19602 5956 19606 6012
rect 19606 5956 19662 6012
rect 19662 5956 19666 6012
rect 19602 5952 19666 5956
rect 19682 6012 19746 6016
rect 19682 5956 19686 6012
rect 19686 5956 19742 6012
rect 19742 5956 19746 6012
rect 19682 5952 19746 5956
rect 19762 6012 19826 6016
rect 19762 5956 19766 6012
rect 19766 5956 19822 6012
rect 19822 5956 19826 6012
rect 19762 5952 19826 5956
rect 26950 6012 27014 6016
rect 26950 5956 26954 6012
rect 26954 5956 27010 6012
rect 27010 5956 27014 6012
rect 26950 5952 27014 5956
rect 27030 6012 27094 6016
rect 27030 5956 27034 6012
rect 27034 5956 27090 6012
rect 27090 5956 27094 6012
rect 27030 5952 27094 5956
rect 27110 6012 27174 6016
rect 27110 5956 27114 6012
rect 27114 5956 27170 6012
rect 27170 5956 27174 6012
rect 27110 5952 27174 5956
rect 27190 6012 27254 6016
rect 27190 5956 27194 6012
rect 27194 5956 27250 6012
rect 27250 5956 27254 6012
rect 27190 5952 27254 5956
rect 5326 5468 5390 5472
rect 5326 5412 5330 5468
rect 5330 5412 5386 5468
rect 5386 5412 5390 5468
rect 5326 5408 5390 5412
rect 5406 5468 5470 5472
rect 5406 5412 5410 5468
rect 5410 5412 5466 5468
rect 5466 5412 5470 5468
rect 5406 5408 5470 5412
rect 5486 5468 5550 5472
rect 5486 5412 5490 5468
rect 5490 5412 5546 5468
rect 5546 5412 5550 5468
rect 5486 5408 5550 5412
rect 5566 5468 5630 5472
rect 5566 5412 5570 5468
rect 5570 5412 5626 5468
rect 5626 5412 5630 5468
rect 5566 5408 5630 5412
rect 12754 5468 12818 5472
rect 12754 5412 12758 5468
rect 12758 5412 12814 5468
rect 12814 5412 12818 5468
rect 12754 5408 12818 5412
rect 12834 5468 12898 5472
rect 12834 5412 12838 5468
rect 12838 5412 12894 5468
rect 12894 5412 12898 5468
rect 12834 5408 12898 5412
rect 12914 5468 12978 5472
rect 12914 5412 12918 5468
rect 12918 5412 12974 5468
rect 12974 5412 12978 5468
rect 12914 5408 12978 5412
rect 12994 5468 13058 5472
rect 12994 5412 12998 5468
rect 12998 5412 13054 5468
rect 13054 5412 13058 5468
rect 12994 5408 13058 5412
rect 20182 5468 20246 5472
rect 20182 5412 20186 5468
rect 20186 5412 20242 5468
rect 20242 5412 20246 5468
rect 20182 5408 20246 5412
rect 20262 5468 20326 5472
rect 20262 5412 20266 5468
rect 20266 5412 20322 5468
rect 20322 5412 20326 5468
rect 20262 5408 20326 5412
rect 20342 5468 20406 5472
rect 20342 5412 20346 5468
rect 20346 5412 20402 5468
rect 20402 5412 20406 5468
rect 20342 5408 20406 5412
rect 20422 5468 20486 5472
rect 20422 5412 20426 5468
rect 20426 5412 20482 5468
rect 20482 5412 20486 5468
rect 20422 5408 20486 5412
rect 27610 5468 27674 5472
rect 27610 5412 27614 5468
rect 27614 5412 27670 5468
rect 27670 5412 27674 5468
rect 27610 5408 27674 5412
rect 27690 5468 27754 5472
rect 27690 5412 27694 5468
rect 27694 5412 27750 5468
rect 27750 5412 27754 5468
rect 27690 5408 27754 5412
rect 27770 5468 27834 5472
rect 27770 5412 27774 5468
rect 27774 5412 27830 5468
rect 27830 5412 27834 5468
rect 27770 5408 27834 5412
rect 27850 5468 27914 5472
rect 27850 5412 27854 5468
rect 27854 5412 27910 5468
rect 27910 5412 27914 5468
rect 27850 5408 27914 5412
rect 4666 4924 4730 4928
rect 4666 4868 4670 4924
rect 4670 4868 4726 4924
rect 4726 4868 4730 4924
rect 4666 4864 4730 4868
rect 4746 4924 4810 4928
rect 4746 4868 4750 4924
rect 4750 4868 4806 4924
rect 4806 4868 4810 4924
rect 4746 4864 4810 4868
rect 4826 4924 4890 4928
rect 4826 4868 4830 4924
rect 4830 4868 4886 4924
rect 4886 4868 4890 4924
rect 4826 4864 4890 4868
rect 4906 4924 4970 4928
rect 4906 4868 4910 4924
rect 4910 4868 4966 4924
rect 4966 4868 4970 4924
rect 4906 4864 4970 4868
rect 12094 4924 12158 4928
rect 12094 4868 12098 4924
rect 12098 4868 12154 4924
rect 12154 4868 12158 4924
rect 12094 4864 12158 4868
rect 12174 4924 12238 4928
rect 12174 4868 12178 4924
rect 12178 4868 12234 4924
rect 12234 4868 12238 4924
rect 12174 4864 12238 4868
rect 12254 4924 12318 4928
rect 12254 4868 12258 4924
rect 12258 4868 12314 4924
rect 12314 4868 12318 4924
rect 12254 4864 12318 4868
rect 12334 4924 12398 4928
rect 12334 4868 12338 4924
rect 12338 4868 12394 4924
rect 12394 4868 12398 4924
rect 12334 4864 12398 4868
rect 19522 4924 19586 4928
rect 19522 4868 19526 4924
rect 19526 4868 19582 4924
rect 19582 4868 19586 4924
rect 19522 4864 19586 4868
rect 19602 4924 19666 4928
rect 19602 4868 19606 4924
rect 19606 4868 19662 4924
rect 19662 4868 19666 4924
rect 19602 4864 19666 4868
rect 19682 4924 19746 4928
rect 19682 4868 19686 4924
rect 19686 4868 19742 4924
rect 19742 4868 19746 4924
rect 19682 4864 19746 4868
rect 19762 4924 19826 4928
rect 19762 4868 19766 4924
rect 19766 4868 19822 4924
rect 19822 4868 19826 4924
rect 19762 4864 19826 4868
rect 26950 4924 27014 4928
rect 26950 4868 26954 4924
rect 26954 4868 27010 4924
rect 27010 4868 27014 4924
rect 26950 4864 27014 4868
rect 27030 4924 27094 4928
rect 27030 4868 27034 4924
rect 27034 4868 27090 4924
rect 27090 4868 27094 4924
rect 27030 4864 27094 4868
rect 27110 4924 27174 4928
rect 27110 4868 27114 4924
rect 27114 4868 27170 4924
rect 27170 4868 27174 4924
rect 27110 4864 27174 4868
rect 27190 4924 27254 4928
rect 27190 4868 27194 4924
rect 27194 4868 27250 4924
rect 27250 4868 27254 4924
rect 27190 4864 27254 4868
rect 5326 4380 5390 4384
rect 5326 4324 5330 4380
rect 5330 4324 5386 4380
rect 5386 4324 5390 4380
rect 5326 4320 5390 4324
rect 5406 4380 5470 4384
rect 5406 4324 5410 4380
rect 5410 4324 5466 4380
rect 5466 4324 5470 4380
rect 5406 4320 5470 4324
rect 5486 4380 5550 4384
rect 5486 4324 5490 4380
rect 5490 4324 5546 4380
rect 5546 4324 5550 4380
rect 5486 4320 5550 4324
rect 5566 4380 5630 4384
rect 5566 4324 5570 4380
rect 5570 4324 5626 4380
rect 5626 4324 5630 4380
rect 5566 4320 5630 4324
rect 12754 4380 12818 4384
rect 12754 4324 12758 4380
rect 12758 4324 12814 4380
rect 12814 4324 12818 4380
rect 12754 4320 12818 4324
rect 12834 4380 12898 4384
rect 12834 4324 12838 4380
rect 12838 4324 12894 4380
rect 12894 4324 12898 4380
rect 12834 4320 12898 4324
rect 12914 4380 12978 4384
rect 12914 4324 12918 4380
rect 12918 4324 12974 4380
rect 12974 4324 12978 4380
rect 12914 4320 12978 4324
rect 12994 4380 13058 4384
rect 12994 4324 12998 4380
rect 12998 4324 13054 4380
rect 13054 4324 13058 4380
rect 12994 4320 13058 4324
rect 20182 4380 20246 4384
rect 20182 4324 20186 4380
rect 20186 4324 20242 4380
rect 20242 4324 20246 4380
rect 20182 4320 20246 4324
rect 20262 4380 20326 4384
rect 20262 4324 20266 4380
rect 20266 4324 20322 4380
rect 20322 4324 20326 4380
rect 20262 4320 20326 4324
rect 20342 4380 20406 4384
rect 20342 4324 20346 4380
rect 20346 4324 20402 4380
rect 20402 4324 20406 4380
rect 20342 4320 20406 4324
rect 20422 4380 20486 4384
rect 20422 4324 20426 4380
rect 20426 4324 20482 4380
rect 20482 4324 20486 4380
rect 20422 4320 20486 4324
rect 27610 4380 27674 4384
rect 27610 4324 27614 4380
rect 27614 4324 27670 4380
rect 27670 4324 27674 4380
rect 27610 4320 27674 4324
rect 27690 4380 27754 4384
rect 27690 4324 27694 4380
rect 27694 4324 27750 4380
rect 27750 4324 27754 4380
rect 27690 4320 27754 4324
rect 27770 4380 27834 4384
rect 27770 4324 27774 4380
rect 27774 4324 27830 4380
rect 27830 4324 27834 4380
rect 27770 4320 27834 4324
rect 27850 4380 27914 4384
rect 27850 4324 27854 4380
rect 27854 4324 27910 4380
rect 27910 4324 27914 4380
rect 27850 4320 27914 4324
rect 4666 3836 4730 3840
rect 4666 3780 4670 3836
rect 4670 3780 4726 3836
rect 4726 3780 4730 3836
rect 4666 3776 4730 3780
rect 4746 3836 4810 3840
rect 4746 3780 4750 3836
rect 4750 3780 4806 3836
rect 4806 3780 4810 3836
rect 4746 3776 4810 3780
rect 4826 3836 4890 3840
rect 4826 3780 4830 3836
rect 4830 3780 4886 3836
rect 4886 3780 4890 3836
rect 4826 3776 4890 3780
rect 4906 3836 4970 3840
rect 4906 3780 4910 3836
rect 4910 3780 4966 3836
rect 4966 3780 4970 3836
rect 4906 3776 4970 3780
rect 12094 3836 12158 3840
rect 12094 3780 12098 3836
rect 12098 3780 12154 3836
rect 12154 3780 12158 3836
rect 12094 3776 12158 3780
rect 12174 3836 12238 3840
rect 12174 3780 12178 3836
rect 12178 3780 12234 3836
rect 12234 3780 12238 3836
rect 12174 3776 12238 3780
rect 12254 3836 12318 3840
rect 12254 3780 12258 3836
rect 12258 3780 12314 3836
rect 12314 3780 12318 3836
rect 12254 3776 12318 3780
rect 12334 3836 12398 3840
rect 12334 3780 12338 3836
rect 12338 3780 12394 3836
rect 12394 3780 12398 3836
rect 12334 3776 12398 3780
rect 19522 3836 19586 3840
rect 19522 3780 19526 3836
rect 19526 3780 19582 3836
rect 19582 3780 19586 3836
rect 19522 3776 19586 3780
rect 19602 3836 19666 3840
rect 19602 3780 19606 3836
rect 19606 3780 19662 3836
rect 19662 3780 19666 3836
rect 19602 3776 19666 3780
rect 19682 3836 19746 3840
rect 19682 3780 19686 3836
rect 19686 3780 19742 3836
rect 19742 3780 19746 3836
rect 19682 3776 19746 3780
rect 19762 3836 19826 3840
rect 19762 3780 19766 3836
rect 19766 3780 19822 3836
rect 19822 3780 19826 3836
rect 19762 3776 19826 3780
rect 26950 3836 27014 3840
rect 26950 3780 26954 3836
rect 26954 3780 27010 3836
rect 27010 3780 27014 3836
rect 26950 3776 27014 3780
rect 27030 3836 27094 3840
rect 27030 3780 27034 3836
rect 27034 3780 27090 3836
rect 27090 3780 27094 3836
rect 27030 3776 27094 3780
rect 27110 3836 27174 3840
rect 27110 3780 27114 3836
rect 27114 3780 27170 3836
rect 27170 3780 27174 3836
rect 27110 3776 27174 3780
rect 27190 3836 27254 3840
rect 27190 3780 27194 3836
rect 27194 3780 27250 3836
rect 27250 3780 27254 3836
rect 27190 3776 27254 3780
rect 5326 3292 5390 3296
rect 5326 3236 5330 3292
rect 5330 3236 5386 3292
rect 5386 3236 5390 3292
rect 5326 3232 5390 3236
rect 5406 3292 5470 3296
rect 5406 3236 5410 3292
rect 5410 3236 5466 3292
rect 5466 3236 5470 3292
rect 5406 3232 5470 3236
rect 5486 3292 5550 3296
rect 5486 3236 5490 3292
rect 5490 3236 5546 3292
rect 5546 3236 5550 3292
rect 5486 3232 5550 3236
rect 5566 3292 5630 3296
rect 5566 3236 5570 3292
rect 5570 3236 5626 3292
rect 5626 3236 5630 3292
rect 5566 3232 5630 3236
rect 12754 3292 12818 3296
rect 12754 3236 12758 3292
rect 12758 3236 12814 3292
rect 12814 3236 12818 3292
rect 12754 3232 12818 3236
rect 12834 3292 12898 3296
rect 12834 3236 12838 3292
rect 12838 3236 12894 3292
rect 12894 3236 12898 3292
rect 12834 3232 12898 3236
rect 12914 3292 12978 3296
rect 12914 3236 12918 3292
rect 12918 3236 12974 3292
rect 12974 3236 12978 3292
rect 12914 3232 12978 3236
rect 12994 3292 13058 3296
rect 12994 3236 12998 3292
rect 12998 3236 13054 3292
rect 13054 3236 13058 3292
rect 12994 3232 13058 3236
rect 20182 3292 20246 3296
rect 20182 3236 20186 3292
rect 20186 3236 20242 3292
rect 20242 3236 20246 3292
rect 20182 3232 20246 3236
rect 20262 3292 20326 3296
rect 20262 3236 20266 3292
rect 20266 3236 20322 3292
rect 20322 3236 20326 3292
rect 20262 3232 20326 3236
rect 20342 3292 20406 3296
rect 20342 3236 20346 3292
rect 20346 3236 20402 3292
rect 20402 3236 20406 3292
rect 20342 3232 20406 3236
rect 20422 3292 20486 3296
rect 20422 3236 20426 3292
rect 20426 3236 20482 3292
rect 20482 3236 20486 3292
rect 20422 3232 20486 3236
rect 27610 3292 27674 3296
rect 27610 3236 27614 3292
rect 27614 3236 27670 3292
rect 27670 3236 27674 3292
rect 27610 3232 27674 3236
rect 27690 3292 27754 3296
rect 27690 3236 27694 3292
rect 27694 3236 27750 3292
rect 27750 3236 27754 3292
rect 27690 3232 27754 3236
rect 27770 3292 27834 3296
rect 27770 3236 27774 3292
rect 27774 3236 27830 3292
rect 27830 3236 27834 3292
rect 27770 3232 27834 3236
rect 27850 3292 27914 3296
rect 27850 3236 27854 3292
rect 27854 3236 27910 3292
rect 27910 3236 27914 3292
rect 27850 3232 27914 3236
rect 4666 2748 4730 2752
rect 4666 2692 4670 2748
rect 4670 2692 4726 2748
rect 4726 2692 4730 2748
rect 4666 2688 4730 2692
rect 4746 2748 4810 2752
rect 4746 2692 4750 2748
rect 4750 2692 4806 2748
rect 4806 2692 4810 2748
rect 4746 2688 4810 2692
rect 4826 2748 4890 2752
rect 4826 2692 4830 2748
rect 4830 2692 4886 2748
rect 4886 2692 4890 2748
rect 4826 2688 4890 2692
rect 4906 2748 4970 2752
rect 4906 2692 4910 2748
rect 4910 2692 4966 2748
rect 4966 2692 4970 2748
rect 4906 2688 4970 2692
rect 12094 2748 12158 2752
rect 12094 2692 12098 2748
rect 12098 2692 12154 2748
rect 12154 2692 12158 2748
rect 12094 2688 12158 2692
rect 12174 2748 12238 2752
rect 12174 2692 12178 2748
rect 12178 2692 12234 2748
rect 12234 2692 12238 2748
rect 12174 2688 12238 2692
rect 12254 2748 12318 2752
rect 12254 2692 12258 2748
rect 12258 2692 12314 2748
rect 12314 2692 12318 2748
rect 12254 2688 12318 2692
rect 12334 2748 12398 2752
rect 12334 2692 12338 2748
rect 12338 2692 12394 2748
rect 12394 2692 12398 2748
rect 12334 2688 12398 2692
rect 19522 2748 19586 2752
rect 19522 2692 19526 2748
rect 19526 2692 19582 2748
rect 19582 2692 19586 2748
rect 19522 2688 19586 2692
rect 19602 2748 19666 2752
rect 19602 2692 19606 2748
rect 19606 2692 19662 2748
rect 19662 2692 19666 2748
rect 19602 2688 19666 2692
rect 19682 2748 19746 2752
rect 19682 2692 19686 2748
rect 19686 2692 19742 2748
rect 19742 2692 19746 2748
rect 19682 2688 19746 2692
rect 19762 2748 19826 2752
rect 19762 2692 19766 2748
rect 19766 2692 19822 2748
rect 19822 2692 19826 2748
rect 19762 2688 19826 2692
rect 26950 2748 27014 2752
rect 26950 2692 26954 2748
rect 26954 2692 27010 2748
rect 27010 2692 27014 2748
rect 26950 2688 27014 2692
rect 27030 2748 27094 2752
rect 27030 2692 27034 2748
rect 27034 2692 27090 2748
rect 27090 2692 27094 2748
rect 27030 2688 27094 2692
rect 27110 2748 27174 2752
rect 27110 2692 27114 2748
rect 27114 2692 27170 2748
rect 27170 2692 27174 2748
rect 27110 2688 27174 2692
rect 27190 2748 27254 2752
rect 27190 2692 27194 2748
rect 27194 2692 27250 2748
rect 27250 2692 27254 2748
rect 27190 2688 27254 2692
rect 5326 2204 5390 2208
rect 5326 2148 5330 2204
rect 5330 2148 5386 2204
rect 5386 2148 5390 2204
rect 5326 2144 5390 2148
rect 5406 2204 5470 2208
rect 5406 2148 5410 2204
rect 5410 2148 5466 2204
rect 5466 2148 5470 2204
rect 5406 2144 5470 2148
rect 5486 2204 5550 2208
rect 5486 2148 5490 2204
rect 5490 2148 5546 2204
rect 5546 2148 5550 2204
rect 5486 2144 5550 2148
rect 5566 2204 5630 2208
rect 5566 2148 5570 2204
rect 5570 2148 5626 2204
rect 5626 2148 5630 2204
rect 5566 2144 5630 2148
rect 12754 2204 12818 2208
rect 12754 2148 12758 2204
rect 12758 2148 12814 2204
rect 12814 2148 12818 2204
rect 12754 2144 12818 2148
rect 12834 2204 12898 2208
rect 12834 2148 12838 2204
rect 12838 2148 12894 2204
rect 12894 2148 12898 2204
rect 12834 2144 12898 2148
rect 12914 2204 12978 2208
rect 12914 2148 12918 2204
rect 12918 2148 12974 2204
rect 12974 2148 12978 2204
rect 12914 2144 12978 2148
rect 12994 2204 13058 2208
rect 12994 2148 12998 2204
rect 12998 2148 13054 2204
rect 13054 2148 13058 2204
rect 12994 2144 13058 2148
rect 20182 2204 20246 2208
rect 20182 2148 20186 2204
rect 20186 2148 20242 2204
rect 20242 2148 20246 2204
rect 20182 2144 20246 2148
rect 20262 2204 20326 2208
rect 20262 2148 20266 2204
rect 20266 2148 20322 2204
rect 20322 2148 20326 2204
rect 20262 2144 20326 2148
rect 20342 2204 20406 2208
rect 20342 2148 20346 2204
rect 20346 2148 20402 2204
rect 20402 2148 20406 2204
rect 20342 2144 20406 2148
rect 20422 2204 20486 2208
rect 20422 2148 20426 2204
rect 20426 2148 20482 2204
rect 20482 2148 20486 2204
rect 20422 2144 20486 2148
rect 27610 2204 27674 2208
rect 27610 2148 27614 2204
rect 27614 2148 27670 2204
rect 27670 2148 27674 2204
rect 27610 2144 27674 2148
rect 27690 2204 27754 2208
rect 27690 2148 27694 2204
rect 27694 2148 27750 2204
rect 27750 2148 27754 2204
rect 27690 2144 27754 2148
rect 27770 2204 27834 2208
rect 27770 2148 27774 2204
rect 27774 2148 27830 2204
rect 27830 2148 27834 2204
rect 27770 2144 27834 2148
rect 27850 2204 27914 2208
rect 27850 2148 27854 2204
rect 27854 2148 27910 2204
rect 27910 2148 27914 2204
rect 27850 2144 27914 2148
<< metal4 >>
rect 4658 28864 4978 29424
rect 4658 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4978 28864
rect 4658 27776 4978 28800
rect 4658 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4978 27776
rect 4658 26688 4978 27712
rect 4658 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4978 26688
rect 4658 26094 4978 26624
rect 4658 25858 4700 26094
rect 4936 25858 4978 26094
rect 4658 25600 4978 25858
rect 4658 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4978 25600
rect 4658 24512 4978 25536
rect 4658 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4978 24512
rect 4658 23424 4978 24448
rect 4658 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4978 23424
rect 4658 22336 4978 23360
rect 4658 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4978 22336
rect 4658 21248 4978 22272
rect 4658 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4978 21248
rect 4658 20160 4978 21184
rect 4658 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4978 20160
rect 4658 19294 4978 20096
rect 4658 19072 4700 19294
rect 4936 19072 4978 19294
rect 4658 19008 4666 19072
rect 4730 19008 4746 19058
rect 4810 19008 4826 19058
rect 4890 19008 4906 19058
rect 4970 19008 4978 19072
rect 4658 17984 4978 19008
rect 4658 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4978 17984
rect 4658 16896 4978 17920
rect 4658 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4978 16896
rect 4658 15808 4978 16832
rect 4658 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4978 15808
rect 4658 14720 4978 15744
rect 4658 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4978 14720
rect 4658 13632 4978 14656
rect 4658 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4978 13632
rect 4658 12544 4978 13568
rect 4658 12480 4666 12544
rect 4730 12494 4746 12544
rect 4810 12494 4826 12544
rect 4890 12494 4906 12544
rect 4970 12480 4978 12544
rect 4658 12258 4700 12480
rect 4936 12258 4978 12480
rect 4658 11456 4978 12258
rect 4658 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4978 11456
rect 4658 10368 4978 11392
rect 4658 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4978 10368
rect 4658 9280 4978 10304
rect 4658 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4978 9280
rect 4658 8192 4978 9216
rect 4658 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4978 8192
rect 4658 7104 4978 8128
rect 4658 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4978 7104
rect 4658 6016 4978 7040
rect 4658 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4978 6016
rect 4658 5694 4978 5952
rect 4658 5458 4700 5694
rect 4936 5458 4978 5694
rect 4658 4928 4978 5458
rect 4658 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4978 4928
rect 4658 3840 4978 4864
rect 4658 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4978 3840
rect 4658 2752 4978 3776
rect 4658 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4978 2752
rect 4658 2128 4978 2688
rect 5318 29408 5638 29424
rect 5318 29344 5326 29408
rect 5390 29344 5406 29408
rect 5470 29344 5486 29408
rect 5550 29344 5566 29408
rect 5630 29344 5638 29408
rect 5318 28320 5638 29344
rect 5318 28256 5326 28320
rect 5390 28256 5406 28320
rect 5470 28256 5486 28320
rect 5550 28256 5566 28320
rect 5630 28256 5638 28320
rect 5318 27232 5638 28256
rect 5318 27168 5326 27232
rect 5390 27168 5406 27232
rect 5470 27168 5486 27232
rect 5550 27168 5566 27232
rect 5630 27168 5638 27232
rect 5318 26754 5638 27168
rect 5318 26518 5360 26754
rect 5596 26518 5638 26754
rect 5318 26144 5638 26518
rect 5318 26080 5326 26144
rect 5390 26080 5406 26144
rect 5470 26080 5486 26144
rect 5550 26080 5566 26144
rect 5630 26080 5638 26144
rect 5318 25056 5638 26080
rect 5318 24992 5326 25056
rect 5390 24992 5406 25056
rect 5470 24992 5486 25056
rect 5550 24992 5566 25056
rect 5630 24992 5638 25056
rect 5318 23968 5638 24992
rect 5318 23904 5326 23968
rect 5390 23904 5406 23968
rect 5470 23904 5486 23968
rect 5550 23904 5566 23968
rect 5630 23904 5638 23968
rect 5318 22880 5638 23904
rect 5318 22816 5326 22880
rect 5390 22816 5406 22880
rect 5470 22816 5486 22880
rect 5550 22816 5566 22880
rect 5630 22816 5638 22880
rect 5318 21792 5638 22816
rect 5318 21728 5326 21792
rect 5390 21728 5406 21792
rect 5470 21728 5486 21792
rect 5550 21728 5566 21792
rect 5630 21728 5638 21792
rect 5318 20704 5638 21728
rect 5318 20640 5326 20704
rect 5390 20640 5406 20704
rect 5470 20640 5486 20704
rect 5550 20640 5566 20704
rect 5630 20640 5638 20704
rect 5318 19954 5638 20640
rect 5318 19718 5360 19954
rect 5596 19718 5638 19954
rect 5318 19616 5638 19718
rect 5318 19552 5326 19616
rect 5390 19552 5406 19616
rect 5470 19552 5486 19616
rect 5550 19552 5566 19616
rect 5630 19552 5638 19616
rect 5318 18528 5638 19552
rect 5318 18464 5326 18528
rect 5390 18464 5406 18528
rect 5470 18464 5486 18528
rect 5550 18464 5566 18528
rect 5630 18464 5638 18528
rect 5318 17440 5638 18464
rect 5318 17376 5326 17440
rect 5390 17376 5406 17440
rect 5470 17376 5486 17440
rect 5550 17376 5566 17440
rect 5630 17376 5638 17440
rect 5318 16352 5638 17376
rect 5318 16288 5326 16352
rect 5390 16288 5406 16352
rect 5470 16288 5486 16352
rect 5550 16288 5566 16352
rect 5630 16288 5638 16352
rect 5318 15264 5638 16288
rect 5318 15200 5326 15264
rect 5390 15200 5406 15264
rect 5470 15200 5486 15264
rect 5550 15200 5566 15264
rect 5630 15200 5638 15264
rect 5318 14176 5638 15200
rect 5318 14112 5326 14176
rect 5390 14112 5406 14176
rect 5470 14112 5486 14176
rect 5550 14112 5566 14176
rect 5630 14112 5638 14176
rect 5318 13154 5638 14112
rect 5318 13088 5360 13154
rect 5596 13088 5638 13154
rect 5318 13024 5326 13088
rect 5630 13024 5638 13088
rect 5318 12918 5360 13024
rect 5596 12918 5638 13024
rect 5318 12000 5638 12918
rect 5318 11936 5326 12000
rect 5390 11936 5406 12000
rect 5470 11936 5486 12000
rect 5550 11936 5566 12000
rect 5630 11936 5638 12000
rect 5318 10912 5638 11936
rect 5318 10848 5326 10912
rect 5390 10848 5406 10912
rect 5470 10848 5486 10912
rect 5550 10848 5566 10912
rect 5630 10848 5638 10912
rect 5318 9824 5638 10848
rect 5318 9760 5326 9824
rect 5390 9760 5406 9824
rect 5470 9760 5486 9824
rect 5550 9760 5566 9824
rect 5630 9760 5638 9824
rect 5318 8736 5638 9760
rect 5318 8672 5326 8736
rect 5390 8672 5406 8736
rect 5470 8672 5486 8736
rect 5550 8672 5566 8736
rect 5630 8672 5638 8736
rect 5318 7648 5638 8672
rect 5318 7584 5326 7648
rect 5390 7584 5406 7648
rect 5470 7584 5486 7648
rect 5550 7584 5566 7648
rect 5630 7584 5638 7648
rect 5318 6560 5638 7584
rect 5318 6496 5326 6560
rect 5390 6496 5406 6560
rect 5470 6496 5486 6560
rect 5550 6496 5566 6560
rect 5630 6496 5638 6560
rect 5318 6354 5638 6496
rect 5318 6118 5360 6354
rect 5596 6118 5638 6354
rect 5318 5472 5638 6118
rect 5318 5408 5326 5472
rect 5390 5408 5406 5472
rect 5470 5408 5486 5472
rect 5550 5408 5566 5472
rect 5630 5408 5638 5472
rect 5318 4384 5638 5408
rect 5318 4320 5326 4384
rect 5390 4320 5406 4384
rect 5470 4320 5486 4384
rect 5550 4320 5566 4384
rect 5630 4320 5638 4384
rect 5318 3296 5638 4320
rect 5318 3232 5326 3296
rect 5390 3232 5406 3296
rect 5470 3232 5486 3296
rect 5550 3232 5566 3296
rect 5630 3232 5638 3296
rect 5318 2208 5638 3232
rect 5318 2144 5326 2208
rect 5390 2144 5406 2208
rect 5470 2144 5486 2208
rect 5550 2144 5566 2208
rect 5630 2144 5638 2208
rect 5318 2128 5638 2144
rect 12086 28864 12406 29424
rect 12086 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12406 28864
rect 12086 27776 12406 28800
rect 12086 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12406 27776
rect 12086 26688 12406 27712
rect 12086 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12406 26688
rect 12086 26094 12406 26624
rect 12086 25858 12128 26094
rect 12364 25858 12406 26094
rect 12086 25600 12406 25858
rect 12086 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12406 25600
rect 12086 24512 12406 25536
rect 12086 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12406 24512
rect 12086 23424 12406 24448
rect 12086 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12406 23424
rect 12086 22336 12406 23360
rect 12086 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12406 22336
rect 12086 21248 12406 22272
rect 12086 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12406 21248
rect 12086 20160 12406 21184
rect 12086 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12406 20160
rect 12086 19294 12406 20096
rect 12086 19072 12128 19294
rect 12364 19072 12406 19294
rect 12086 19008 12094 19072
rect 12158 19008 12174 19058
rect 12238 19008 12254 19058
rect 12318 19008 12334 19058
rect 12398 19008 12406 19072
rect 12086 17984 12406 19008
rect 12086 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12406 17984
rect 12086 16896 12406 17920
rect 12086 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12406 16896
rect 12086 15808 12406 16832
rect 12086 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12406 15808
rect 12086 14720 12406 15744
rect 12086 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12406 14720
rect 12086 13632 12406 14656
rect 12086 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12406 13632
rect 12086 12544 12406 13568
rect 12086 12480 12094 12544
rect 12158 12494 12174 12544
rect 12238 12494 12254 12544
rect 12318 12494 12334 12544
rect 12398 12480 12406 12544
rect 12086 12258 12128 12480
rect 12364 12258 12406 12480
rect 12086 11456 12406 12258
rect 12086 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12406 11456
rect 12086 10368 12406 11392
rect 12086 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12406 10368
rect 12086 9280 12406 10304
rect 12086 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12406 9280
rect 12086 8192 12406 9216
rect 12086 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12406 8192
rect 12086 7104 12406 8128
rect 12086 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12406 7104
rect 12086 6016 12406 7040
rect 12086 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12406 6016
rect 12086 5694 12406 5952
rect 12086 5458 12128 5694
rect 12364 5458 12406 5694
rect 12086 4928 12406 5458
rect 12086 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12406 4928
rect 12086 3840 12406 4864
rect 12086 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12406 3840
rect 12086 2752 12406 3776
rect 12086 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12406 2752
rect 12086 2128 12406 2688
rect 12746 29408 13066 29424
rect 12746 29344 12754 29408
rect 12818 29344 12834 29408
rect 12898 29344 12914 29408
rect 12978 29344 12994 29408
rect 13058 29344 13066 29408
rect 12746 28320 13066 29344
rect 12746 28256 12754 28320
rect 12818 28256 12834 28320
rect 12898 28256 12914 28320
rect 12978 28256 12994 28320
rect 13058 28256 13066 28320
rect 12746 27232 13066 28256
rect 12746 27168 12754 27232
rect 12818 27168 12834 27232
rect 12898 27168 12914 27232
rect 12978 27168 12994 27232
rect 13058 27168 13066 27232
rect 12746 26754 13066 27168
rect 12746 26518 12788 26754
rect 13024 26518 13066 26754
rect 12746 26144 13066 26518
rect 12746 26080 12754 26144
rect 12818 26080 12834 26144
rect 12898 26080 12914 26144
rect 12978 26080 12994 26144
rect 13058 26080 13066 26144
rect 12746 25056 13066 26080
rect 12746 24992 12754 25056
rect 12818 24992 12834 25056
rect 12898 24992 12914 25056
rect 12978 24992 12994 25056
rect 13058 24992 13066 25056
rect 12746 23968 13066 24992
rect 12746 23904 12754 23968
rect 12818 23904 12834 23968
rect 12898 23904 12914 23968
rect 12978 23904 12994 23968
rect 13058 23904 13066 23968
rect 12746 22880 13066 23904
rect 12746 22816 12754 22880
rect 12818 22816 12834 22880
rect 12898 22816 12914 22880
rect 12978 22816 12994 22880
rect 13058 22816 13066 22880
rect 12746 21792 13066 22816
rect 12746 21728 12754 21792
rect 12818 21728 12834 21792
rect 12898 21728 12914 21792
rect 12978 21728 12994 21792
rect 13058 21728 13066 21792
rect 12746 20704 13066 21728
rect 12746 20640 12754 20704
rect 12818 20640 12834 20704
rect 12898 20640 12914 20704
rect 12978 20640 12994 20704
rect 13058 20640 13066 20704
rect 12746 19954 13066 20640
rect 12746 19718 12788 19954
rect 13024 19718 13066 19954
rect 12746 19616 13066 19718
rect 12746 19552 12754 19616
rect 12818 19552 12834 19616
rect 12898 19552 12914 19616
rect 12978 19552 12994 19616
rect 13058 19552 13066 19616
rect 12746 18528 13066 19552
rect 12746 18464 12754 18528
rect 12818 18464 12834 18528
rect 12898 18464 12914 18528
rect 12978 18464 12994 18528
rect 13058 18464 13066 18528
rect 12746 17440 13066 18464
rect 12746 17376 12754 17440
rect 12818 17376 12834 17440
rect 12898 17376 12914 17440
rect 12978 17376 12994 17440
rect 13058 17376 13066 17440
rect 12746 16352 13066 17376
rect 12746 16288 12754 16352
rect 12818 16288 12834 16352
rect 12898 16288 12914 16352
rect 12978 16288 12994 16352
rect 13058 16288 13066 16352
rect 12746 15264 13066 16288
rect 12746 15200 12754 15264
rect 12818 15200 12834 15264
rect 12898 15200 12914 15264
rect 12978 15200 12994 15264
rect 13058 15200 13066 15264
rect 12746 14176 13066 15200
rect 12746 14112 12754 14176
rect 12818 14112 12834 14176
rect 12898 14112 12914 14176
rect 12978 14112 12994 14176
rect 13058 14112 13066 14176
rect 12746 13154 13066 14112
rect 12746 13088 12788 13154
rect 13024 13088 13066 13154
rect 12746 13024 12754 13088
rect 13058 13024 13066 13088
rect 12746 12918 12788 13024
rect 13024 12918 13066 13024
rect 12746 12000 13066 12918
rect 12746 11936 12754 12000
rect 12818 11936 12834 12000
rect 12898 11936 12914 12000
rect 12978 11936 12994 12000
rect 13058 11936 13066 12000
rect 12746 10912 13066 11936
rect 12746 10848 12754 10912
rect 12818 10848 12834 10912
rect 12898 10848 12914 10912
rect 12978 10848 12994 10912
rect 13058 10848 13066 10912
rect 12746 9824 13066 10848
rect 12746 9760 12754 9824
rect 12818 9760 12834 9824
rect 12898 9760 12914 9824
rect 12978 9760 12994 9824
rect 13058 9760 13066 9824
rect 12746 8736 13066 9760
rect 12746 8672 12754 8736
rect 12818 8672 12834 8736
rect 12898 8672 12914 8736
rect 12978 8672 12994 8736
rect 13058 8672 13066 8736
rect 12746 7648 13066 8672
rect 12746 7584 12754 7648
rect 12818 7584 12834 7648
rect 12898 7584 12914 7648
rect 12978 7584 12994 7648
rect 13058 7584 13066 7648
rect 12746 6560 13066 7584
rect 12746 6496 12754 6560
rect 12818 6496 12834 6560
rect 12898 6496 12914 6560
rect 12978 6496 12994 6560
rect 13058 6496 13066 6560
rect 12746 6354 13066 6496
rect 12746 6118 12788 6354
rect 13024 6118 13066 6354
rect 12746 5472 13066 6118
rect 12746 5408 12754 5472
rect 12818 5408 12834 5472
rect 12898 5408 12914 5472
rect 12978 5408 12994 5472
rect 13058 5408 13066 5472
rect 12746 4384 13066 5408
rect 12746 4320 12754 4384
rect 12818 4320 12834 4384
rect 12898 4320 12914 4384
rect 12978 4320 12994 4384
rect 13058 4320 13066 4384
rect 12746 3296 13066 4320
rect 12746 3232 12754 3296
rect 12818 3232 12834 3296
rect 12898 3232 12914 3296
rect 12978 3232 12994 3296
rect 13058 3232 13066 3296
rect 12746 2208 13066 3232
rect 12746 2144 12754 2208
rect 12818 2144 12834 2208
rect 12898 2144 12914 2208
rect 12978 2144 12994 2208
rect 13058 2144 13066 2208
rect 12746 2128 13066 2144
rect 19514 28864 19834 29424
rect 19514 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19834 28864
rect 19514 27776 19834 28800
rect 19514 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19834 27776
rect 19514 26688 19834 27712
rect 19514 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19834 26688
rect 19514 26094 19834 26624
rect 19514 25858 19556 26094
rect 19792 25858 19834 26094
rect 19514 25600 19834 25858
rect 19514 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19834 25600
rect 19514 24512 19834 25536
rect 19514 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19834 24512
rect 19514 23424 19834 24448
rect 19514 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19834 23424
rect 19514 22336 19834 23360
rect 19514 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19834 22336
rect 19514 21248 19834 22272
rect 19514 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19834 21248
rect 19514 20160 19834 21184
rect 19514 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19834 20160
rect 19514 19294 19834 20096
rect 19514 19072 19556 19294
rect 19792 19072 19834 19294
rect 19514 19008 19522 19072
rect 19586 19008 19602 19058
rect 19666 19008 19682 19058
rect 19746 19008 19762 19058
rect 19826 19008 19834 19072
rect 19514 17984 19834 19008
rect 19514 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19834 17984
rect 19514 16896 19834 17920
rect 19514 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19834 16896
rect 19514 15808 19834 16832
rect 19514 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19834 15808
rect 19514 14720 19834 15744
rect 19514 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19834 14720
rect 19514 13632 19834 14656
rect 19514 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19834 13632
rect 19514 12544 19834 13568
rect 19514 12480 19522 12544
rect 19586 12494 19602 12544
rect 19666 12494 19682 12544
rect 19746 12494 19762 12544
rect 19826 12480 19834 12544
rect 19514 12258 19556 12480
rect 19792 12258 19834 12480
rect 19514 11456 19834 12258
rect 19514 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19834 11456
rect 19514 10368 19834 11392
rect 19514 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19834 10368
rect 19514 9280 19834 10304
rect 19514 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19834 9280
rect 19514 8192 19834 9216
rect 19514 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19834 8192
rect 19514 7104 19834 8128
rect 19514 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19834 7104
rect 19514 6016 19834 7040
rect 19514 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19834 6016
rect 19514 5694 19834 5952
rect 19514 5458 19556 5694
rect 19792 5458 19834 5694
rect 19514 4928 19834 5458
rect 19514 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19834 4928
rect 19514 3840 19834 4864
rect 19514 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19834 3840
rect 19514 2752 19834 3776
rect 19514 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19834 2752
rect 19514 2128 19834 2688
rect 20174 29408 20494 29424
rect 20174 29344 20182 29408
rect 20246 29344 20262 29408
rect 20326 29344 20342 29408
rect 20406 29344 20422 29408
rect 20486 29344 20494 29408
rect 20174 28320 20494 29344
rect 20174 28256 20182 28320
rect 20246 28256 20262 28320
rect 20326 28256 20342 28320
rect 20406 28256 20422 28320
rect 20486 28256 20494 28320
rect 20174 27232 20494 28256
rect 20174 27168 20182 27232
rect 20246 27168 20262 27232
rect 20326 27168 20342 27232
rect 20406 27168 20422 27232
rect 20486 27168 20494 27232
rect 20174 26754 20494 27168
rect 20174 26518 20216 26754
rect 20452 26518 20494 26754
rect 20174 26144 20494 26518
rect 20174 26080 20182 26144
rect 20246 26080 20262 26144
rect 20326 26080 20342 26144
rect 20406 26080 20422 26144
rect 20486 26080 20494 26144
rect 20174 25056 20494 26080
rect 20174 24992 20182 25056
rect 20246 24992 20262 25056
rect 20326 24992 20342 25056
rect 20406 24992 20422 25056
rect 20486 24992 20494 25056
rect 20174 23968 20494 24992
rect 20174 23904 20182 23968
rect 20246 23904 20262 23968
rect 20326 23904 20342 23968
rect 20406 23904 20422 23968
rect 20486 23904 20494 23968
rect 20174 22880 20494 23904
rect 20174 22816 20182 22880
rect 20246 22816 20262 22880
rect 20326 22816 20342 22880
rect 20406 22816 20422 22880
rect 20486 22816 20494 22880
rect 20174 21792 20494 22816
rect 20174 21728 20182 21792
rect 20246 21728 20262 21792
rect 20326 21728 20342 21792
rect 20406 21728 20422 21792
rect 20486 21728 20494 21792
rect 20174 20704 20494 21728
rect 20174 20640 20182 20704
rect 20246 20640 20262 20704
rect 20326 20640 20342 20704
rect 20406 20640 20422 20704
rect 20486 20640 20494 20704
rect 20174 19954 20494 20640
rect 20174 19718 20216 19954
rect 20452 19718 20494 19954
rect 20174 19616 20494 19718
rect 20174 19552 20182 19616
rect 20246 19552 20262 19616
rect 20326 19552 20342 19616
rect 20406 19552 20422 19616
rect 20486 19552 20494 19616
rect 20174 18528 20494 19552
rect 20174 18464 20182 18528
rect 20246 18464 20262 18528
rect 20326 18464 20342 18528
rect 20406 18464 20422 18528
rect 20486 18464 20494 18528
rect 20174 17440 20494 18464
rect 20174 17376 20182 17440
rect 20246 17376 20262 17440
rect 20326 17376 20342 17440
rect 20406 17376 20422 17440
rect 20486 17376 20494 17440
rect 20174 16352 20494 17376
rect 20174 16288 20182 16352
rect 20246 16288 20262 16352
rect 20326 16288 20342 16352
rect 20406 16288 20422 16352
rect 20486 16288 20494 16352
rect 20174 15264 20494 16288
rect 20174 15200 20182 15264
rect 20246 15200 20262 15264
rect 20326 15200 20342 15264
rect 20406 15200 20422 15264
rect 20486 15200 20494 15264
rect 20174 14176 20494 15200
rect 20174 14112 20182 14176
rect 20246 14112 20262 14176
rect 20326 14112 20342 14176
rect 20406 14112 20422 14176
rect 20486 14112 20494 14176
rect 20174 13154 20494 14112
rect 20174 13088 20216 13154
rect 20452 13088 20494 13154
rect 20174 13024 20182 13088
rect 20486 13024 20494 13088
rect 20174 12918 20216 13024
rect 20452 12918 20494 13024
rect 20174 12000 20494 12918
rect 20174 11936 20182 12000
rect 20246 11936 20262 12000
rect 20326 11936 20342 12000
rect 20406 11936 20422 12000
rect 20486 11936 20494 12000
rect 20174 10912 20494 11936
rect 20174 10848 20182 10912
rect 20246 10848 20262 10912
rect 20326 10848 20342 10912
rect 20406 10848 20422 10912
rect 20486 10848 20494 10912
rect 20174 9824 20494 10848
rect 20174 9760 20182 9824
rect 20246 9760 20262 9824
rect 20326 9760 20342 9824
rect 20406 9760 20422 9824
rect 20486 9760 20494 9824
rect 20174 8736 20494 9760
rect 20174 8672 20182 8736
rect 20246 8672 20262 8736
rect 20326 8672 20342 8736
rect 20406 8672 20422 8736
rect 20486 8672 20494 8736
rect 20174 7648 20494 8672
rect 20174 7584 20182 7648
rect 20246 7584 20262 7648
rect 20326 7584 20342 7648
rect 20406 7584 20422 7648
rect 20486 7584 20494 7648
rect 20174 6560 20494 7584
rect 20174 6496 20182 6560
rect 20246 6496 20262 6560
rect 20326 6496 20342 6560
rect 20406 6496 20422 6560
rect 20486 6496 20494 6560
rect 20174 6354 20494 6496
rect 20174 6118 20216 6354
rect 20452 6118 20494 6354
rect 20174 5472 20494 6118
rect 20174 5408 20182 5472
rect 20246 5408 20262 5472
rect 20326 5408 20342 5472
rect 20406 5408 20422 5472
rect 20486 5408 20494 5472
rect 20174 4384 20494 5408
rect 20174 4320 20182 4384
rect 20246 4320 20262 4384
rect 20326 4320 20342 4384
rect 20406 4320 20422 4384
rect 20486 4320 20494 4384
rect 20174 3296 20494 4320
rect 20174 3232 20182 3296
rect 20246 3232 20262 3296
rect 20326 3232 20342 3296
rect 20406 3232 20422 3296
rect 20486 3232 20494 3296
rect 20174 2208 20494 3232
rect 20174 2144 20182 2208
rect 20246 2144 20262 2208
rect 20326 2144 20342 2208
rect 20406 2144 20422 2208
rect 20486 2144 20494 2208
rect 20174 2128 20494 2144
rect 26942 28864 27262 29424
rect 26942 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27262 28864
rect 26942 27776 27262 28800
rect 26942 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27262 27776
rect 26942 26688 27262 27712
rect 26942 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27262 26688
rect 26942 26094 27262 26624
rect 26942 25858 26984 26094
rect 27220 25858 27262 26094
rect 26942 25600 27262 25858
rect 26942 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27262 25600
rect 26942 24512 27262 25536
rect 26942 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27262 24512
rect 26942 23424 27262 24448
rect 26942 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27262 23424
rect 26942 22336 27262 23360
rect 26942 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27262 22336
rect 26942 21248 27262 22272
rect 26942 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27262 21248
rect 26942 20160 27262 21184
rect 26942 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27262 20160
rect 26942 19294 27262 20096
rect 26942 19072 26984 19294
rect 27220 19072 27262 19294
rect 26942 19008 26950 19072
rect 27014 19008 27030 19058
rect 27094 19008 27110 19058
rect 27174 19008 27190 19058
rect 27254 19008 27262 19072
rect 26942 17984 27262 19008
rect 26942 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27262 17984
rect 26942 16896 27262 17920
rect 26942 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27262 16896
rect 26942 15808 27262 16832
rect 26942 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27262 15808
rect 26942 14720 27262 15744
rect 26942 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27262 14720
rect 26942 13632 27262 14656
rect 26942 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27262 13632
rect 26942 12544 27262 13568
rect 26942 12480 26950 12544
rect 27014 12494 27030 12544
rect 27094 12494 27110 12544
rect 27174 12494 27190 12544
rect 27254 12480 27262 12544
rect 26942 12258 26984 12480
rect 27220 12258 27262 12480
rect 26942 11456 27262 12258
rect 26942 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27262 11456
rect 26942 10368 27262 11392
rect 26942 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27262 10368
rect 26942 9280 27262 10304
rect 26942 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27262 9280
rect 26942 8192 27262 9216
rect 26942 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27262 8192
rect 26942 7104 27262 8128
rect 26942 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27262 7104
rect 26942 6016 27262 7040
rect 26942 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27262 6016
rect 26942 5694 27262 5952
rect 26942 5458 26984 5694
rect 27220 5458 27262 5694
rect 26942 4928 27262 5458
rect 26942 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27262 4928
rect 26942 3840 27262 4864
rect 26942 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27262 3840
rect 26942 2752 27262 3776
rect 26942 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27262 2752
rect 26942 2128 27262 2688
rect 27602 29408 27922 29424
rect 27602 29344 27610 29408
rect 27674 29344 27690 29408
rect 27754 29344 27770 29408
rect 27834 29344 27850 29408
rect 27914 29344 27922 29408
rect 27602 28320 27922 29344
rect 27602 28256 27610 28320
rect 27674 28256 27690 28320
rect 27754 28256 27770 28320
rect 27834 28256 27850 28320
rect 27914 28256 27922 28320
rect 27602 27232 27922 28256
rect 27602 27168 27610 27232
rect 27674 27168 27690 27232
rect 27754 27168 27770 27232
rect 27834 27168 27850 27232
rect 27914 27168 27922 27232
rect 27602 26754 27922 27168
rect 27602 26518 27644 26754
rect 27880 26518 27922 26754
rect 27602 26144 27922 26518
rect 27602 26080 27610 26144
rect 27674 26080 27690 26144
rect 27754 26080 27770 26144
rect 27834 26080 27850 26144
rect 27914 26080 27922 26144
rect 27602 25056 27922 26080
rect 27602 24992 27610 25056
rect 27674 24992 27690 25056
rect 27754 24992 27770 25056
rect 27834 24992 27850 25056
rect 27914 24992 27922 25056
rect 27602 23968 27922 24992
rect 27602 23904 27610 23968
rect 27674 23904 27690 23968
rect 27754 23904 27770 23968
rect 27834 23904 27850 23968
rect 27914 23904 27922 23968
rect 27602 22880 27922 23904
rect 27602 22816 27610 22880
rect 27674 22816 27690 22880
rect 27754 22816 27770 22880
rect 27834 22816 27850 22880
rect 27914 22816 27922 22880
rect 27602 21792 27922 22816
rect 27602 21728 27610 21792
rect 27674 21728 27690 21792
rect 27754 21728 27770 21792
rect 27834 21728 27850 21792
rect 27914 21728 27922 21792
rect 27602 20704 27922 21728
rect 27602 20640 27610 20704
rect 27674 20640 27690 20704
rect 27754 20640 27770 20704
rect 27834 20640 27850 20704
rect 27914 20640 27922 20704
rect 27602 19954 27922 20640
rect 27602 19718 27644 19954
rect 27880 19718 27922 19954
rect 27602 19616 27922 19718
rect 27602 19552 27610 19616
rect 27674 19552 27690 19616
rect 27754 19552 27770 19616
rect 27834 19552 27850 19616
rect 27914 19552 27922 19616
rect 27602 18528 27922 19552
rect 27602 18464 27610 18528
rect 27674 18464 27690 18528
rect 27754 18464 27770 18528
rect 27834 18464 27850 18528
rect 27914 18464 27922 18528
rect 27602 17440 27922 18464
rect 27602 17376 27610 17440
rect 27674 17376 27690 17440
rect 27754 17376 27770 17440
rect 27834 17376 27850 17440
rect 27914 17376 27922 17440
rect 27602 16352 27922 17376
rect 27602 16288 27610 16352
rect 27674 16288 27690 16352
rect 27754 16288 27770 16352
rect 27834 16288 27850 16352
rect 27914 16288 27922 16352
rect 27602 15264 27922 16288
rect 27602 15200 27610 15264
rect 27674 15200 27690 15264
rect 27754 15200 27770 15264
rect 27834 15200 27850 15264
rect 27914 15200 27922 15264
rect 27602 14176 27922 15200
rect 27602 14112 27610 14176
rect 27674 14112 27690 14176
rect 27754 14112 27770 14176
rect 27834 14112 27850 14176
rect 27914 14112 27922 14176
rect 27602 13154 27922 14112
rect 27602 13088 27644 13154
rect 27880 13088 27922 13154
rect 27602 13024 27610 13088
rect 27914 13024 27922 13088
rect 27602 12918 27644 13024
rect 27880 12918 27922 13024
rect 27602 12000 27922 12918
rect 27602 11936 27610 12000
rect 27674 11936 27690 12000
rect 27754 11936 27770 12000
rect 27834 11936 27850 12000
rect 27914 11936 27922 12000
rect 27602 10912 27922 11936
rect 27602 10848 27610 10912
rect 27674 10848 27690 10912
rect 27754 10848 27770 10912
rect 27834 10848 27850 10912
rect 27914 10848 27922 10912
rect 27602 9824 27922 10848
rect 27602 9760 27610 9824
rect 27674 9760 27690 9824
rect 27754 9760 27770 9824
rect 27834 9760 27850 9824
rect 27914 9760 27922 9824
rect 27602 8736 27922 9760
rect 27602 8672 27610 8736
rect 27674 8672 27690 8736
rect 27754 8672 27770 8736
rect 27834 8672 27850 8736
rect 27914 8672 27922 8736
rect 27602 7648 27922 8672
rect 27602 7584 27610 7648
rect 27674 7584 27690 7648
rect 27754 7584 27770 7648
rect 27834 7584 27850 7648
rect 27914 7584 27922 7648
rect 27602 6560 27922 7584
rect 27602 6496 27610 6560
rect 27674 6496 27690 6560
rect 27754 6496 27770 6560
rect 27834 6496 27850 6560
rect 27914 6496 27922 6560
rect 27602 6354 27922 6496
rect 27602 6118 27644 6354
rect 27880 6118 27922 6354
rect 27602 5472 27922 6118
rect 27602 5408 27610 5472
rect 27674 5408 27690 5472
rect 27754 5408 27770 5472
rect 27834 5408 27850 5472
rect 27914 5408 27922 5472
rect 27602 4384 27922 5408
rect 27602 4320 27610 4384
rect 27674 4320 27690 4384
rect 27754 4320 27770 4384
rect 27834 4320 27850 4384
rect 27914 4320 27922 4384
rect 27602 3296 27922 4320
rect 27602 3232 27610 3296
rect 27674 3232 27690 3296
rect 27754 3232 27770 3296
rect 27834 3232 27850 3296
rect 27914 3232 27922 3296
rect 27602 2208 27922 3232
rect 27602 2144 27610 2208
rect 27674 2144 27690 2208
rect 27754 2144 27770 2208
rect 27834 2144 27850 2208
rect 27914 2144 27922 2208
rect 27602 2128 27922 2144
<< via4 >>
rect 4700 25858 4936 26094
rect 4700 19072 4936 19294
rect 4700 19058 4730 19072
rect 4730 19058 4746 19072
rect 4746 19058 4810 19072
rect 4810 19058 4826 19072
rect 4826 19058 4890 19072
rect 4890 19058 4906 19072
rect 4906 19058 4936 19072
rect 4700 12480 4730 12494
rect 4730 12480 4746 12494
rect 4746 12480 4810 12494
rect 4810 12480 4826 12494
rect 4826 12480 4890 12494
rect 4890 12480 4906 12494
rect 4906 12480 4936 12494
rect 4700 12258 4936 12480
rect 4700 5458 4936 5694
rect 5360 26518 5596 26754
rect 5360 19718 5596 19954
rect 5360 13088 5596 13154
rect 5360 13024 5390 13088
rect 5390 13024 5406 13088
rect 5406 13024 5470 13088
rect 5470 13024 5486 13088
rect 5486 13024 5550 13088
rect 5550 13024 5566 13088
rect 5566 13024 5596 13088
rect 5360 12918 5596 13024
rect 5360 6118 5596 6354
rect 12128 25858 12364 26094
rect 12128 19072 12364 19294
rect 12128 19058 12158 19072
rect 12158 19058 12174 19072
rect 12174 19058 12238 19072
rect 12238 19058 12254 19072
rect 12254 19058 12318 19072
rect 12318 19058 12334 19072
rect 12334 19058 12364 19072
rect 12128 12480 12158 12494
rect 12158 12480 12174 12494
rect 12174 12480 12238 12494
rect 12238 12480 12254 12494
rect 12254 12480 12318 12494
rect 12318 12480 12334 12494
rect 12334 12480 12364 12494
rect 12128 12258 12364 12480
rect 12128 5458 12364 5694
rect 12788 26518 13024 26754
rect 12788 19718 13024 19954
rect 12788 13088 13024 13154
rect 12788 13024 12818 13088
rect 12818 13024 12834 13088
rect 12834 13024 12898 13088
rect 12898 13024 12914 13088
rect 12914 13024 12978 13088
rect 12978 13024 12994 13088
rect 12994 13024 13024 13088
rect 12788 12918 13024 13024
rect 12788 6118 13024 6354
rect 19556 25858 19792 26094
rect 19556 19072 19792 19294
rect 19556 19058 19586 19072
rect 19586 19058 19602 19072
rect 19602 19058 19666 19072
rect 19666 19058 19682 19072
rect 19682 19058 19746 19072
rect 19746 19058 19762 19072
rect 19762 19058 19792 19072
rect 19556 12480 19586 12494
rect 19586 12480 19602 12494
rect 19602 12480 19666 12494
rect 19666 12480 19682 12494
rect 19682 12480 19746 12494
rect 19746 12480 19762 12494
rect 19762 12480 19792 12494
rect 19556 12258 19792 12480
rect 19556 5458 19792 5694
rect 20216 26518 20452 26754
rect 20216 19718 20452 19954
rect 20216 13088 20452 13154
rect 20216 13024 20246 13088
rect 20246 13024 20262 13088
rect 20262 13024 20326 13088
rect 20326 13024 20342 13088
rect 20342 13024 20406 13088
rect 20406 13024 20422 13088
rect 20422 13024 20452 13088
rect 20216 12918 20452 13024
rect 20216 6118 20452 6354
rect 26984 25858 27220 26094
rect 26984 19072 27220 19294
rect 26984 19058 27014 19072
rect 27014 19058 27030 19072
rect 27030 19058 27094 19072
rect 27094 19058 27110 19072
rect 27110 19058 27174 19072
rect 27174 19058 27190 19072
rect 27190 19058 27220 19072
rect 26984 12480 27014 12494
rect 27014 12480 27030 12494
rect 27030 12480 27094 12494
rect 27094 12480 27110 12494
rect 27110 12480 27174 12494
rect 27174 12480 27190 12494
rect 27190 12480 27220 12494
rect 26984 12258 27220 12480
rect 26984 5458 27220 5694
rect 27644 26518 27880 26754
rect 27644 19718 27880 19954
rect 27644 13088 27880 13154
rect 27644 13024 27674 13088
rect 27674 13024 27690 13088
rect 27690 13024 27754 13088
rect 27754 13024 27770 13088
rect 27770 13024 27834 13088
rect 27834 13024 27850 13088
rect 27850 13024 27880 13088
rect 27644 12918 27880 13024
rect 27644 6118 27880 6354
<< metal5 >>
rect 1056 26754 30868 26796
rect 1056 26518 5360 26754
rect 5596 26518 12788 26754
rect 13024 26518 20216 26754
rect 20452 26518 27644 26754
rect 27880 26518 30868 26754
rect 1056 26476 30868 26518
rect 1056 26094 30868 26136
rect 1056 25858 4700 26094
rect 4936 25858 12128 26094
rect 12364 25858 19556 26094
rect 19792 25858 26984 26094
rect 27220 25858 30868 26094
rect 1056 25816 30868 25858
rect 1056 19954 30868 19996
rect 1056 19718 5360 19954
rect 5596 19718 12788 19954
rect 13024 19718 20216 19954
rect 20452 19718 27644 19954
rect 27880 19718 30868 19954
rect 1056 19676 30868 19718
rect 1056 19294 30868 19336
rect 1056 19058 4700 19294
rect 4936 19058 12128 19294
rect 12364 19058 19556 19294
rect 19792 19058 26984 19294
rect 27220 19058 30868 19294
rect 1056 19016 30868 19058
rect 1056 13154 30868 13196
rect 1056 12918 5360 13154
rect 5596 12918 12788 13154
rect 13024 12918 20216 13154
rect 20452 12918 27644 13154
rect 27880 12918 30868 13154
rect 1056 12876 30868 12918
rect 1056 12494 30868 12536
rect 1056 12258 4700 12494
rect 4936 12258 12128 12494
rect 12364 12258 19556 12494
rect 19792 12258 26984 12494
rect 27220 12258 30868 12494
rect 1056 12216 30868 12258
rect 1056 6354 30868 6396
rect 1056 6118 5360 6354
rect 5596 6118 12788 6354
rect 13024 6118 20216 6354
rect 20452 6118 27644 6354
rect 27880 6118 30868 6354
rect 1056 6076 30868 6118
rect 1056 5694 30868 5736
rect 1056 5458 4700 5694
rect 4936 5458 12128 5694
rect 12364 5458 19556 5694
rect 19792 5458 26984 5694
rect 27220 5458 30868 5694
rect 1056 5416 30868 5458
use sky130_fd_sc_hd__clkbuf_4  _0588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0589_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13524 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0590_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0591_
timestamp 1694700623
transform 1 0 15364 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19044 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0593_
timestamp 1694700623
transform -1 0 18676 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 25116 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0595_
timestamp 1694700623
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9384 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0597_
timestamp 1694700623
transform 1 0 8280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0598_
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0599_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0600_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9108 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0601_
timestamp 1694700623
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0602_
timestamp 1694700623
transform 1 0 6440 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_2  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7636 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0604_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0605_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0606_
timestamp 1694700623
transform 1 0 5428 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0607_
timestamp 1694700623
transform 1 0 5428 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6992 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0609_
timestamp 1694700623
transform 1 0 6072 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0610_
timestamp 1694700623
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0611_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6900 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0612_
timestamp 1694700623
transform 1 0 10396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0613_
timestamp 1694700623
transform 1 0 11408 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0614_
timestamp 1694700623
transform 1 0 10488 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0616_
timestamp 1694700623
transform -1 0 6440 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0617_
timestamp 1694700623
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7084 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0620_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8096 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _0621_
timestamp 1694700623
transform 1 0 6532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0622_
timestamp 1694700623
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0623_
timestamp 1694700623
transform 1 0 6624 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9108 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1694700623
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0626_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8004 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_4  _0627_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7268 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_1  _0628_
timestamp 1694700623
transform 1 0 13248 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 1694700623
transform 1 0 13800 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0630_
timestamp 1694700623
transform -1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0631_
timestamp 1694700623
transform -1 0 14720 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1694700623
transform 1 0 14168 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0633_
timestamp 1694700623
transform -1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0634_
timestamp 1694700623
transform -1 0 16376 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0635_
timestamp 1694700623
transform -1 0 15640 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0636_
timestamp 1694700623
transform -1 0 14904 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0637_
timestamp 1694700623
transform -1 0 15456 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0638_
timestamp 1694700623
transform 1 0 12052 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0639_
timestamp 1694700623
transform -1 0 13432 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0640_
timestamp 1694700623
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0641_
timestamp 1694700623
transform 1 0 6624 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0642_
timestamp 1694700623
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0643_
timestamp 1694700623
transform 1 0 9016 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0644_
timestamp 1694700623
transform 1 0 9016 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0645_
timestamp 1694700623
transform -1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0646_
timestamp 1694700623
transform -1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0647_
timestamp 1694700623
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0648_
timestamp 1694700623
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0649_
timestamp 1694700623
transform -1 0 14352 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0650_
timestamp 1694700623
transform 1 0 14260 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0651_
timestamp 1694700623
transform 1 0 14076 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1694700623
transform -1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0654_
timestamp 1694700623
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13984 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0657_
timestamp 1694700623
transform 1 0 13156 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0658_
timestamp 1694700623
transform -1 0 13892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_2  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _0661_
timestamp 1694700623
transform -1 0 22080 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1694700623
transform -1 0 25852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1694700623
transform 1 0 26312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0664_
timestamp 1694700623
transform 1 0 24564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0665_
timestamp 1694700623
transform 1 0 23460 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1694700623
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0667_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 24932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1694700623
transform 1 0 25392 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0669_
timestamp 1694700623
transform 1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0670_
timestamp 1694700623
transform 1 0 24840 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0671_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0672_
timestamp 1694700623
transform -1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0673_
timestamp 1694700623
transform -1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0674_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14076 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0675_
timestamp 1694700623
transform 1 0 16928 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0676_
timestamp 1694700623
transform 1 0 16836 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0677_
timestamp 1694700623
transform -1 0 17848 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0678_
timestamp 1694700623
transform -1 0 21344 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0679_
timestamp 1694700623
transform 1 0 22540 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22908 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 18400 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0682_
timestamp 1694700623
transform 1 0 18676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0683_
timestamp 1694700623
transform 1 0 10672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 24288 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_2  _0685_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19872 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0686_
timestamp 1694700623
transform 1 0 13984 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 23736 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0688_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 23736 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0689_
timestamp 1694700623
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1694700623
transform 1 0 25852 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0691_
timestamp 1694700623
transform -1 0 26312 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0692_
timestamp 1694700623
transform 1 0 18124 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0693_
timestamp 1694700623
transform -1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 1694700623
transform 1 0 22632 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 1694700623
transform -1 0 21620 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0696_
timestamp 1694700623
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0697_
timestamp 1694700623
transform 1 0 19504 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0698_
timestamp 1694700623
transform -1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0699_
timestamp 1694700623
transform 1 0 20148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0700_
timestamp 1694700623
transform 1 0 19412 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0701_
timestamp 1694700623
transform -1 0 17848 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0702_
timestamp 1694700623
transform -1 0 17572 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1694700623
transform 1 0 14536 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0704_
timestamp 1694700623
transform -1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0705_
timestamp 1694700623
transform 1 0 12604 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1694700623
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15364 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0708_
timestamp 1694700623
transform -1 0 15640 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1694700623
transform 1 0 14628 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0710_
timestamp 1694700623
transform -1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 1694700623
transform 1 0 12144 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 1694700623
transform -1 0 11408 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0713_
timestamp 1694700623
transform -1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0714_
timestamp 1694700623
transform 1 0 14904 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0715_
timestamp 1694700623
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1694700623
transform 1 0 12972 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0717_
timestamp 1694700623
transform 1 0 11592 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0718_
timestamp 1694700623
transform -1 0 17940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0719_
timestamp 1694700623
transform -1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0720_
timestamp 1694700623
transform 1 0 15364 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0721_
timestamp 1694700623
transform 1 0 17572 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0722_
timestamp 1694700623
transform 1 0 16928 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1694700623
transform -1 0 17296 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0724_
timestamp 1694700623
transform -1 0 17572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1694700623
transform -1 0 14076 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 1694700623
transform 1 0 15364 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0727_
timestamp 1694700623
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0728_
timestamp 1694700623
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 1694700623
transform 1 0 12696 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0730_
timestamp 1694700623
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0731_
timestamp 1694700623
transform 1 0 14904 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0732_
timestamp 1694700623
transform -1 0 15456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0733_
timestamp 1694700623
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 1694700623
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0735_
timestamp 1694700623
transform 1 0 13800 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1694700623
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _0737_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10488 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _0738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0739_
timestamp 1694700623
transform 1 0 14628 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0740_
timestamp 1694700623
transform -1 0 15640 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0741_
timestamp 1694700623
transform -1 0 16468 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0742_
timestamp 1694700623
transform -1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1694700623
transform 1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0744_
timestamp 1694700623
transform 1 0 12328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0745_
timestamp 1694700623
transform 1 0 12880 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _0746_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1694700623
transform 1 0 11500 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0748_
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1694700623
transform 1 0 9384 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0750_
timestamp 1694700623
transform -1 0 9384 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 1694700623
transform -1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0752_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 1694700623
transform -1 0 10672 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0754_
timestamp 1694700623
transform 1 0 8280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1694700623
transform 1 0 6992 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0756_
timestamp 1694700623
transform 1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1694700623
transform -1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_4  _0758_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15088 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _0759_
timestamp 1694700623
transform 1 0 10212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0760_
timestamp 1694700623
transform 1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0761_
timestamp 1694700623
transform 1 0 7912 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1694700623
transform 1 0 4324 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0763_
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0764_
timestamp 1694700623
transform -1 0 9752 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1694700623
transform 1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0766_
timestamp 1694700623
transform -1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0767_
timestamp 1694700623
transform -1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1694700623
transform 1 0 10028 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1694700623
transform 1 0 10580 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0770_
timestamp 1694700623
transform 1 0 9752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1694700623
transform 1 0 4140 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0772_
timestamp 1694700623
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0773_
timestamp 1694700623
transform 1 0 9752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1694700623
transform 1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0775_
timestamp 1694700623
transform -1 0 10304 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1694700623
transform -1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0777_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9752 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0778_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10396 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1694700623
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0780_
timestamp 1694700623
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1694700623
transform -1 0 9568 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1694700623
transform 1 0 7544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0783_
timestamp 1694700623
transform 1 0 7820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0784_
timestamp 1694700623
transform -1 0 8096 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0785_
timestamp 1694700623
transform 1 0 7728 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0786_
timestamp 1694700623
transform -1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1694700623
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0788_
timestamp 1694700623
transform 1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0789_
timestamp 1694700623
transform 1 0 8096 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1694700623
transform 1 0 9108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0791_
timestamp 1694700623
transform -1 0 9844 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0792_
timestamp 1694700623
transform 1 0 8280 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1694700623
transform 1 0 3128 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0794_
timestamp 1694700623
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0795_
timestamp 1694700623
transform 1 0 8924 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1694700623
transform -1 0 9384 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1694700623
transform -1 0 8740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0798_
timestamp 1694700623
transform -1 0 7084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 1694700623
transform 1 0 6808 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0800_
timestamp 1694700623
transform 1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0802_
timestamp 1694700623
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1694700623
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0804_
timestamp 1694700623
transform 1 0 6900 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0805_
timestamp 1694700623
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1694700623
transform 1 0 4692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 1694700623
transform 1 0 4140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0808_
timestamp 1694700623
transform -1 0 10396 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0809_
timestamp 1694700623
transform 1 0 10948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0810_
timestamp 1694700623
transform -1 0 12144 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0811_
timestamp 1694700623
transform 1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1694700623
transform 1 0 9200 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 1694700623
transform -1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0814_
timestamp 1694700623
transform -1 0 13524 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0815_
timestamp 1694700623
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0816_
timestamp 1694700623
transform 1 0 11684 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0817_
timestamp 1694700623
transform -1 0 13616 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1694700623
transform -1 0 12696 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0819_
timestamp 1694700623
transform -1 0 15732 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1694700623
transform -1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0821_
timestamp 1694700623
transform -1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0822_
timestamp 1694700623
transform 1 0 12512 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1694700623
transform 1 0 6440 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0825_
timestamp 1694700623
transform -1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0826_
timestamp 1694700623
transform 1 0 10488 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1694700623
transform -1 0 12512 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1694700623
transform -1 0 11868 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0829_
timestamp 1694700623
transform -1 0 9476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1694700623
transform -1 0 7912 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1694700623
transform 1 0 6716 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0832_
timestamp 1694700623
transform 1 0 5244 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0833_
timestamp 1694700623
transform 1 0 4140 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0834_
timestamp 1694700623
transform 1 0 3864 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1694700623
transform -1 0 5704 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0836_
timestamp 1694700623
transform -1 0 4968 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0837_
timestamp 1694700623
transform 1 0 18032 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0838_
timestamp 1694700623
transform -1 0 12696 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0839_
timestamp 1694700623
transform -1 0 5244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0840_
timestamp 1694700623
transform -1 0 13248 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1694700623
transform 1 0 6992 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0842_
timestamp 1694700623
transform 1 0 7728 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0843_
timestamp 1694700623
transform -1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0844_
timestamp 1694700623
transform 1 0 9476 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0845_
timestamp 1694700623
transform -1 0 10028 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0846_
timestamp 1694700623
transform -1 0 9568 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1694700623
transform -1 0 8648 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0848_
timestamp 1694700623
transform 1 0 7452 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0849_
timestamp 1694700623
transform -1 0 12604 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1694700623
transform 1 0 9568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0852_
timestamp 1694700623
transform -1 0 6256 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7728 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7176 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1694700623
transform 1 0 4600 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1694700623
transform 1 0 5244 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0857_
timestamp 1694700623
transform 1 0 6348 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0858_
timestamp 1694700623
transform 1 0 6348 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0859_
timestamp 1694700623
transform -1 0 8280 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0860_
timestamp 1694700623
transform -1 0 6992 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0861_
timestamp 1694700623
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0862_
timestamp 1694700623
transform 1 0 6900 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1694700623
transform 1 0 7360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0864_
timestamp 1694700623
transform 1 0 7268 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0865_
timestamp 1694700623
transform -1 0 9936 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0866_
timestamp 1694700623
transform -1 0 8648 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0867_
timestamp 1694700623
transform 1 0 8372 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1694700623
transform 1 0 8924 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0869_
timestamp 1694700623
transform -1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0870_
timestamp 1694700623
transform -1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1694700623
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0872_
timestamp 1694700623
transform -1 0 11776 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0873_
timestamp 1694700623
transform 1 0 10672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1694700623
transform -1 0 10856 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0875_
timestamp 1694700623
transform 1 0 10396 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1694700623
transform 1 0 10396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0877_
timestamp 1694700623
transform 1 0 10120 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1694700623
transform -1 0 12052 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1694700623
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0880_
timestamp 1694700623
transform 1 0 10764 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1694700623
transform 1 0 9936 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0882_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14904 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1694700623
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0884_
timestamp 1694700623
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0885_
timestamp 1694700623
transform -1 0 13892 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1694700623
transform -1 0 13984 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 1694700623
transform -1 0 14904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 1694700623
transform 1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1694700623
transform -1 0 16008 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1694700623
transform -1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 1694700623
transform 1 0 4324 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1694700623
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 1694700623
transform 1 0 3864 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1694700623
transform 1 0 3128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1694700623
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1694700623
transform 1 0 5520 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 1694700623
transform 1 0 9384 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1694700623
transform 1 0 8188 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0900_
timestamp 1694700623
transform 1 0 12328 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1694700623
transform -1 0 12144 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0902_
timestamp 1694700623
transform -1 0 19780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0903_
timestamp 1694700623
transform -1 0 22724 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0904_
timestamp 1694700623
transform 1 0 28704 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0905_
timestamp 1694700623
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1694700623
transform -1 0 29440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0907_
timestamp 1694700623
transform 1 0 22264 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0908_
timestamp 1694700623
transform 1 0 22816 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0909_
timestamp 1694700623
transform 1 0 24656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0910_
timestamp 1694700623
transform 1 0 22724 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1694700623
transform -1 0 25668 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0912_
timestamp 1694700623
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0913_
timestamp 1694700623
transform 1 0 25116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0914_
timestamp 1694700623
transform -1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0915_
timestamp 1694700623
transform 1 0 27232 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0916_
timestamp 1694700623
transform 1 0 27784 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0917_
timestamp 1694700623
transform -1 0 27968 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0918_
timestamp 1694700623
transform 1 0 26128 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0919_
timestamp 1694700623
transform 1 0 23644 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1694700623
transform -1 0 25668 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 25668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0922_
timestamp 1694700623
transform 1 0 23368 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1694700623
transform 1 0 24196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0924_
timestamp 1694700623
transform 1 0 24104 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0925_
timestamp 1694700623
transform -1 0 24656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0926_
timestamp 1694700623
transform 1 0 24472 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1694700623
transform 1 0 25484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0928_
timestamp 1694700623
transform -1 0 25852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0929_
timestamp 1694700623
transform 1 0 26772 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0930_
timestamp 1694700623
transform -1 0 26864 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0931_
timestamp 1694700623
transform 1 0 28244 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0932_
timestamp 1694700623
transform 1 0 27692 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0933_
timestamp 1694700623
transform 1 0 29808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0934_
timestamp 1694700623
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0935_
timestamp 1694700623
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0936_
timestamp 1694700623
transform 1 0 28704 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0937_
timestamp 1694700623
transform 1 0 27600 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0938_
timestamp 1694700623
transform 1 0 27600 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0939_
timestamp 1694700623
transform -1 0 29440 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1694700623
transform -1 0 29348 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0941_
timestamp 1694700623
transform -1 0 29440 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0942_
timestamp 1694700623
transform 1 0 29256 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0943_
timestamp 1694700623
transform -1 0 28704 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0944_
timestamp 1694700623
transform 1 0 28152 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0945_
timestamp 1694700623
transform 1 0 21896 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0946_
timestamp 1694700623
transform 1 0 22448 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 23552 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0948_
timestamp 1694700623
transform -1 0 19504 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0949_
timestamp 1694700623
transform -1 0 19780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0950_
timestamp 1694700623
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1694700623
transform 1 0 19044 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1694700623
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp 1694700623
transform 1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0955_
timestamp 1694700623
transform 1 0 16008 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0956_
timestamp 1694700623
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16928 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0958_
timestamp 1694700623
transform -1 0 22356 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0959_
timestamp 1694700623
transform 1 0 19228 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0960_
timestamp 1694700623
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0961_
timestamp 1694700623
transform -1 0 27876 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0962_
timestamp 1694700623
transform -1 0 27416 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0963_
timestamp 1694700623
transform -1 0 21620 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0964_
timestamp 1694700623
transform -1 0 19044 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0965_
timestamp 1694700623
transform 1 0 15732 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0966_
timestamp 1694700623
transform -1 0 17480 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0967_
timestamp 1694700623
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0968_
timestamp 1694700623
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 1694700623
transform 1 0 16192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1694700623
transform 1 0 18584 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0971_
timestamp 1694700623
transform -1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0972_
timestamp 1694700623
transform -1 0 19228 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1694700623
transform 1 0 19228 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0974_
timestamp 1694700623
transform 1 0 17848 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0975_
timestamp 1694700623
transform 1 0 17204 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1694700623
transform 1 0 16744 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1694700623
transform -1 0 21436 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0978_
timestamp 1694700623
transform -1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0979_
timestamp 1694700623
transform 1 0 19504 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0981_
timestamp 1694700623
transform -1 0 20608 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0982_
timestamp 1694700623
transform -1 0 19136 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0983_
timestamp 1694700623
transform 1 0 17480 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0984_
timestamp 1694700623
transform 1 0 17204 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1694700623
transform 1 0 16928 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0986_
timestamp 1694700623
transform -1 0 23000 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1694700623
transform -1 0 24012 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1694700623
transform -1 0 23184 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0989_
timestamp 1694700623
transform 1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1694700623
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1694700623
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1694700623
transform 1 0 27416 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1694700623
transform -1 0 26956 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1694700623
transform 1 0 28888 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0995_
timestamp 1694700623
transform 1 0 28520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0996_
timestamp 1694700623
transform 1 0 28612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0997_
timestamp 1694700623
transform -1 0 30176 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0998_
timestamp 1694700623
transform 1 0 25944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1694700623
transform 1 0 23552 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1694700623
transform 1 0 23000 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 29348 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1002_
timestamp 1694700623
transform 1 0 26772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1003_
timestamp 1694700623
transform 1 0 27048 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1004_
timestamp 1694700623
transform -1 0 28152 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1694700623
transform 1 0 25116 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1694700623
transform 1 0 24932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1007_
timestamp 1694700623
transform 1 0 28244 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1694700623
transform -1 0 27968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1009_
timestamp 1694700623
transform 1 0 27416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1010_
timestamp 1694700623
transform -1 0 30360 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1011_
timestamp 1694700623
transform -1 0 30084 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1012_
timestamp 1694700623
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 1694700623
transform 1 0 24748 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1694700623
transform 1 0 24472 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1694700623
transform 1 0 28520 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1016_
timestamp 1694700623
transform 1 0 27968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 1694700623
transform 1 0 28060 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1018_
timestamp 1694700623
transform 1 0 27784 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1694700623
transform 1 0 25760 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1694700623
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1694700623
transform 1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1022_
timestamp 1694700623
transform 1 0 24472 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1694700623
transform -1 0 24472 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1024_
timestamp 1694700623
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1025_
timestamp 1694700623
transform -1 0 25944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1026_
timestamp 1694700623
transform -1 0 26588 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1027_
timestamp 1694700623
transform -1 0 28336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1028_
timestamp 1694700623
transform 1 0 27140 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1029_
timestamp 1694700623
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp 1694700623
transform 1 0 25576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1694700623
transform 1 0 25024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1032_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22908 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1033_
timestamp 1694700623
transform -1 0 24012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1034_
timestamp 1694700623
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1035_
timestamp 1694700623
transform 1 0 22264 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1694700623
transform 1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1037_
timestamp 1694700623
transform 1 0 23092 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1038_
timestamp 1694700623
transform -1 0 24196 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp 1694700623
transform 1 0 23460 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1694700623
transform -1 0 23276 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1041_
timestamp 1694700623
transform 1 0 21344 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1042_
timestamp 1694700623
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1043_
timestamp 1694700623
transform -1 0 25208 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1044_
timestamp 1694700623
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1045_
timestamp 1694700623
transform 1 0 19688 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1694700623
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1047_
timestamp 1694700623
transform -1 0 25484 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1048_
timestamp 1694700623
transform -1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1049_
timestamp 1694700623
transform 1 0 21252 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1050_
timestamp 1694700623
transform -1 0 22724 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1694700623
transform 1 0 21252 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1694700623
transform 1 0 20056 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 22908 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1054_
timestamp 1694700623
transform 1 0 24472 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1055_
timestamp 1694700623
transform -1 0 25852 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1056_
timestamp 1694700623
transform 1 0 21988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1057_
timestamp 1694700623
transform -1 0 21712 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1694700623
transform -1 0 21988 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1059_
timestamp 1694700623
transform 1 0 14628 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1060_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15272 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_4  _1061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11868 0 1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1694700623
transform -1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1064_
timestamp 1694700623
transform -1 0 11868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1065_
timestamp 1694700623
transform -1 0 12328 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1066_
timestamp 1694700623
transform -1 0 12880 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1068_
timestamp 1694700623
transform -1 0 6992 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1069_
timestamp 1694700623
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1070_
timestamp 1694700623
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1071_
timestamp 1694700623
transform -1 0 5428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1072_
timestamp 1694700623
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1073_
timestamp 1694700623
transform -1 0 6256 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1074_
timestamp 1694700623
transform -1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1075_
timestamp 1694700623
transform -1 0 8004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1076_
timestamp 1694700623
transform -1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1077_
timestamp 1694700623
transform -1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1078_
timestamp 1694700623
transform -1 0 19780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1079_
timestamp 1694700623
transform 1 0 19780 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1080_
timestamp 1694700623
transform -1 0 19136 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _1081_
timestamp 1694700623
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1082_
timestamp 1694700623
transform 1 0 17664 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1083_
timestamp 1694700623
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1084_
timestamp 1694700623
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1085_
timestamp 1694700623
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1086_
timestamp 1694700623
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1087_
timestamp 1694700623
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1088_
timestamp 1694700623
transform 1 0 19044 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1089_
timestamp 1694700623
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1090_
timestamp 1694700623
transform 1 0 18584 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _1091_
timestamp 1694700623
transform 1 0 19228 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1092_
timestamp 1694700623
transform 1 0 19688 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1093_
timestamp 1694700623
transform 1 0 20148 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1094_
timestamp 1694700623
transform 1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand4b_2  _1095_
timestamp 1694700623
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1096_
timestamp 1694700623
transform -1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1097_
timestamp 1694700623
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1098_
timestamp 1694700623
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1099_
timestamp 1694700623
transform 1 0 22540 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1100_
timestamp 1694700623
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1101_
timestamp 1694700623
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1102_
timestamp 1694700623
transform -1 0 21712 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1103_
timestamp 1694700623
transform 1 0 19872 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1104_
timestamp 1694700623
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4b_2  _1105_
timestamp 1694700623
transform -1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1106_
timestamp 1694700623
transform 1 0 14812 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1107_
timestamp 1694700623
transform 1 0 15272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1108_
timestamp 1694700623
transform 1 0 14076 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1694700623
transform -1 0 14536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1694700623
transform -1 0 15640 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1694700623
transform 1 0 15272 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1694700623
transform 1 0 14904 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1113_
timestamp 1694700623
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1114_
timestamp 1694700623
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1115_
timestamp 1694700623
transform 1 0 16376 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1118_
timestamp 1694700623
transform -1 0 13340 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1119_
timestamp 1694700623
transform 1 0 12512 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1120_
timestamp 1694700623
transform -1 0 9568 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1121_
timestamp 1694700623
transform -1 0 8188 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1122_
timestamp 1694700623
transform -1 0 5336 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1123_
timestamp 1694700623
transform -1 0 5796 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1124_
timestamp 1694700623
transform 1 0 10580 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1125_
timestamp 1694700623
transform 1 0 23184 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1694700623
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1694700623
transform -1 0 21712 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1694700623
transform -1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1694700623
transform 1 0 23828 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1694700623
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1694700623
transform 1 0 24748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1694700623
transform 1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1694700623
transform 1 0 25300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1694700623
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1694700623
transform -1 0 22448 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1136_
timestamp 1694700623
transform -1 0 11408 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1694700623
transform 1 0 18032 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1694700623
transform 1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1694700623
transform 1 0 16652 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1694700623
transform -1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1694700623
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1694700623
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1694700623
transform -1 0 3680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1694700623
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1694700623
transform 1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1694700623
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1147_
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1694700623
transform 1 0 14536 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1149_
timestamp 1694700623
transform -1 0 19780 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1150_
timestamp 1694700623
transform 1 0 17480 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1694700623
transform -1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1694700623
transform 1 0 15456 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1694700623
transform -1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1694700623
transform 1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1155_
timestamp 1694700623
transform -1 0 18032 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1694700623
transform -1 0 17204 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1694700623
transform -1 0 12972 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1158_
timestamp 1694700623
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1159_
timestamp 1694700623
transform 1 0 14536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1160_
timestamp 1694700623
transform -1 0 15732 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1161_
timestamp 1694700623
transform 1 0 15272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1694700623
transform -1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1694700623
transform -1 0 11960 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1694700623
transform 1 0 9292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1694700623
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1694700623
transform -1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1167_
timestamp 1694700623
transform -1 0 11408 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1694700623
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1694700623
transform 1 0 11040 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1694700623
transform 1 0 4416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1694700623
transform -1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1694700623
transform -1 0 3220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1694700623
transform -1 0 3404 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1694700623
transform -1 0 3404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1694700623
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1694700623
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1177_
timestamp 1694700623
transform 1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1694700623
transform -1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1694700623
transform -1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1694700623
transform -1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1694700623
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1694700623
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1694700623
transform 1 0 20148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1694700623
transform 1 0 22356 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1694700623
transform 1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21988 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19596 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1189_
timestamp 1694700623
transform 1 0 19228 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1694700623
transform 1 0 23736 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1694700623
transform 1 0 24472 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1694700623
transform 1 0 23920 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1694700623
transform 1 0 24012 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1694700623
transform 1 0 24472 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1694700623
transform 1 0 22448 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1694700623
transform 1 0 20332 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1197_
timestamp 1694700623
transform 1 0 16652 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1198_
timestamp 1694700623
transform 1 0 16192 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15640 0 1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1200_
timestamp 1694700623
transform 1 0 12144 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1201_
timestamp 1694700623
transform 1 0 7544 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1202_
timestamp 1694700623
transform 1 0 5060 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1203_
timestamp 1694700623
transform 1 0 2668 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1204_
timestamp 1694700623
transform 1 0 2484 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1205_
timestamp 1694700623
transform 1 0 16008 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1206_
timestamp 1694700623
transform 1 0 14076 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1207_
timestamp 1694700623
transform 1 0 13524 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 20700 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1694700623
transform 1 0 12788 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1694700623
transform 1 0 14536 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1211_
timestamp 1694700623
transform 1 0 14444 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1694700623
transform 1 0 13892 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1213_
timestamp 1694700623
transform 1 0 16652 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1214_
timestamp 1694700623
transform 1 0 17204 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1215_
timestamp 1694700623
transform 1 0 11592 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1216_
timestamp 1694700623
transform -1 0 14536 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1217_
timestamp 1694700623
transform 1 0 14812 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1218_
timestamp 1694700623
transform 1 0 16652 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_2  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12328 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1220_
timestamp 1694700623
transform -1 0 10948 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1222_
timestamp 1694700623
transform 1 0 4140 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1223_
timestamp 1694700623
transform -1 0 5796 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1224_
timestamp 1694700623
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1225_
timestamp 1694700623
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1226_
timestamp 1694700623
transform 1 0 6440 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1227_
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1228_
timestamp 1694700623
transform -1 0 10488 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1229_
timestamp 1694700623
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1230_
timestamp 1694700623
transform -1 0 18400 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1231_
timestamp 1694700623
transform -1 0 18308 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1232_
timestamp 1694700623
transform -1 0 19136 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1233_
timestamp 1694700623
transform -1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1234_
timestamp 1694700623
transform -1 0 15732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1235_
timestamp 1694700623
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1236_
timestamp 1694700623
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1237_
timestamp 1694700623
transform 1 0 22356 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1238_
timestamp 1694700623
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1239_
timestamp 1694700623
transform 1 0 19780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1240_
timestamp 1694700623
transform 1 0 20608 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1241_
timestamp 1694700623
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1242_
timestamp 1694700623
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1243_
timestamp 1694700623
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1244_
timestamp 1694700623
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1245_
timestamp 1694700623
transform 1 0 25576 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1246_
timestamp 1694700623
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1247_
timestamp 1694700623
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1248_
timestamp 1694700623
transform -1 0 21160 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1249_
timestamp 1694700623
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1250_
timestamp 1694700623
transform 1 0 14628 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1251_
timestamp 1694700623
transform -1 0 18492 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1252_
timestamp 1694700623
transform 1 0 18308 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1694700623
transform 1 0 10396 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 1694700623
transform 1 0 10580 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1255_
timestamp 1694700623
transform -1 0 10396 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1256_
timestamp 1694700623
transform -1 0 6532 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1257_
timestamp 1694700623
transform 1 0 6348 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1258_
timestamp 1694700623
transform 1 0 10488 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 1694700623
transform 1 0 9200 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1694700623
transform 1 0 3772 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1694700623
transform 1 0 2024 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1694700623
transform 1 0 1840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 1694700623
transform 1 0 1840 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1264_
timestamp 1694700623
transform 1 0 1748 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1694700623
transform 1 0 2300 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1266_
timestamp 1694700623
transform 1 0 3404 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 1694700623
transform 1 0 5704 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1694700623
transform 1 0 10488 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1269_
timestamp 1694700623
transform 1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1270_
timestamp 1694700623
transform 1 0 15364 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1271_
timestamp 1694700623
transform 1 0 17296 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 1694700623
transform 1 0 11132 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1274_
timestamp 1694700623
transform 1 0 19136 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1275_
timestamp 1694700623
transform 1 0 21804 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1276_
timestamp 1694700623
transform 1 0 23644 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  _1277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12052 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1278_
timestamp 1694700623
transform 1 0 9476 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1279_
timestamp 1694700623
transform 1 0 6532 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1280_
timestamp 1694700623
transform -1 0 5888 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1281_
timestamp 1694700623
transform 1 0 4324 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1282_
timestamp 1694700623
transform 1 0 4692 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1283_
timestamp 1694700623
transform 1 0 4692 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1284_
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1285_
timestamp 1694700623
transform 1 0 5152 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1286_
timestamp 1694700623
transform 1 0 7452 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1287_
timestamp 1694700623
transform -1 0 13524 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1288_
timestamp 1694700623
transform 1 0 17204 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1289_
timestamp 1694700623
transform 1 0 17112 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1290_
timestamp 1694700623
transform 1 0 18124 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1291_
timestamp 1694700623
transform 1 0 16652 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1292_
timestamp 1694700623
transform 1 0 14168 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1293_
timestamp 1694700623
transform 1 0 19688 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1294_
timestamp 1694700623
transform -1 0 22632 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1295_
timestamp 1694700623
transform -1 0 24012 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1296_
timestamp 1694700623
transform 1 0 19964 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1297_
timestamp 1694700623
transform 1 0 19320 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1298_
timestamp 1694700623
transform 1 0 20424 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1299_
timestamp 1694700623
transform -1 0 23736 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1300_
timestamp 1694700623
transform 1 0 26312 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1301_
timestamp 1694700623
transform 1 0 25576 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1302_
timestamp 1694700623
transform 1 0 25576 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1303_
timestamp 1694700623
transform 1 0 24840 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1304_
timestamp 1694700623
transform 1 0 23644 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1305_
timestamp 1694700623
transform 1 0 20976 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1306_
timestamp 1694700623
transform 1 0 19780 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1307_
timestamp 1694700623
transform 1 0 19228 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1308_
timestamp 1694700623
transform 1 0 14260 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12236 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clock
timestamp 1694700623
transform -1 0 8464 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clock
timestamp 1694700623
transform -1 0 9476 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clock
timestamp 1694700623
transform 1 0 18584 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clock
timestamp 1694700623
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1694700623
transform -1 0 13248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1694700623
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout12
timestamp 1694700623
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1694700623
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1694700623
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1694700623
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1694700623
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1694700623
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1694700623
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1694700623
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1694700623
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1694700623
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1694700623
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1694700623
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1694700623
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1694700623
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1694700623
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1694700623
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1694700623
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1694700623
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1694700623
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1694700623
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1694700623
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1694700623
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1694700623
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1694700623
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1694700623
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1694700623
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1694700623
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1694700623
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1694700623
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_317
timestamp 1694700623
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1694700623
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1694700623
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1694700623
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1694700623
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1694700623
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1694700623
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1694700623
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1694700623
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1694700623
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1694700623
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1694700623
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1694700623
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1694700623
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1694700623
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1694700623
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1694700623
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1694700623
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1694700623
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1694700623
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1694700623
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1694700623
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1694700623
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1694700623
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1694700623
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1694700623
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1694700623
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1694700623
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1694700623
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_317
timestamp 1694700623
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1694700623
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1694700623
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1694700623
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1694700623
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1694700623
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1694700623
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1694700623
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1694700623
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1694700623
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1694700623
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1694700623
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1694700623
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1694700623
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1694700623
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1694700623
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1694700623
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1694700623
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1694700623
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1694700623
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1694700623
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1694700623
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1694700623
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1694700623
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1694700623
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1694700623
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1694700623
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1694700623
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1694700623
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1694700623
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_309
timestamp 1694700623
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_317
timestamp 1694700623
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1694700623
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1694700623
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1694700623
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1694700623
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1694700623
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1694700623
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1694700623
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1694700623
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1694700623
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1694700623
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1694700623
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1694700623
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1694700623
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1694700623
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1694700623
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1694700623
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1694700623
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1694700623
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1694700623
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1694700623
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1694700623
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1694700623
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1694700623
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1694700623
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1694700623
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1694700623
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1694700623
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1694700623
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1694700623
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1694700623
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_317
timestamp 1694700623
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1694700623
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1694700623
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1694700623
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1694700623
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1694700623
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1694700623
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1694700623
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1694700623
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1694700623
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1694700623
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1694700623
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1694700623
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1694700623
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1694700623
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1694700623
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1694700623
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1694700623
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1694700623
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1694700623
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1694700623
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1694700623
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1694700623
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1694700623
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1694700623
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1694700623
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1694700623
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1694700623
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1694700623
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_309
timestamp 1694700623
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_317
timestamp 1694700623
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1694700623
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1694700623
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1694700623
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1694700623
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1694700623
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1694700623
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1694700623
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1694700623
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1694700623
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_116
timestamp 1694700623
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_126
timestamp 1694700623
transform 1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_134
timestamp 1694700623
transform 1 0 13432 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_144
timestamp 1694700623
transform 1 0 14352 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_154
timestamp 1694700623
transform 1 0 15272 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1694700623
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1694700623
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1694700623
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1694700623
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1694700623
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1694700623
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1694700623
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1694700623
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1694700623
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1694700623
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1694700623
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1694700623
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1694700623
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1694700623
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1694700623
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_317
timestamp 1694700623
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1694700623
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1694700623
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_49
timestamp 1694700623
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_70
timestamp 1694700623
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1694700623
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_92
timestamp 1694700623
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_100
timestamp 1694700623
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_129
timestamp 1694700623
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1694700623
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_156
timestamp 1694700623
transform 1 0 15456 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1694700623
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1694700623
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_197
timestamp 1694700623
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_202
timestamp 1694700623
transform 1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_206
timestamp 1694700623
transform 1 0 20056 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_210
timestamp 1694700623
transform 1 0 20424 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_222
timestamp 1694700623
transform 1 0 21528 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_230
timestamp 1694700623
transform 1 0 22264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_234
timestamp 1694700623
transform 1 0 22632 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_242
timestamp 1694700623
transform 1 0 23368 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_246
timestamp 1694700623
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1694700623
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1694700623
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1694700623
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1694700623
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1694700623
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1694700623
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_309
timestamp 1694700623
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_317
timestamp 1694700623
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1694700623
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1694700623
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1694700623
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_116
timestamp 1694700623
transform 1 0 11776 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_128
timestamp 1694700623
transform 1 0 12880 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_140
timestamp 1694700623
transform 1 0 13984 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_152
timestamp 1694700623
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_159
timestamp 1694700623
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1694700623
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_169
timestamp 1694700623
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_175
timestamp 1694700623
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_188
timestamp 1694700623
transform 1 0 18400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_217
timestamp 1694700623
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1694700623
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_265
timestamp 1694700623
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1694700623
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1694700623
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1694700623
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1694700623
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_317
timestamp 1694700623
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1694700623
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1694700623
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_53
timestamp 1694700623
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_59
timestamp 1694700623
transform 1 0 6532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_63
timestamp 1694700623
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_73
timestamp 1694700623
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1694700623
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_92
timestamp 1694700623
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_104
timestamp 1694700623
transform 1 0 10672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_112
timestamp 1694700623
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_122
timestamp 1694700623
transform 1 0 12328 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_128
timestamp 1694700623
transform 1 0 12880 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_167
timestamp 1694700623
transform 1 0 16468 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_209
timestamp 1694700623
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_246
timestamp 1694700623
transform 1 0 23736 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1694700623
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1694700623
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1694700623
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1694700623
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1694700623
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1694700623
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_309
timestamp 1694700623
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_317
timestamp 1694700623
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1694700623
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_23
timestamp 1694700623
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1694700623
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1694700623
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1694700623
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_77
timestamp 1694700623
transform 1 0 8188 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_86
timestamp 1694700623
transform 1 0 9016 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_98
timestamp 1694700623
transform 1 0 10120 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1694700623
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_148
timestamp 1694700623
transform 1 0 14720 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_154
timestamp 1694700623
transform 1 0 15272 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_163
timestamp 1694700623
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1694700623
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1694700623
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_177
timestamp 1694700623
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_190
timestamp 1694700623
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_194
timestamp 1694700623
transform 1 0 18952 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_216
timestamp 1694700623
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_246
timestamp 1694700623
transform 1 0 23736 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_254
timestamp 1694700623
transform 1 0 24472 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_267
timestamp 1694700623
transform 1 0 25668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1694700623
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1694700623
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1694700623
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1694700623
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_317
timestamp 1694700623
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1694700623
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1694700623
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_74
timestamp 1694700623
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1694700623
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_93
timestamp 1694700623
transform 1 0 9660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_111
timestamp 1694700623
transform 1 0 11316 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_135
timestamp 1694700623
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1694700623
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_153
timestamp 1694700623
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_176
timestamp 1694700623
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_192
timestamp 1694700623
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_221
timestamp 1694700623
transform 1 0 21436 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_227
timestamp 1694700623
transform 1 0 21988 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1694700623
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_253
timestamp 1694700623
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_261
timestamp 1694700623
transform 1 0 25116 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_270
timestamp 1694700623
transform 1 0 25944 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_282
timestamp 1694700623
transform 1 0 27048 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_294
timestamp 1694700623
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_306
timestamp 1694700623
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_309
timestamp 1694700623
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_317
timestamp 1694700623
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1694700623
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1694700623
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1694700623
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1694700623
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1694700623
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_66
timestamp 1694700623
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_70
timestamp 1694700623
transform 1 0 7544 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_91
timestamp 1694700623
transform 1 0 9476 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1694700623
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1694700623
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_113
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_121
timestamp 1694700623
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_126
timestamp 1694700623
transform 1 0 12696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_134
timestamp 1694700623
transform 1 0 13432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_148
timestamp 1694700623
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1694700623
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_172
timestamp 1694700623
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_195
timestamp 1694700623
transform 1 0 19044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_201
timestamp 1694700623
transform 1 0 19596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1694700623
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_256
timestamp 1694700623
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_274
timestamp 1694700623
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1694700623
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1694700623
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1694700623
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_317
timestamp 1694700623
transform 1 0 30268 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_15
timestamp 1694700623
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_22
timestamp 1694700623
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_49
timestamp 1694700623
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_61
timestamp 1694700623
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_75
timestamp 1694700623
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1694700623
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_89
timestamp 1694700623
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_95
timestamp 1694700623
transform 1 0 9844 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_107
timestamp 1694700623
transform 1 0 10948 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_119
timestamp 1694700623
transform 1 0 12052 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1694700623
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1694700623
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1694700623
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_149
timestamp 1694700623
transform 1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_156
timestamp 1694700623
transform 1 0 15456 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_168
timestamp 1694700623
transform 1 0 16560 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_174
timestamp 1694700623
transform 1 0 17112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_187
timestamp 1694700623
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1694700623
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1694700623
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_209
timestamp 1694700623
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_228
timestamp 1694700623
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_232
timestamp 1694700623
transform 1 0 22448 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_238
timestamp 1694700623
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1694700623
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_253
timestamp 1694700623
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_261
timestamp 1694700623
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1694700623
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1694700623
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1694700623
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1694700623
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_309
timestamp 1694700623
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_317
timestamp 1694700623
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 1694700623
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_42
timestamp 1694700623
transform 1 0 4968 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_90
timestamp 1694700623
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_101
timestamp 1694700623
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1694700623
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_134
timestamp 1694700623
transform 1 0 13432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_146
timestamp 1694700623
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 1694700623
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1694700623
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1694700623
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_180
timestamp 1694700623
transform 1 0 17664 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_192
timestamp 1694700623
transform 1 0 18768 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_204
timestamp 1694700623
transform 1 0 19872 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_216
timestamp 1694700623
transform 1 0 20976 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_225
timestamp 1694700623
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_252
timestamp 1694700623
transform 1 0 24288 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_265
timestamp 1694700623
transform 1 0 25484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_274
timestamp 1694700623
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1694700623
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1694700623
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1694700623
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_317
timestamp 1694700623
transform 1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1694700623
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1694700623
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1694700623
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_53
timestamp 1694700623
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_57
timestamp 1694700623
transform 1 0 6348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_70
timestamp 1694700623
transform 1 0 7544 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1694700623
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_88
timestamp 1694700623
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_96
timestamp 1694700623
transform 1 0 9936 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_104
timestamp 1694700623
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_116
timestamp 1694700623
transform 1 0 11776 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_122
timestamp 1694700623
transform 1 0 12328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1694700623
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_141
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_153
timestamp 1694700623
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_162
timestamp 1694700623
transform 1 0 16008 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_166
timestamp 1694700623
transform 1 0 16376 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_223
timestamp 1694700623
transform 1 0 21620 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_231
timestamp 1694700623
transform 1 0 22356 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_236
timestamp 1694700623
transform 1 0 22816 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 1694700623
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1694700623
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_260
timestamp 1694700623
transform 1 0 25024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_266
timestamp 1694700623
transform 1 0 25576 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_271
timestamp 1694700623
transform 1 0 26036 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_283
timestamp 1694700623
transform 1 0 27140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_295
timestamp 1694700623
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1694700623
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_309
timestamp 1694700623
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_317
timestamp 1694700623
transform 1 0 30268 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_15
timestamp 1694700623
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_20
timestamp 1694700623
transform 1 0 2944 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_25
timestamp 1694700623
transform 1 0 3404 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_31
timestamp 1694700623
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_70
timestamp 1694700623
transform 1 0 7544 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_102
timestamp 1694700623
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1694700623
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_125
timestamp 1694700623
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_130
timestamp 1694700623
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_140
timestamp 1694700623
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_155
timestamp 1694700623
transform 1 0 15364 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_159
timestamp 1694700623
transform 1 0 15732 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_166
timestamp 1694700623
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_169
timestamp 1694700623
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_175
timestamp 1694700623
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_179
timestamp 1694700623
transform 1 0 17572 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_183
timestamp 1694700623
transform 1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_207
timestamp 1694700623
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1694700623
transform 1 0 21436 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1694700623
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_249
timestamp 1694700623
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_256
timestamp 1694700623
transform 1 0 24656 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_267
timestamp 1694700623
transform 1 0 25668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1694700623
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1694700623
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1694700623
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1694700623
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_317
timestamp 1694700623
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1694700623
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_38
timestamp 1694700623
transform 1 0 4600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_66
timestamp 1694700623
transform 1 0 7176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_93
timestamp 1694700623
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_107
timestamp 1694700623
transform 1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_115
timestamp 1694700623
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_129
timestamp 1694700623
transform 1 0 12972 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1694700623
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp 1694700623
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_149
timestamp 1694700623
transform 1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_158
timestamp 1694700623
transform 1 0 15640 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_165
timestamp 1694700623
transform 1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_171
timestamp 1694700623
transform 1 0 16836 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_177
timestamp 1694700623
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_181
timestamp 1694700623
transform 1 0 17756 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1694700623
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_204
timestamp 1694700623
transform 1 0 19872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_226
timestamp 1694700623
transform 1 0 21896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_235
timestamp 1694700623
transform 1 0 22724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_243
timestamp 1694700623
transform 1 0 23460 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_253
timestamp 1694700623
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_269
timestamp 1694700623
transform 1 0 25852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_281
timestamp 1694700623
transform 1 0 26956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_293
timestamp 1694700623
transform 1 0 28060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1694700623
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1694700623
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_317
timestamp 1694700623
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_15
timestamp 1694700623
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_21
timestamp 1694700623
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_25
timestamp 1694700623
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_37
timestamp 1694700623
transform 1 0 4508 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_43
timestamp 1694700623
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_64
timestamp 1694700623
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_76
timestamp 1694700623
transform 1 0 8096 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_88
timestamp 1694700623
transform 1 0 9200 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_99
timestamp 1694700623
transform 1 0 10212 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_107
timestamp 1694700623
transform 1 0 10948 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_139
timestamp 1694700623
transform 1 0 13892 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_151
timestamp 1694700623
transform 1 0 14996 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_163
timestamp 1694700623
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1694700623
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_182
timestamp 1694700623
transform 1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_209
timestamp 1694700623
transform 1 0 20332 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_225
timestamp 1694700623
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_248
timestamp 1694700623
transform 1 0 23920 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_254
timestamp 1694700623
transform 1 0 24472 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_266
timestamp 1694700623
transform 1 0 25576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1694700623
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1694700623
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1694700623
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1694700623
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_317
timestamp 1694700623
transform 1 0 30268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1694700623
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_38
timestamp 1694700623
transform 1 0 4600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_60
timestamp 1694700623
transform 1 0 6624 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_71
timestamp 1694700623
transform 1 0 7636 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1694700623
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_95
timestamp 1694700623
transform 1 0 9844 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_107
timestamp 1694700623
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_119
timestamp 1694700623
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_131
timestamp 1694700623
transform 1 0 13156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1694700623
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1694700623
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_157
timestamp 1694700623
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_169
timestamp 1694700623
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 1694700623
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_183
timestamp 1694700623
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1694700623
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_221
timestamp 1694700623
transform 1 0 21436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_227
timestamp 1694700623
transform 1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_235
timestamp 1694700623
transform 1 0 22724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_241
timestamp 1694700623
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1694700623
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1694700623
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1694700623
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1694700623
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1694700623
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1694700623
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1694700623
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_309
timestamp 1694700623
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_317
timestamp 1694700623
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1694700623
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_19
timestamp 1694700623
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_31
timestamp 1694700623
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_47
timestamp 1694700623
transform 1 0 5428 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_80
timestamp 1694700623
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_100
timestamp 1694700623
transform 1 0 10304 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_117
timestamp 1694700623
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_122
timestamp 1694700623
transform 1 0 12328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_134
timestamp 1694700623
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_144
timestamp 1694700623
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1694700623
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1694700623
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_182
timestamp 1694700623
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_210
timestamp 1694700623
transform 1 0 20424 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_218
timestamp 1694700623
transform 1 0 21160 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1694700623
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1694700623
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_246
timestamp 1694700623
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_250
timestamp 1694700623
transform 1 0 24104 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_268
timestamp 1694700623
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_272
timestamp 1694700623
transform 1 0 26128 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1694700623
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1694700623
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1694700623
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_317
timestamp 1694700623
transform 1 0 30268 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1694700623
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1694700623
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1694700623
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_51
timestamp 1694700623
transform 1 0 5796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_65
timestamp 1694700623
transform 1 0 7084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1694700623
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1694700623
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1694700623
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1694700623
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_149
timestamp 1694700623
transform 1 0 14812 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_157
timestamp 1694700623
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_169
timestamp 1694700623
transform 1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_174
timestamp 1694700623
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1694700623
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1694700623
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_197
timestamp 1694700623
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_248
timestamp 1694700623
transform 1 0 23920 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1694700623
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_262
timestamp 1694700623
transform 1 0 25208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_267
timestamp 1694700623
transform 1 0 25668 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_280
timestamp 1694700623
transform 1 0 26864 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_292
timestamp 1694700623
transform 1 0 27968 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_304
timestamp 1694700623
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1694700623
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_317
timestamp 1694700623
transform 1 0 30268 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_13
timestamp 1694700623
transform 1 0 2300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_17
timestamp 1694700623
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_64
timestamp 1694700623
transform 1 0 6992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_76
timestamp 1694700623
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_85
timestamp 1694700623
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_100
timestamp 1694700623
transform 1 0 10304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1694700623
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_122
timestamp 1694700623
transform 1 0 12328 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_128
timestamp 1694700623
transform 1 0 12880 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_135
timestamp 1694700623
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_145
timestamp 1694700623
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_159
timestamp 1694700623
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1694700623
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_202
timestamp 1694700623
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_215
timestamp 1694700623
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1694700623
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1694700623
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_242
timestamp 1694700623
transform 1 0 23368 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_254
timestamp 1694700623
transform 1 0 24472 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_262
timestamp 1694700623
transform 1 0 25208 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_270
timestamp 1694700623
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_277
timestamp 1694700623
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1694700623
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1694700623
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1694700623
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_317
timestamp 1694700623
transform 1 0 30268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 1694700623
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_44
timestamp 1694700623
transform 1 0 5152 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_64
timestamp 1694700623
transform 1 0 6992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1694700623
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_101
timestamp 1694700623
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_128
timestamp 1694700623
transform 1 0 12880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1694700623
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_163
timestamp 1694700623
transform 1 0 16100 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_176
timestamp 1694700623
transform 1 0 17296 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 1694700623
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_209
timestamp 1694700623
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_217
timestamp 1694700623
transform 1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_227
timestamp 1694700623
transform 1 0 21988 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_242
timestamp 1694700623
transform 1 0 23368 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1694700623
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_275
timestamp 1694700623
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_292
timestamp 1694700623
transform 1 0 27968 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_304
timestamp 1694700623
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_309
timestamp 1694700623
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_317
timestamp 1694700623
transform 1 0 30268 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_15
timestamp 1694700623
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_21
timestamp 1694700623
transform 1 0 3036 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_31
timestamp 1694700623
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_43
timestamp 1694700623
transform 1 0 5060 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_51
timestamp 1694700623
transform 1 0 5796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1694700623
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_81
timestamp 1694700623
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_89
timestamp 1694700623
transform 1 0 9292 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_146
timestamp 1694700623
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_156
timestamp 1694700623
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_163
timestamp 1694700623
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1694700623
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 1694700623
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 1694700623
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1694700623
transform 1 0 19596 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_211
timestamp 1694700623
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1694700623
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_235
timestamp 1694700623
transform 1 0 22724 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_247
timestamp 1694700623
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_259
timestamp 1694700623
transform 1 0 24932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_265
timestamp 1694700623
transform 1 0 25484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1694700623
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_281
timestamp 1694700623
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_296
timestamp 1694700623
transform 1 0 28336 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_308
timestamp 1694700623
transform 1 0 29440 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1694700623
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1694700623
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_58
timestamp 1694700623
transform 1 0 6440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_80
timestamp 1694700623
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_91
timestamp 1694700623
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_107
timestamp 1694700623
transform 1 0 10948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_150
timestamp 1694700623
transform 1 0 14904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_182
timestamp 1694700623
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_191
timestamp 1694700623
transform 1 0 18676 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_217
timestamp 1694700623
transform 1 0 21068 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_223
timestamp 1694700623
transform 1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_229
timestamp 1694700623
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1694700623
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1694700623
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_267
timestamp 1694700623
transform 1 0 25668 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_271
timestamp 1694700623
transform 1 0 26036 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_276
timestamp 1694700623
transform 1 0 26496 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_282
timestamp 1694700623
transform 1 0 27048 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1694700623
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1694700623
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1694700623
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_309
timestamp 1694700623
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_317
timestamp 1694700623
transform 1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1694700623
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_46
timestamp 1694700623
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_64
timestamp 1694700623
transform 1 0 6992 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_72
timestamp 1694700623
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_86
timestamp 1694700623
transform 1 0 9016 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_98
timestamp 1694700623
transform 1 0 10120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1694700623
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1694700623
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1694700623
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_175
timestamp 1694700623
transform 1 0 17204 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_195
timestamp 1694700623
transform 1 0 19044 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_203
timestamp 1694700623
transform 1 0 19780 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_209
timestamp 1694700623
transform 1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1694700623
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_237
timestamp 1694700623
transform 1 0 22908 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_241
timestamp 1694700623
transform 1 0 23276 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_250
timestamp 1694700623
transform 1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_258
timestamp 1694700623
transform 1 0 24840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_275
timestamp 1694700623
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1694700623
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_296
timestamp 1694700623
transform 1 0 28336 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_308
timestamp 1694700623
transform 1 0 29440 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1694700623
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_38
timestamp 1694700623
transform 1 0 4600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_46
timestamp 1694700623
transform 1 0 5336 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_53
timestamp 1694700623
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_61
timestamp 1694700623
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_69
timestamp 1694700623
transform 1 0 7452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_77
timestamp 1694700623
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1694700623
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1694700623
transform 1 0 11316 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_118
timestamp 1694700623
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_144
timestamp 1694700623
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_152
timestamp 1694700623
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_159
timestamp 1694700623
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_171
timestamp 1694700623
transform 1 0 16836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_183
timestamp 1694700623
transform 1 0 17940 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_204
timestamp 1694700623
transform 1 0 19872 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_253
timestamp 1694700623
transform 1 0 24380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1694700623
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1694700623
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_317
timestamp 1694700623
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1694700623
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_27
timestamp 1694700623
transform 1 0 3588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp 1694700623
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_63
timestamp 1694700623
transform 1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_70
timestamp 1694700623
transform 1 0 7544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_82
timestamp 1694700623
transform 1 0 8648 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 1694700623
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1694700623
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1694700623
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1694700623
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_184
timestamp 1694700623
transform 1 0 18032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_196
timestamp 1694700623
transform 1 0 19136 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_201
timestamp 1694700623
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_205
timestamp 1694700623
transform 1 0 19964 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_218
timestamp 1694700623
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_266
timestamp 1694700623
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1694700623
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_281
timestamp 1694700623
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_291
timestamp 1694700623
transform 1 0 27876 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_303
timestamp 1694700623
transform 1 0 28980 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_315
timestamp 1694700623
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_319
timestamp 1694700623
transform 1 0 30452 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1694700623
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1694700623
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1694700623
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_49
timestamp 1694700623
transform 1 0 5612 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_53
timestamp 1694700623
transform 1 0 5980 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_70
timestamp 1694700623
transform 1 0 7544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_90
timestamp 1694700623
transform 1 0 9384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_98
timestamp 1694700623
transform 1 0 10120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_117
timestamp 1694700623
transform 1 0 11868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_123
timestamp 1694700623
transform 1 0 12420 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_132
timestamp 1694700623
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1694700623
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_153
timestamp 1694700623
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_161
timestamp 1694700623
transform 1 0 15916 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_218
timestamp 1694700623
transform 1 0 21160 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_230
timestamp 1694700623
transform 1 0 22264 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1694700623
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1694700623
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_253
timestamp 1694700623
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_260
timestamp 1694700623
transform 1 0 25024 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_295
timestamp 1694700623
transform 1 0 28244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_299
timestamp 1694700623
transform 1 0 28612 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1694700623
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_315
timestamp 1694700623
transform 1 0 30084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_319
timestamp 1694700623
transform 1 0 30452 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1694700623
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_15
timestamp 1694700623
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_37
timestamp 1694700623
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_49
timestamp 1694700623
transform 1 0 5612 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1694700623
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_65
timestamp 1694700623
transform 1 0 7084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_77
timestamp 1694700623
transform 1 0 8188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_101
timestamp 1694700623
transform 1 0 10396 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_108
timestamp 1694700623
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_120
timestamp 1694700623
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_131
timestamp 1694700623
transform 1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_151
timestamp 1694700623
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_169
timestamp 1694700623
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_173
timestamp 1694700623
transform 1 0 17020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_185
timestamp 1694700623
transform 1 0 18124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_197
timestamp 1694700623
transform 1 0 19228 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1694700623
transform 1 0 19596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_220
timestamp 1694700623
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_237
timestamp 1694700623
transform 1 0 22908 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_245
timestamp 1694700623
transform 1 0 23644 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_277
timestamp 1694700623
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_298
timestamp 1694700623
transform 1 0 28520 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_304
timestamp 1694700623
transform 1 0 29072 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_308
timestamp 1694700623
transform 1 0 29440 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_7
timestamp 1694700623
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_19
timestamp 1694700623
transform 1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1694700623
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_39
timestamp 1694700623
transform 1 0 4692 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_63
timestamp 1694700623
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_75
timestamp 1694700623
transform 1 0 8004 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1694700623
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1694700623
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_109
timestamp 1694700623
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_144
timestamp 1694700623
transform 1 0 14352 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_166
timestamp 1694700623
transform 1 0 16376 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_180
timestamp 1694700623
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_185
timestamp 1694700623
transform 1 0 18124 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_189
timestamp 1694700623
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_203
timestamp 1694700623
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_213
timestamp 1694700623
transform 1 0 20700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_225
timestamp 1694700623
transform 1 0 21804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1694700623
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1694700623
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_256
timestamp 1694700623
transform 1 0 24656 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_268
timestamp 1694700623
transform 1 0 25760 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_280
timestamp 1694700623
transform 1 0 26864 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_289
timestamp 1694700623
transform 1 0 27692 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_297
timestamp 1694700623
transform 1 0 28428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_301
timestamp 1694700623
transform 1 0 28796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1694700623
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_309
timestamp 1694700623
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_317
timestamp 1694700623
transform 1 0 30268 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 1694700623
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_19
timestamp 1694700623
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_31
timestamp 1694700623
transform 1 0 3956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_35
timestamp 1694700623
transform 1 0 4324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_44
timestamp 1694700623
transform 1 0 5152 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1694700623
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1694700623
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_66
timestamp 1694700623
transform 1 0 7176 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_99
timestamp 1694700623
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1694700623
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_113
timestamp 1694700623
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1694700623
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_126
timestamp 1694700623
transform 1 0 12696 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_132
timestamp 1694700623
transform 1 0 13248 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_141
timestamp 1694700623
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1694700623
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_169
timestamp 1694700623
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_178
timestamp 1694700623
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_200
timestamp 1694700623
transform 1 0 19504 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1694700623
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_245
timestamp 1694700623
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_269
timestamp 1694700623
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_293
timestamp 1694700623
transform 1 0 28060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_301
timestamp 1694700623
transform 1 0 28796 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_318
timestamp 1694700623
transform 1 0 30360 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1694700623
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_19
timestamp 1694700623
transform 1 0 2852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_24
timestamp 1694700623
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_32
timestamp 1694700623
transform 1 0 4048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_38
timestamp 1694700623
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_46
timestamp 1694700623
transform 1 0 5336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_58
timestamp 1694700623
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1694700623
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_100
timestamp 1694700623
transform 1 0 10304 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_116
timestamp 1694700623
transform 1 0 11776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_131
timestamp 1694700623
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1694700623
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1694700623
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_153
timestamp 1694700623
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_161
timestamp 1694700623
transform 1 0 15916 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_167
timestamp 1694700623
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_171
timestamp 1694700623
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1694700623
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_189
timestamp 1694700623
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1694700623
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_200
timestamp 1694700623
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_249
timestamp 1694700623
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_253
timestamp 1694700623
transform 1 0 24380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_287
timestamp 1694700623
transform 1 0 27508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1694700623
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_309
timestamp 1694700623
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_317
timestamp 1694700623
transform 1 0 30268 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1694700623
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1694700623
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1694700623
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1694700623
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_74
timestamp 1694700623
transform 1 0 7912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_86
timestamp 1694700623
transform 1 0 9016 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_98
timestamp 1694700623
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1694700623
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_116
timestamp 1694700623
transform 1 0 11776 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_133
timestamp 1694700623
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_162
timestamp 1694700623
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1694700623
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_178
timestamp 1694700623
transform 1 0 17480 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_202
timestamp 1694700623
transform 1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_218
timestamp 1694700623
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_249
timestamp 1694700623
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_257
timestamp 1694700623
transform 1 0 24748 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1694700623
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1694700623
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1694700623
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1694700623
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_293
timestamp 1694700623
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_297
timestamp 1694700623
transform 1 0 28428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_318
timestamp 1694700623
transform 1 0 30360 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1694700623
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1694700623
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1694700623
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1694700623
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_52
timestamp 1694700623
transform 1 0 5888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_65
timestamp 1694700623
transform 1 0 7084 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_74
timestamp 1694700623
transform 1 0 7912 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1694700623
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_103
timestamp 1694700623
transform 1 0 10580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1694700623
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_132
timestamp 1694700623
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_141
timestamp 1694700623
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_181
timestamp 1694700623
transform 1 0 17756 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_187
timestamp 1694700623
transform 1 0 18308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_224
timestamp 1694700623
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1694700623
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1694700623
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_257
timestamp 1694700623
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_300
timestamp 1694700623
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_309
timestamp 1694700623
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_317
timestamp 1694700623
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 1694700623
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 1694700623
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_31
timestamp 1694700623
transform 1 0 3956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_37
timestamp 1694700623
transform 1 0 4508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1694700623
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1694700623
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_64
timestamp 1694700623
transform 1 0 6992 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_70
timestamp 1694700623
transform 1 0 7544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_97
timestamp 1694700623
transform 1 0 10028 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1694700623
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1694700623
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_125
timestamp 1694700623
transform 1 0 12604 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_143
timestamp 1694700623
transform 1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_158
timestamp 1694700623
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1694700623
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_172
timestamp 1694700623
transform 1 0 16928 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_212
timestamp 1694700623
transform 1 0 20608 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1694700623
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1694700623
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_240
timestamp 1694700623
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_244
timestamp 1694700623
transform 1 0 23552 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1694700623
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_291
timestamp 1694700623
transform 1 0 27876 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_303
timestamp 1694700623
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_315
timestamp 1694700623
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_319
timestamp 1694700623
transform 1 0 30452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1694700623
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1694700623
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1694700623
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_29
timestamp 1694700623
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_42
timestamp 1694700623
transform 1 0 4968 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_54
timestamp 1694700623
transform 1 0 6072 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_66
timestamp 1694700623
transform 1 0 7176 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_78
timestamp 1694700623
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_96
timestamp 1694700623
transform 1 0 9936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_100
timestamp 1694700623
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_104
timestamp 1694700623
transform 1 0 10672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_112
timestamp 1694700623
transform 1 0 11408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_119
timestamp 1694700623
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1694700623
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_141
timestamp 1694700623
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_159
timestamp 1694700623
transform 1 0 15732 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_171
timestamp 1694700623
transform 1 0 16836 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_187
timestamp 1694700623
transform 1 0 18308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_204
timestamp 1694700623
transform 1 0 19872 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_210
timestamp 1694700623
transform 1 0 20424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_214
timestamp 1694700623
transform 1 0 20792 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_238
timestamp 1694700623
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1694700623
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_265
timestamp 1694700623
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_269
timestamp 1694700623
transform 1 0 25852 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_281
timestamp 1694700623
transform 1 0 26956 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_287
timestamp 1694700623
transform 1 0 27508 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_294
timestamp 1694700623
transform 1 0 28152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_298
timestamp 1694700623
transform 1 0 28520 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1694700623
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_316
timestamp 1694700623
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1694700623
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1694700623
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_27
timestamp 1694700623
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_37
timestamp 1694700623
transform 1 0 4508 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_50
timestamp 1694700623
transform 1 0 5704 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_78
timestamp 1694700623
transform 1 0 8280 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_87
timestamp 1694700623
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_91
timestamp 1694700623
transform 1 0 9476 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_130
timestamp 1694700623
transform 1 0 13064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_142
timestamp 1694700623
transform 1 0 14168 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_189
timestamp 1694700623
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_193
timestamp 1694700623
transform 1 0 18860 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_206
timestamp 1694700623
transform 1 0 20056 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_212
timestamp 1694700623
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1694700623
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1694700623
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_237
timestamp 1694700623
transform 1 0 22908 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_241
timestamp 1694700623
transform 1 0 23276 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_253
timestamp 1694700623
transform 1 0 24380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_270
timestamp 1694700623
transform 1 0 25944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_287
timestamp 1694700623
transform 1 0 27508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_291
timestamp 1694700623
transform 1 0 27876 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_308
timestamp 1694700623
transform 1 0 29440 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1694700623
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1694700623
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1694700623
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1694700623
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1694700623
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_53
timestamp 1694700623
transform 1 0 5980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_67
timestamp 1694700623
transform 1 0 7268 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_82
timestamp 1694700623
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1694700623
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_92
timestamp 1694700623
transform 1 0 9568 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_104
timestamp 1694700623
transform 1 0 10672 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_112
timestamp 1694700623
transform 1 0 11408 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_127
timestamp 1694700623
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_136
timestamp 1694700623
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_141
timestamp 1694700623
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_149
timestamp 1694700623
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_153
timestamp 1694700623
transform 1 0 15180 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_160
timestamp 1694700623
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_172
timestamp 1694700623
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_184
timestamp 1694700623
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1694700623
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_253
timestamp 1694700623
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_262
timestamp 1694700623
transform 1 0 25208 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_266
timestamp 1694700623
transform 1 0 25576 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_278
timestamp 1694700623
transform 1 0 26680 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_286
timestamp 1694700623
transform 1 0 27416 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_294
timestamp 1694700623
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1694700623
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_309
timestamp 1694700623
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_317
timestamp 1694700623
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1694700623
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1694700623
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1694700623
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1694700623
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_47
timestamp 1694700623
transform 1 0 5428 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_53
timestamp 1694700623
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_64
timestamp 1694700623
transform 1 0 6992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_72
timestamp 1694700623
transform 1 0 7728 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_78
timestamp 1694700623
transform 1 0 8280 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_90
timestamp 1694700623
transform 1 0 9384 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_103
timestamp 1694700623
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1694700623
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1694700623
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_125
timestamp 1694700623
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_133
timestamp 1694700623
transform 1 0 13340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_138
timestamp 1694700623
transform 1 0 13800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_150
timestamp 1694700623
transform 1 0 14904 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1694700623
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1694700623
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_181
timestamp 1694700623
transform 1 0 17756 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_203
timestamp 1694700623
transform 1 0 19780 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_211
timestamp 1694700623
transform 1 0 20516 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_215
timestamp 1694700623
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1694700623
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1694700623
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_237
timestamp 1694700623
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_246
timestamp 1694700623
transform 1 0 23736 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_274
timestamp 1694700623
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1694700623
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1694700623
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1694700623
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_317
timestamp 1694700623
transform 1 0 30268 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1694700623
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1694700623
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1694700623
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_29
timestamp 1694700623
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_35
timestamp 1694700623
transform 1 0 4324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_66
timestamp 1694700623
transform 1 0 7176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1694700623
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_92
timestamp 1694700623
transform 1 0 9568 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_100
timestamp 1694700623
transform 1 0 10304 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_124
timestamp 1694700623
transform 1 0 12512 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_132
timestamp 1694700623
transform 1 0 13248 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_136
timestamp 1694700623
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1694700623
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_172
timestamp 1694700623
transform 1 0 16928 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1694700623
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1694700623
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1694700623
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1694700623
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1694700623
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1694700623
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1694700623
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1694700623
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1694700623
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1694700623
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1694700623
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1694700623
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1694700623
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_309
timestamp 1694700623
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_317
timestamp 1694700623
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1694700623
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1694700623
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1694700623
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1694700623
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1694700623
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1694700623
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_108
timestamp 1694700623
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_113
timestamp 1694700623
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_122
timestamp 1694700623
transform 1 0 12328 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_126
timestamp 1694700623
transform 1 0 12696 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_150
timestamp 1694700623
transform 1 0 14904 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_162
timestamp 1694700623
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_196
timestamp 1694700623
transform 1 0 19136 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_208
timestamp 1694700623
transform 1 0 20240 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_220
timestamp 1694700623
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1694700623
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1694700623
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1694700623
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1694700623
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1694700623
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1694700623
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1694700623
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1694700623
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1694700623
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_317
timestamp 1694700623
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1694700623
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1694700623
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1694700623
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1694700623
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1694700623
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1694700623
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1694700623
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1694700623
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1694700623
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_85
timestamp 1694700623
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_92
timestamp 1694700623
transform 1 0 9568 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_100
timestamp 1694700623
transform 1 0 10304 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_123
timestamp 1694700623
transform 1 0 12420 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1694700623
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1694700623
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_153
timestamp 1694700623
transform 1 0 15180 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_159
timestamp 1694700623
transform 1 0 15732 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_171
timestamp 1694700623
transform 1 0 16836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_177
timestamp 1694700623
transform 1 0 17388 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_193
timestamp 1694700623
transform 1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_213
timestamp 1694700623
transform 1 0 20700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_225
timestamp 1694700623
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_237
timestamp 1694700623
transform 1 0 22908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_249
timestamp 1694700623
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1694700623
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1694700623
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1694700623
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1694700623
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1694700623
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1694700623
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1694700623
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_317
timestamp 1694700623
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1694700623
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1694700623
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1694700623
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1694700623
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1694700623
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1694700623
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1694700623
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1694700623
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1694700623
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1694700623
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1694700623
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1694700623
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_113
timestamp 1694700623
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_165
timestamp 1694700623
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_185
timestamp 1694700623
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_203
timestamp 1694700623
transform 1 0 19780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_215
timestamp 1694700623
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1694700623
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1694700623
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1694700623
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1694700623
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1694700623
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1694700623
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1694700623
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1694700623
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1694700623
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1694700623
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_317
timestamp 1694700623
transform 1 0 30268 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1694700623
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1694700623
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1694700623
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1694700623
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1694700623
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1694700623
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1694700623
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1694700623
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1694700623
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1694700623
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1694700623
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1694700623
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1694700623
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1694700623
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1694700623
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_173
timestamp 1694700623
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_191
timestamp 1694700623
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1694700623
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_205
timestamp 1694700623
transform 1 0 19964 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_217
timestamp 1694700623
transform 1 0 21068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_229
timestamp 1694700623
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_241
timestamp 1694700623
transform 1 0 23276 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_249
timestamp 1694700623
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1694700623
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1694700623
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1694700623
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1694700623
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1694700623
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1694700623
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_309
timestamp 1694700623
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_317
timestamp 1694700623
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1694700623
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1694700623
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1694700623
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1694700623
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1694700623
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1694700623
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1694700623
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1694700623
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1694700623
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1694700623
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1694700623
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1694700623
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1694700623
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1694700623
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_137
timestamp 1694700623
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_145
timestamp 1694700623
transform 1 0 14444 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_149
timestamp 1694700623
transform 1 0 14812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_153
timestamp 1694700623
transform 1 0 15180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_157
timestamp 1694700623
transform 1 0 15548 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_165
timestamp 1694700623
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_169
timestamp 1694700623
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_175
timestamp 1694700623
transform 1 0 17204 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_192
timestamp 1694700623
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_204
timestamp 1694700623
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_216
timestamp 1694700623
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1694700623
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1694700623
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1694700623
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1694700623
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1694700623
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1694700623
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1694700623
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1694700623
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1694700623
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_317
timestamp 1694700623
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1694700623
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1694700623
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1694700623
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1694700623
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1694700623
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1694700623
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1694700623
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1694700623
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1694700623
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1694700623
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1694700623
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1694700623
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1694700623
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1694700623
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1694700623
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1694700623
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1694700623
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1694700623
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1694700623
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1694700623
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1694700623
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1694700623
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1694700623
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1694700623
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1694700623
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1694700623
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1694700623
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1694700623
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1694700623
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1694700623
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1694700623
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1694700623
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1694700623
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_309
timestamp 1694700623
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_317
timestamp 1694700623
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1694700623
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1694700623
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1694700623
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1694700623
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1694700623
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1694700623
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1694700623
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1694700623
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1694700623
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1694700623
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1694700623
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1694700623
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1694700623
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1694700623
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1694700623
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1694700623
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1694700623
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1694700623
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1694700623
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1694700623
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1694700623
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1694700623
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1694700623
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1694700623
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1694700623
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1694700623
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1694700623
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1694700623
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1694700623
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1694700623
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1694700623
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1694700623
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1694700623
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_317
timestamp 1694700623
transform 1 0 30268 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1694700623
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1694700623
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1694700623
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1694700623
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1694700623
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1694700623
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1694700623
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1694700623
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1694700623
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1694700623
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1694700623
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1694700623
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1694700623
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1694700623
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1694700623
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1694700623
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1694700623
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1694700623
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1694700623
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1694700623
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1694700623
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1694700623
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1694700623
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1694700623
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1694700623
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1694700623
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1694700623
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1694700623
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1694700623
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1694700623
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1694700623
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1694700623
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1694700623
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_309
timestamp 1694700623
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_317
timestamp 1694700623
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1694700623
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1694700623
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_27
timestamp 1694700623
transform 1 0 3588 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_29
timestamp 1694700623
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_41
timestamp 1694700623
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1694700623
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1694700623
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1694700623
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_81
timestamp 1694700623
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_85
timestamp 1694700623
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_97
timestamp 1694700623
transform 1 0 10028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1694700623
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1694700623
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_125
timestamp 1694700623
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_135
timestamp 1694700623
transform 1 0 13524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_139
timestamp 1694700623
transform 1 0 13892 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_141
timestamp 1694700623
transform 1 0 14076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_153
timestamp 1694700623
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 1694700623
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1694700623
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1694700623
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_181
timestamp 1694700623
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_191
timestamp 1694700623
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_195
timestamp 1694700623
transform 1 0 19044 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_197
timestamp 1694700623
transform 1 0 19228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_209
timestamp 1694700623
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1694700623
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1694700623
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1694700623
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_249
timestamp 1694700623
transform 1 0 24012 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_253
timestamp 1694700623
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_265
timestamp 1694700623
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 1694700623
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1694700623
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1694700623
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_305
timestamp 1694700623
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_309
timestamp 1694700623
transform 1 0 29532 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_317
timestamp 1694700623
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1694700623
transform -1 0 18860 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1694700623
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1694700623
transform -1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1694700623
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1694700623
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1694700623
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1694700623
transform -1 0 19228 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1694700623
transform -1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1694700623
transform -1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1694700623
transform -1 0 18768 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1694700623
transform -1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1694700623
transform -1 0 8280 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1694700623
transform -1 0 7544 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1694700623
transform 1 0 9568 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1694700623
transform -1 0 5152 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1694700623
transform -1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1694700623
transform -1 0 14076 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output2
timestamp 1694700623
transform -1 0 18676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 1694700623
transform 1 0 12972 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1694700623
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1694700623
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1694700623
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1694700623
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1694700623
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 1694700623
transform -1 0 16100 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_50
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_51
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_52
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_53
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_54
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_55
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_56
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_57
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_58
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_59
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_60
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_61
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_62
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_63
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_64
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_65
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_66
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_67
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_68
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_69
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_70
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_71
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_72
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_73
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_74
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_75
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_76
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_77
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_78
timestamp 1694700623
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1694700623
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_79
timestamp 1694700623
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1694700623
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_80
timestamp 1694700623
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1694700623
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_81
timestamp 1694700623
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1694700623
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_82
timestamp 1694700623
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1694700623
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_83
timestamp 1694700623
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1694700623
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_84
timestamp 1694700623
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1694700623
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_85
timestamp 1694700623
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1694700623
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_86
timestamp 1694700623
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1694700623
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_87
timestamp 1694700623
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1694700623
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_88
timestamp 1694700623
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1694700623
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_89
timestamp 1694700623
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1694700623
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_90
timestamp 1694700623
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1694700623
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_91
timestamp 1694700623
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1694700623
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_92
timestamp 1694700623
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1694700623
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_93
timestamp 1694700623
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1694700623
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_94
timestamp 1694700623
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1694700623
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_95
timestamp 1694700623
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1694700623
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_96
timestamp 1694700623
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1694700623
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_97
timestamp 1694700623
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1694700623
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_98
timestamp 1694700623
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1694700623
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_99
timestamp 1694700623
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1694700623
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1694700623
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1694700623
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1694700623
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1694700623
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1694700623
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1694700623
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp 1694700623
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_113
timestamp 1694700623
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_114
timestamp 1694700623
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_115
timestamp 1694700623
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_118
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_119
timestamp 1694700623
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_120
timestamp 1694700623
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_121
timestamp 1694700623
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_123
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp 1694700623
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_125
timestamp 1694700623
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_126
timestamp 1694700623
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_128
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_129
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_130
timestamp 1694700623
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_131
timestamp 1694700623
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_132
timestamp 1694700623
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_133
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_134
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_135
timestamp 1694700623
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_136
timestamp 1694700623
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_137
timestamp 1694700623
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_138
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_139
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_140
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_141
timestamp 1694700623
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_142
timestamp 1694700623
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_143
timestamp 1694700623
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_144
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_145
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_146
timestamp 1694700623
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_147
timestamp 1694700623
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_148
timestamp 1694700623
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_149
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_150
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_151
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_152
timestamp 1694700623
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_153
timestamp 1694700623
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_154
timestamp 1694700623
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_155
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_156
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_157
timestamp 1694700623
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_158
timestamp 1694700623
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_159
timestamp 1694700623
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_160
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_161
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_162
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_163
timestamp 1694700623
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_164
timestamp 1694700623
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_165
timestamp 1694700623
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_166
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_167
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_168
timestamp 1694700623
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_169
timestamp 1694700623
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_170
timestamp 1694700623
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_171
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_172
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_173
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_174
timestamp 1694700623
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_175
timestamp 1694700623
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_176
timestamp 1694700623
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_177
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_178
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_179
timestamp 1694700623
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_180
timestamp 1694700623
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_181
timestamp 1694700623
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_182
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_183
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_184
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_185
timestamp 1694700623
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_186
timestamp 1694700623
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_187
timestamp 1694700623
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_188
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_189
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_190
timestamp 1694700623
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_191
timestamp 1694700623
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_192
timestamp 1694700623
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_193
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_194
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_195
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_196
timestamp 1694700623
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_197
timestamp 1694700623
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_198
timestamp 1694700623
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_199
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_200
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_201
timestamp 1694700623
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_202
timestamp 1694700623
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_203
timestamp 1694700623
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_204
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_205
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_206
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_207
timestamp 1694700623
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_208
timestamp 1694700623
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_209
timestamp 1694700623
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_210
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_211
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_212
timestamp 1694700623
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_213
timestamp 1694700623
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_214
timestamp 1694700623
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_215
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_216
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_217
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_218
timestamp 1694700623
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_219
timestamp 1694700623
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_220
timestamp 1694700623
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_221
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_222
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_223
timestamp 1694700623
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_224
timestamp 1694700623
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_225
timestamp 1694700623
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_226
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_227
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_228
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_229
timestamp 1694700623
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_230
timestamp 1694700623
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_231
timestamp 1694700623
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_232
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_233
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_234
timestamp 1694700623
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_235
timestamp 1694700623
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_236
timestamp 1694700623
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_237
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_238
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_239
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_240
timestamp 1694700623
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_241
timestamp 1694700623
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_242
timestamp 1694700623
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_243
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_244
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_245
timestamp 1694700623
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_246
timestamp 1694700623
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_247
timestamp 1694700623
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_248
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_249
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_250
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_251
timestamp 1694700623
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_252
timestamp 1694700623
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_253
timestamp 1694700623
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_254
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_255
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_256
timestamp 1694700623
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_257
timestamp 1694700623
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_258
timestamp 1694700623
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_259
timestamp 1694700623
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_260
timestamp 1694700623
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_261
timestamp 1694700623
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_262
timestamp 1694700623
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_263
timestamp 1694700623
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_264
timestamp 1694700623
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_265
timestamp 1694700623
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_266
timestamp 1694700623
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_267
timestamp 1694700623
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_268
timestamp 1694700623
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_269
timestamp 1694700623
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_270
timestamp 1694700623
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_271
timestamp 1694700623
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_272
timestamp 1694700623
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_273
timestamp 1694700623
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_274
timestamp 1694700623
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_275
timestamp 1694700623
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_276
timestamp 1694700623
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_277
timestamp 1694700623
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_278
timestamp 1694700623
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_279
timestamp 1694700623
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_280
timestamp 1694700623
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_281
timestamp 1694700623
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_282
timestamp 1694700623
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_283
timestamp 1694700623
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_284
timestamp 1694700623
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_285
timestamp 1694700623
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_286
timestamp 1694700623
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_287
timestamp 1694700623
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_288
timestamp 1694700623
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_289
timestamp 1694700623
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_290
timestamp 1694700623
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_291
timestamp 1694700623
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_292
timestamp 1694700623
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_293
timestamp 1694700623
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_294
timestamp 1694700623
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_295
timestamp 1694700623
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_296
timestamp 1694700623
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_297
timestamp 1694700623
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_298
timestamp 1694700623
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_299
timestamp 1694700623
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_300
timestamp 1694700623
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_301
timestamp 1694700623
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_302
timestamp 1694700623
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_303
timestamp 1694700623
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_304
timestamp 1694700623
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_305
timestamp 1694700623
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_306
timestamp 1694700623
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_307
timestamp 1694700623
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_308
timestamp 1694700623
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_309
timestamp 1694700623
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_310
timestamp 1694700623
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_311
timestamp 1694700623
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_312
timestamp 1694700623
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_313
timestamp 1694700623
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_314
timestamp 1694700623
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_315
timestamp 1694700623
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_316
timestamp 1694700623
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_317
timestamp 1694700623
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_318
timestamp 1694700623
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_319
timestamp 1694700623
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_320
timestamp 1694700623
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_321
timestamp 1694700623
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_322
timestamp 1694700623
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_323
timestamp 1694700623
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_324
timestamp 1694700623
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_325
timestamp 1694700623
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_326
timestamp 1694700623
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_327
timestamp 1694700623
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_328
timestamp 1694700623
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_329
timestamp 1694700623
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_330
timestamp 1694700623
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_331
timestamp 1694700623
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_332
timestamp 1694700623
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_333
timestamp 1694700623
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_334
timestamp 1694700623
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_335
timestamp 1694700623
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_336
timestamp 1694700623
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_337
timestamp 1694700623
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_338
timestamp 1694700623
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_339
timestamp 1694700623
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_340
timestamp 1694700623
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_341
timestamp 1694700623
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_342
timestamp 1694700623
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_343
timestamp 1694700623
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_344
timestamp 1694700623
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_345
timestamp 1694700623
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_346
timestamp 1694700623
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_347
timestamp 1694700623
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_348
timestamp 1694700623
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_349
timestamp 1694700623
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_350
timestamp 1694700623
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_351
timestamp 1694700623
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_352
timestamp 1694700623
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_353
timestamp 1694700623
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_354
timestamp 1694700623
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_355
timestamp 1694700623
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_356
timestamp 1694700623
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_357
timestamp 1694700623
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_358
timestamp 1694700623
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_359
timestamp 1694700623
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_360
timestamp 1694700623
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_361
timestamp 1694700623
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_362
timestamp 1694700623
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_363
timestamp 1694700623
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_364
timestamp 1694700623
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_365
timestamp 1694700623
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_366
timestamp 1694700623
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_367
timestamp 1694700623
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_368
timestamp 1694700623
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_369
timestamp 1694700623
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_370
timestamp 1694700623
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_371
timestamp 1694700623
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_372
timestamp 1694700623
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_373
timestamp 1694700623
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_374
timestamp 1694700623
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_375
timestamp 1694700623
transform 1 0 3680 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_376
timestamp 1694700623
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_377
timestamp 1694700623
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_378
timestamp 1694700623
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_379
timestamp 1694700623
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_380
timestamp 1694700623
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_381
timestamp 1694700623
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_382
timestamp 1694700623
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_383
timestamp 1694700623
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_384
timestamp 1694700623
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_385
timestamp 1694700623
transform 1 0 29440 0 -1 29376
box -38 -48 130 592
<< labels >>
flabel metal4 s 5318 2128 5638 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12746 2128 13066 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 20174 2128 20494 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27602 2128 27922 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6076 30868 6396 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12876 30868 13196 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 19676 30868 19996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 26476 30868 26796 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4658 2128 4978 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12086 2128 12406 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19514 2128 19834 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26942 2128 27262 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5416 30868 5736 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12216 30868 12536 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 19016 30868 19336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 25816 30868 26136 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 clock
port 2 nsew signal input
flabel metal2 s 18050 31200 18106 32000 0 FreeSans 224 90 0 0 logisim_clock_tree_0_out
port 3 nsew signal tristate
flabel metal2 s 12898 31200 12954 32000 0 FreeSans 224 90 0 0 ram_addr_o[0]
port 4 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 ram_addr_o[1]
port 5 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 ram_addr_o[2]
port 6 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 ram_addr_o[3]
port 7 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 ram_addr_o[4]
port 8 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 ram_data_io[0]
port 9 nsew signal bidirectional
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 ram_data_io[10]
port 10 nsew signal bidirectional
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 ram_data_io[11]
port 11 nsew signal bidirectional
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 ram_data_io[12]
port 12 nsew signal bidirectional
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 ram_data_io[13]
port 13 nsew signal bidirectional
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 ram_data_io[14]
port 14 nsew signal bidirectional
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 ram_data_io[15]
port 15 nsew signal bidirectional
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 ram_data_io[16]
port 16 nsew signal bidirectional
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 ram_data_io[17]
port 17 nsew signal bidirectional
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 ram_data_io[18]
port 18 nsew signal bidirectional
flabel metal3 s 31200 10888 32000 11008 0 FreeSans 480 0 0 0 ram_data_io[19]
port 19 nsew signal bidirectional
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 ram_data_io[1]
port 20 nsew signal bidirectional
flabel metal3 s 31200 13608 32000 13728 0 FreeSans 480 0 0 0 ram_data_io[20]
port 21 nsew signal bidirectional
flabel metal3 s 31200 15648 32000 15768 0 FreeSans 480 0 0 0 ram_data_io[21]
port 22 nsew signal bidirectional
flabel metal3 s 31200 17008 32000 17128 0 FreeSans 480 0 0 0 ram_data_io[22]
port 23 nsew signal bidirectional
flabel metal3 s 31200 16328 32000 16448 0 FreeSans 480 0 0 0 ram_data_io[23]
port 24 nsew signal bidirectional
flabel metal3 s 31200 18368 32000 18488 0 FreeSans 480 0 0 0 ram_data_io[24]
port 25 nsew signal bidirectional
flabel metal3 s 31200 19728 32000 19848 0 FreeSans 480 0 0 0 ram_data_io[25]
port 26 nsew signal bidirectional
flabel metal3 s 31200 21088 32000 21208 0 FreeSans 480 0 0 0 ram_data_io[26]
port 27 nsew signal bidirectional
flabel metal3 s 31200 21768 32000 21888 0 FreeSans 480 0 0 0 ram_data_io[27]
port 28 nsew signal bidirectional
flabel metal3 s 31200 20408 32000 20528 0 FreeSans 480 0 0 0 ram_data_io[28]
port 29 nsew signal bidirectional
flabel metal2 s 20626 31200 20682 32000 0 FreeSans 224 90 0 0 ram_data_io[29]
port 30 nsew signal bidirectional
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 ram_data_io[2]
port 31 nsew signal bidirectional
flabel metal3 s 31200 17688 32000 17808 0 FreeSans 480 0 0 0 ram_data_io[30]
port 32 nsew signal bidirectional
flabel metal2 s 14830 31200 14886 32000 0 FreeSans 224 90 0 0 ram_data_io[31]
port 33 nsew signal bidirectional
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 ram_data_io[3]
port 34 nsew signal bidirectional
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 ram_data_io[4]
port 35 nsew signal bidirectional
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 ram_data_io[5]
port 36 nsew signal bidirectional
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 ram_data_io[6]
port 37 nsew signal bidirectional
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 ram_data_io[7]
port 38 nsew signal bidirectional
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 ram_data_io[8]
port 39 nsew signal bidirectional
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 ram_data_io[9]
port 40 nsew signal bidirectional
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 ram_rw_en_o
port 41 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 reset_i
port 42 nsew signal input
flabel metal2 s 15474 31200 15530 32000 0 FreeSans 224 90 0 0 stop_lamp_o
port 43 nsew signal tristate
rlabel metal1 15962 29376 15962 29376 0 VGND
rlabel metal1 15962 28832 15962 28832 0 VPWR
rlabel metal1 18763 23766 18763 23766 0 _0000_
rlabel metal2 23046 11934 23046 11934 0 _0001_
rlabel metal1 21305 12206 21305 12206 0 _0002_
rlabel metal2 20194 15640 20194 15640 0 _0003_
rlabel metal1 24564 16150 24564 16150 0 _0004_
rlabel metal2 25438 16354 25438 16354 0 _0005_
rlabel metal2 24886 18088 24886 18088 0 _0006_
rlabel metal2 24978 19822 24978 19822 0 _0007_
rlabel metal2 25438 23528 25438 23528 0 _0008_
rlabel metal1 23552 23494 23552 23494 0 _0009_
rlabel metal1 22087 23018 22087 23018 0 _0010_
rlabel metal1 18124 22202 18124 22202 0 _0011_
rlabel metal2 17066 17442 17066 17442 0 _0012_
rlabel metal1 16698 21318 16698 21318 0 _0013_
rlabel metal1 13945 18666 13945 18666 0 _0014_
rlabel metal1 8648 18938 8648 18938 0 _0015_
rlabel metal2 6118 18530 6118 18530 0 _0016_
rlabel metal2 3542 18462 3542 18462 0 _0017_
rlabel metal2 3910 20230 3910 20230 0 _0018_
rlabel metal2 17066 15640 17066 15640 0 _0019_
rlabel metal1 15831 16150 15831 16150 0 _0020_
rlabel metal1 14628 16762 14628 16762 0 _0021_
rlabel metal1 14497 24786 14497 24786 0 _0022_
rlabel metal2 15594 23970 15594 23970 0 _0023_
rlabel metal1 15732 22950 15732 22950 0 _0024_
rlabel metal1 15647 20502 15647 20502 0 _0025_
rlabel metal1 12151 24106 12151 24106 0 _0026_
rlabel metal1 11868 24922 11868 24922 0 _0027_
rlabel metal2 9430 24990 9430 24990 0 _0028_
rlabel metal1 5796 23834 5796 23834 0 _0029_
rlabel metal2 8418 24582 8418 24582 0 _0030_
rlabel metal1 11224 15334 11224 15334 0 _0031_
rlabel metal1 10955 16490 10955 16490 0 _0032_
rlabel metal2 4554 17442 4554 17442 0 _0033_
rlabel metal1 3726 16014 3726 16014 0 _0034_
rlabel metal1 3128 14042 3128 14042 0 _0035_
rlabel metal2 3266 12036 3266 12036 0 _0036_
rlabel metal1 3220 10778 3220 10778 0 _0037_
rlabel metal1 3542 9146 3542 9146 0 _0038_
rlabel metal2 4186 7582 4186 7582 0 _0039_
rlabel metal2 6762 6120 6762 6120 0 _0040_
rlabel metal1 11592 5338 11592 5338 0 _0041_
rlabel metal1 17809 5610 17809 5610 0 _0042_
rlabel metal2 16790 8058 16790 8058 0 _0043_
rlabel metal1 19097 9962 19097 9962 0 _0044_
rlabel metal2 12190 13056 12190 13056 0 _0045_
rlabel metal2 12466 11560 12466 11560 0 _0046_
rlabel metal1 20240 5882 20240 5882 0 _0047_
rlabel metal1 22540 5882 22540 5882 0 _0048_
rlabel metal1 24012 5882 24012 5882 0 _0049_
rlabel metal2 21942 11968 21942 11968 0 _0050_
rlabel metal1 20056 11866 20056 11866 0 _0051_
rlabel metal1 19448 15674 19448 15674 0 _0052_
rlabel metal2 23230 16626 23230 16626 0 _0053_
rlabel metal1 24978 16218 24978 16218 0 _0054_
rlabel metal1 24242 18360 24242 18360 0 _0055_
rlabel metal1 24334 19448 24334 19448 0 _0056_
rlabel metal1 24932 23290 24932 23290 0 _0057_
rlabel metal1 22908 22746 22908 22746 0 _0058_
rlabel metal1 20608 23018 20608 23018 0 _0059_
rlabel metal2 16974 22372 16974 22372 0 _0060_
rlabel metal1 16560 17714 16560 17714 0 _0061_
rlabel metal1 16100 20570 16100 20570 0 _0062_
rlabel metal1 12374 18802 12374 18802 0 _0063_
rlabel metal1 7912 19414 7912 19414 0 _0064_
rlabel metal1 5382 18632 5382 18632 0 _0065_
rlabel metal1 3082 18326 3082 18326 0 _0066_
rlabel metal1 2944 20026 2944 20026 0 _0067_
rlabel metal1 16192 15130 16192 15130 0 _0068_
rlabel metal1 14628 16014 14628 16014 0 _0069_
rlabel metal1 13984 16762 13984 16762 0 _0070_
rlabel metal1 19232 25194 19232 25194 0 _0071_
rlabel metal1 14950 21114 14950 21114 0 _0072_
rlabel metal1 17424 26350 17424 26350 0 _0073_
rlabel metal2 12834 25670 12834 25670 0 _0074_
rlabel metal1 14459 25942 14459 25942 0 _0075_
rlabel metal1 15267 25874 15267 25874 0 _0076_
rlabel metal1 10626 23834 10626 23834 0 _0077_
rlabel metal2 10994 25058 10994 25058 0 _0078_
rlabel metal1 9798 24378 9798 24378 0 _0079_
rlabel metal1 6302 23834 6302 23834 0 _0080_
rlabel metal1 6624 24378 6624 24378 0 _0081_
rlabel metal1 10987 14586 10987 14586 0 _0082_
rlabel metal1 9338 16490 9338 16490 0 _0083_
rlabel metal1 4140 17306 4140 17306 0 _0084_
rlabel metal1 2438 15674 2438 15674 0 _0085_
rlabel metal1 2300 14042 2300 14042 0 _0086_
rlabel metal1 2392 12274 2392 12274 0 _0087_
rlabel metal1 2392 10778 2392 10778 0 _0088_
rlabel metal2 2622 9316 2622 9316 0 _0089_
rlabel metal1 3772 7446 3772 7446 0 _0090_
rlabel metal1 6065 5882 6065 5882 0 _0091_
rlabel metal1 11178 5746 11178 5746 0 _0092_
rlabel metal2 16330 5916 16330 5916 0 _0093_
rlabel metal1 15548 7786 15548 7786 0 _0094_
rlabel metal1 17572 9962 17572 9962 0 _0095_
rlabel metal1 11546 12954 11546 12954 0 _0096_
rlabel metal1 11592 11662 11592 11662 0 _0097_
rlabel metal2 19458 6052 19458 6052 0 _0098_
rlabel metal1 21574 6188 21574 6188 0 _0099_
rlabel metal1 23966 6392 23966 6392 0 _0100_
rlabel metal2 19458 15164 19458 15164 0 _0101_
rlabel metal1 13708 21522 13708 21522 0 _0102_
rlabel metal1 14674 20842 14674 20842 0 _0103_
rlabel metal1 13340 19414 13340 19414 0 _0104_
rlabel metal1 18630 15470 18630 15470 0 _0105_
rlabel metal1 21666 14994 21666 14994 0 _0106_
rlabel metal1 25668 7990 25668 7990 0 _0107_
rlabel metal1 23782 8534 23782 8534 0 _0108_
rlabel metal1 9200 10030 9200 10030 0 _0109_
rlabel metal1 8970 10064 8970 10064 0 _0110_
rlabel metal1 9660 9962 9660 9962 0 _0111_
rlabel metal1 10258 10574 10258 10574 0 _0112_
rlabel metal2 8326 10880 8326 10880 0 _0113_
rlabel metal1 6854 12614 6854 12614 0 _0114_
rlabel metal1 7038 12138 7038 12138 0 _0115_
rlabel metal1 7958 12172 7958 12172 0 _0116_
rlabel metal1 6394 15130 6394 15130 0 _0117_
rlabel metal1 7866 20468 7866 20468 0 _0118_
rlabel metal2 6578 16252 6578 16252 0 _0119_
rlabel metal1 6210 16048 6210 16048 0 _0120_
rlabel metal2 7498 15130 7498 15130 0 _0121_
rlabel metal1 6670 17850 6670 17850 0 _0122_
rlabel metal2 6854 17476 6854 17476 0 _0123_
rlabel metal1 7130 17612 7130 17612 0 _0124_
rlabel metal1 11362 17646 11362 17646 0 _0125_
rlabel metal1 11868 17646 11868 17646 0 _0126_
rlabel metal2 11086 17952 11086 17952 0 _0127_
rlabel metal1 7222 17748 7222 17748 0 _0128_
rlabel metal1 5980 15674 5980 15674 0 _0129_
rlabel metal2 6946 16422 6946 16422 0 _0130_
rlabel metal2 7406 15708 7406 15708 0 _0131_
rlabel metal1 8050 13838 8050 13838 0 _0132_
rlabel metal2 7590 13396 7590 13396 0 _0133_
rlabel metal1 7866 13260 7866 13260 0 _0134_
rlabel metal1 8234 10608 8234 10608 0 _0135_
rlabel metal2 9154 10948 9154 10948 0 _0136_
rlabel metal1 9568 10642 9568 10642 0 _0137_
rlabel metal1 8970 10540 8970 10540 0 _0138_
rlabel metal1 8234 10778 8234 10778 0 _0139_
rlabel metal1 12972 10030 12972 10030 0 _0140_
rlabel metal1 14352 12206 14352 12206 0 _0141_
rlabel metal1 15226 13294 15226 13294 0 _0142_
rlabel metal1 14674 10676 14674 10676 0 _0143_
rlabel metal1 12834 9588 12834 9588 0 _0144_
rlabel metal1 14490 10234 14490 10234 0 _0145_
rlabel metal1 15640 11322 15640 11322 0 _0146_
rlabel metal1 15042 10506 15042 10506 0 _0147_
rlabel metal2 14858 10506 14858 10506 0 _0148_
rlabel metal1 13478 10200 13478 10200 0 _0149_
rlabel metal2 14858 5372 14858 5372 0 _0150_
rlabel metal1 12604 5338 12604 5338 0 _0151_
rlabel metal2 13662 7582 13662 7582 0 _0152_
rlabel metal1 7866 7888 7866 7888 0 _0153_
rlabel metal1 7544 7854 7544 7854 0 _0154_
rlabel metal1 7682 8058 7682 8058 0 _0155_
rlabel metal1 9936 6766 9936 6766 0 _0156_
rlabel metal1 9706 6834 9706 6834 0 _0157_
rlabel metal1 10488 7854 10488 7854 0 _0158_
rlabel metal2 12466 8262 12466 8262 0 _0159_
rlabel metal2 12558 9248 12558 9248 0 _0160_
rlabel metal1 13892 10642 13892 10642 0 _0161_
rlabel metal1 14628 12954 14628 12954 0 _0162_
rlabel metal2 14950 9588 14950 9588 0 _0163_
rlabel metal1 13892 10710 13892 10710 0 _0164_
rlabel metal1 14076 6834 14076 6834 0 _0165_
rlabel metal2 13754 6596 13754 6596 0 _0166_
rlabel metal1 14582 5746 14582 5746 0 _0167_
rlabel metal1 14030 6766 14030 6766 0 _0168_
rlabel metal2 13386 9027 13386 9027 0 _0169_
rlabel metal1 13616 10234 13616 10234 0 _0170_
rlabel metal1 13432 10642 13432 10642 0 _0171_
rlabel metal1 12558 10064 12558 10064 0 _0172_
rlabel metal1 19550 10098 19550 10098 0 _0173_
rlabel metal1 20884 9010 20884 9010 0 _0174_
rlabel metal1 25208 9146 25208 9146 0 _0175_
rlabel metal1 26082 8874 26082 8874 0 _0176_
rlabel metal1 25254 7786 25254 7786 0 _0177_
rlabel metal1 26174 8466 26174 8466 0 _0178_
rlabel viali 25622 8465 25622 8465 0 _0179_
rlabel metal2 24794 9384 24794 9384 0 _0180_
rlabel metal1 26036 9554 26036 9554 0 _0181_
rlabel metal1 25438 9588 25438 9588 0 _0182_
rlabel metal1 24472 9554 24472 9554 0 _0183_
rlabel metal1 9798 13906 9798 13906 0 _0184_
rlabel metal1 9384 12614 9384 12614 0 _0185_
rlabel metal1 13018 6800 13018 6800 0 _0186_
rlabel metal2 16054 8262 16054 8262 0 _0187_
rlabel metal1 17802 12920 17802 12920 0 _0188_
rlabel metal1 17802 11628 17802 11628 0 _0189_
rlabel metal1 17434 11832 17434 11832 0 _0190_
rlabel metal1 22494 8942 22494 8942 0 _0191_
rlabel metal1 22816 9486 22816 9486 0 _0192_
rlabel metal1 23506 9520 23506 9520 0 _0193_
rlabel metal2 18814 14756 18814 14756 0 _0194_
rlabel metal1 16790 14858 16790 14858 0 _0195_
rlabel metal1 17066 12784 17066 12784 0 _0196_
rlabel metal1 23736 7514 23736 7514 0 _0197_
rlabel metal1 14076 14994 14076 14994 0 _0198_
rlabel metal1 20838 7242 20838 7242 0 _0199_
rlabel metal1 23598 6766 23598 6766 0 _0200_
rlabel metal1 22678 9622 22678 9622 0 _0201_
rlabel metal1 26220 9146 26220 9146 0 _0202_
rlabel metal1 24886 9418 24886 9418 0 _0203_
rlabel via2 8694 13821 8694 13821 0 _0204_
rlabel metal1 23000 6766 23000 6766 0 _0205_
rlabel metal2 21390 6460 21390 6460 0 _0206_
rlabel viali 20653 10030 20653 10030 0 _0207_
rlabel metal1 20217 9962 20217 9962 0 _0208_
rlabel metal2 20654 8704 20654 8704 0 _0209_
rlabel metal1 19780 5678 19780 5678 0 _0210_
rlabel metal1 17204 12682 17204 12682 0 _0211_
rlabel metal1 17250 11730 17250 11730 0 _0212_
rlabel metal1 15088 12750 15088 12750 0 _0213_
rlabel metal1 12834 9350 12834 9350 0 _0214_
rlabel metal2 12650 10166 12650 10166 0 _0215_
rlabel metal2 15134 10676 15134 10676 0 _0216_
rlabel metal2 15226 13090 15226 13090 0 _0217_
rlabel metal1 15272 12274 15272 12274 0 _0218_
rlabel metal1 16031 11798 16031 11798 0 _0219_
rlabel metal1 12650 11220 12650 11220 0 _0220_
rlabel metal1 11684 11254 11684 11254 0 _0221_
rlabel metal1 16882 12886 16882 12886 0 _0222_
rlabel metal1 17079 12886 17079 12886 0 _0223_
rlabel metal2 16698 13124 16698 13124 0 _0224_
rlabel metal2 13110 13056 13110 13056 0 _0225_
rlabel metal2 17158 10030 17158 10030 0 _0226_
rlabel metal1 15272 10098 15272 10098 0 _0227_
rlabel metal1 17033 9622 17033 9622 0 _0228_
rlabel metal1 18032 15130 18032 15130 0 _0229_
rlabel metal1 16882 9690 16882 9690 0 _0230_
rlabel metal1 17296 10234 17296 10234 0 _0231_
rlabel metal1 15410 7344 15410 7344 0 _0232_
rlabel metal1 15548 7174 15548 7174 0 _0233_
rlabel metal2 15962 7990 15962 7990 0 _0234_
rlabel metal1 13110 9010 13110 9010 0 _0235_
rlabel metal1 15883 8534 15883 8534 0 _0236_
rlabel metal1 15594 8466 15594 8466 0 _0237_
rlabel metal1 15088 8602 15088 8602 0 _0238_
rlabel metal1 18078 19278 18078 19278 0 _0239_
rlabel metal1 15502 6426 15502 6426 0 _0240_
rlabel metal1 14214 5338 14214 5338 0 _0241_
rlabel metal1 10580 8330 10580 8330 0 _0242_
rlabel metal1 13478 5746 13478 5746 0 _0243_
rlabel metal2 14766 5338 14766 5338 0 _0244_
rlabel metal2 15226 6086 15226 6086 0 _0245_
rlabel metal1 15778 6766 15778 6766 0 _0246_
rlabel metal1 16238 6290 16238 6290 0 _0247_
rlabel metal2 13110 7174 13110 7174 0 _0248_
rlabel metal1 13110 5882 13110 5882 0 _0249_
rlabel metal2 12926 6970 12926 6970 0 _0250_
rlabel metal2 5290 16932 5290 16932 0 _0251_
rlabel metal1 11638 6290 11638 6290 0 _0252_
rlabel metal1 9660 9146 9660 9146 0 _0253_
rlabel metal1 8602 8058 8602 8058 0 _0254_
rlabel metal1 8510 7446 8510 7446 0 _0255_
rlabel metal1 10580 7922 10580 7922 0 _0256_
rlabel metal1 9453 7446 9453 7446 0 _0257_
rlabel metal1 7912 6766 7912 6766 0 _0258_
rlabel metal1 6486 6732 6486 6732 0 _0259_
rlabel metal2 8142 8228 8142 8228 0 _0260_
rlabel via2 13754 15453 13754 15453 0 _0261_
rlabel metal1 8444 8568 8444 8568 0 _0262_
rlabel metal1 8510 8398 8510 8398 0 _0263_
rlabel metal1 5612 7718 5612 7718 0 _0264_
rlabel metal1 4002 7820 4002 7820 0 _0265_
rlabel metal1 9798 9486 9798 9486 0 _0266_
rlabel metal1 10166 10676 10166 10676 0 _0267_
rlabel metal2 10074 10285 10074 10285 0 _0268_
rlabel metal1 10074 10098 10074 10098 0 _0269_
rlabel metal2 10626 9724 10626 9724 0 _0270_
rlabel metal1 10488 9486 10488 9486 0 _0271_
rlabel metal1 7222 9350 7222 9350 0 _0272_
rlabel metal1 3082 8976 3082 8976 0 _0273_
rlabel metal1 10902 11152 10902 11152 0 _0274_
rlabel metal1 9936 12886 9936 12886 0 _0275_
rlabel metal1 9430 12954 9430 12954 0 _0276_
rlabel metal1 9852 11866 9852 11866 0 _0277_
rlabel metal1 10396 11118 10396 11118 0 _0278_
rlabel metal1 4462 11118 4462 11118 0 _0279_
rlabel metal1 2898 10676 2898 10676 0 _0280_
rlabel metal1 9200 12818 9200 12818 0 _0281_
rlabel metal1 7958 14042 7958 14042 0 _0282_
rlabel via1 7958 13821 7958 13821 0 _0283_
rlabel metal2 7866 12716 7866 12716 0 _0284_
rlabel metal1 8533 12818 8533 12818 0 _0285_
rlabel metal1 5520 12070 5520 12070 0 _0286_
rlabel metal1 3312 12410 3312 12410 0 _0287_
rlabel metal1 8510 13974 8510 13974 0 _0288_
rlabel metal1 9414 13974 9414 13974 0 _0289_
rlabel metal1 8786 13906 8786 13906 0 _0290_
rlabel metal1 8326 14008 8326 14008 0 _0291_
rlabel metal1 2691 13906 2691 13906 0 _0292_
rlabel metal1 9522 18190 9522 18190 0 _0293_
rlabel metal1 8556 17578 8556 17578 0 _0294_
rlabel metal2 8142 16252 8142 16252 0 _0295_
rlabel metal2 7038 17340 7038 17340 0 _0296_
rlabel via1 8431 16082 8431 16082 0 _0297_
rlabel metal1 6854 15946 6854 15946 0 _0298_
rlabel metal2 2714 15946 2714 15946 0 _0299_
rlabel metal1 8050 17578 8050 17578 0 _0300_
rlabel viali 8339 17646 8339 17646 0 _0301_
rlabel metal1 6532 17238 6532 17238 0 _0302_
rlabel metal1 4370 17204 4370 17204 0 _0303_
rlabel metal1 9614 18292 9614 18292 0 _0304_
rlabel metal2 11454 18054 11454 18054 0 _0305_
rlabel metal1 11224 18122 11224 18122 0 _0306_
rlabel metal1 9660 17306 9660 17306 0 _0307_
rlabel metal1 9016 16558 9016 16558 0 _0308_
rlabel metal2 11914 14790 11914 14790 0 _0309_
rlabel metal1 12949 15062 12949 15062 0 _0310_
rlabel metal1 13156 22610 13156 22610 0 _0311_
rlabel metal2 12466 20179 12466 20179 0 _0312_
rlabel metal1 14766 20978 14766 20978 0 _0313_
rlabel metal1 13110 20400 13110 20400 0 _0314_
rlabel metal1 8142 23222 8142 23222 0 _0315_
rlabel metal2 12282 22848 12282 22848 0 _0316_
rlabel metal1 10718 23698 10718 23698 0 _0317_
rlabel metal2 6716 20910 6716 20910 0 _0318_
rlabel metal1 9246 19788 9246 19788 0 _0319_
rlabel metal1 11316 20434 11316 20434 0 _0320_
rlabel metal2 11822 22542 11822 22542 0 _0321_
rlabel metal2 10994 20706 10994 20706 0 _0322_
rlabel metal1 7498 20978 7498 20978 0 _0323_
rlabel metal1 7406 20502 7406 20502 0 _0324_
rlabel metal1 5789 20910 5789 20910 0 _0325_
rlabel metal1 4830 21658 4830 21658 0 _0326_
rlabel metal2 4186 22372 4186 22372 0 _0327_
rlabel metal1 4692 22066 4692 22066 0 _0328_
rlabel metal1 5014 22542 5014 22542 0 _0329_
rlabel metal1 4968 22202 4968 22202 0 _0330_
rlabel metal1 19228 16694 19228 16694 0 _0331_
rlabel metal1 6256 21522 6256 21522 0 _0332_
rlabel metal1 7314 22644 7314 22644 0 _0333_
rlabel metal1 8211 22474 8211 22474 0 _0334_
rlabel metal1 7452 23018 7452 23018 0 _0335_
rlabel metal1 7728 22746 7728 22746 0 _0336_
rlabel metal1 9384 21998 9384 21998 0 _0337_
rlabel metal1 10028 21046 10028 21046 0 _0338_
rlabel metal1 8556 20910 8556 20910 0 _0339_
rlabel metal1 8878 23018 8878 23018 0 _0340_
rlabel metal1 8326 22950 8326 22950 0 _0341_
rlabel metal2 7498 22678 7498 22678 0 _0342_
rlabel metal1 6348 22202 6348 22202 0 _0343_
rlabel metal1 7071 22542 7071 22542 0 _0344_
rlabel metal1 6302 22678 6302 22678 0 _0345_
rlabel metal1 7682 22542 7682 22542 0 _0346_
rlabel metal1 7038 22746 7038 22746 0 _0347_
rlabel metal1 5244 20978 5244 20978 0 _0348_
rlabel metal1 6164 21114 6164 21114 0 _0349_
rlabel metal1 7038 21658 7038 21658 0 _0350_
rlabel metal1 6486 23290 6486 23290 0 _0351_
rlabel metal1 6762 23800 6762 23800 0 _0352_
rlabel metal1 8832 22202 8832 22202 0 _0353_
rlabel metal1 7360 20434 7360 20434 0 _0354_
rlabel metal2 7590 20774 7590 20774 0 _0355_
rlabel metal1 8050 20910 8050 20910 0 _0356_
rlabel metal1 8418 20944 8418 20944 0 _0357_
rlabel metal1 8326 21114 8326 21114 0 _0358_
rlabel metal1 9108 22746 9108 22746 0 _0359_
rlabel metal1 10534 20944 10534 20944 0 _0360_
rlabel metal2 10534 21318 10534 21318 0 _0361_
rlabel metal2 11546 20740 11546 20740 0 _0362_
rlabel metal2 11178 20434 11178 20434 0 _0363_
rlabel metal1 10764 21114 10764 21114 0 _0364_
rlabel metal1 10396 21658 10396 21658 0 _0365_
rlabel metal1 10810 22066 10810 22066 0 _0366_
rlabel metal1 11270 22644 11270 22644 0 _0367_
rlabel metal1 11684 22202 11684 22202 0 _0368_
rlabel metal1 11454 22610 11454 22610 0 _0369_
rlabel metal2 10810 23256 10810 23256 0 _0370_
rlabel metal2 13846 21148 13846 21148 0 _0371_
rlabel metal1 7038 19210 7038 19210 0 _0372_
rlabel metal1 14122 14858 14122 14858 0 _0373_
rlabel metal1 14950 15674 14950 15674 0 _0374_
rlabel metal1 15916 14994 15916 14994 0 _0375_
rlabel metal1 3266 19856 3266 19856 0 _0376_
rlabel metal1 3358 18700 3358 18700 0 _0377_
rlabel metal1 6072 19346 6072 19346 0 _0378_
rlabel metal1 9430 19278 9430 19278 0 _0379_
rlabel metal1 12144 18394 12144 18394 0 _0380_
rlabel metal1 17480 18734 17480 18734 0 _0381_
rlabel metal1 18630 20876 18630 20876 0 _0382_
rlabel metal2 30130 18836 30130 18836 0 _0383_
rlabel metal2 30038 18054 30038 18054 0 _0384_
rlabel metal1 29164 18666 29164 18666 0 _0385_
rlabel metal1 23736 13974 23736 13974 0 _0386_
rlabel metal1 23138 13872 23138 13872 0 _0387_
rlabel metal1 25070 13294 25070 13294 0 _0388_
rlabel metal2 24702 12988 24702 12988 0 _0389_
rlabel metal1 25898 13498 25898 13498 0 _0390_
rlabel metal1 25576 14586 25576 14586 0 _0391_
rlabel metal1 25668 15130 25668 15130 0 _0392_
rlabel metal1 26036 14246 26036 14246 0 _0393_
rlabel metal2 27738 14688 27738 14688 0 _0394_
rlabel metal1 28106 14382 28106 14382 0 _0395_
rlabel metal2 25898 14756 25898 14756 0 _0396_
rlabel metal2 26542 13566 26542 13566 0 _0397_
rlabel metal1 25622 11050 25622 11050 0 _0398_
rlabel metal1 25070 10778 25070 10778 0 _0399_
rlabel metal1 25898 12852 25898 12852 0 _0400_
rlabel metal1 24794 14314 24794 14314 0 _0401_
rlabel metal1 24288 10642 24288 10642 0 _0402_
rlabel metal1 24564 9962 24564 9962 0 _0403_
rlabel metal1 24564 10778 24564 10778 0 _0404_
rlabel metal1 25254 12750 25254 12750 0 _0405_
rlabel metal2 25622 13668 25622 13668 0 _0406_
rlabel metal1 26496 14450 26496 14450 0 _0407_
rlabel metal2 26358 13770 26358 13770 0 _0408_
rlabel metal1 28566 18700 28566 18700 0 _0409_
rlabel metal2 29486 20230 29486 20230 0 _0410_
rlabel metal1 28474 20434 28474 20434 0 _0411_
rlabel metal1 29762 19958 29762 19958 0 _0412_
rlabel metal1 28934 22576 28934 22576 0 _0413_
rlabel metal1 27416 22610 27416 22610 0 _0414_
rlabel metal1 29532 21998 29532 21998 0 _0415_
rlabel metal1 29026 22474 29026 22474 0 _0416_
rlabel metal1 29394 22644 29394 22644 0 _0417_
rlabel metal2 29302 22168 29302 22168 0 _0418_
rlabel metal1 29026 20910 29026 20910 0 _0419_
rlabel metal1 25254 21114 25254 21114 0 _0420_
rlabel via1 28934 20230 28934 20230 0 _0421_
rlabel metal1 28428 20910 28428 20910 0 _0422_
rlabel metal1 23690 20978 23690 20978 0 _0423_
rlabel metal1 22494 20808 22494 20808 0 _0424_
rlabel metal1 22954 20876 22954 20876 0 _0425_
rlabel metal2 18722 21556 18722 21556 0 _0426_
rlabel metal2 18814 20638 18814 20638 0 _0427_
rlabel metal1 18906 20944 18906 20944 0 _0428_
rlabel metal2 19090 19142 19090 19142 0 _0429_
rlabel metal2 19458 19652 19458 19652 0 _0430_
rlabel metal1 19412 20502 19412 20502 0 _0431_
rlabel metal1 17572 20026 17572 20026 0 _0432_
rlabel metal1 17112 19754 17112 19754 0 _0433_
rlabel metal1 16790 19890 16790 19890 0 _0434_
rlabel metal2 17618 19108 17618 19108 0 _0435_
rlabel metal1 17480 19346 17480 19346 0 _0436_
rlabel metal1 21482 10438 21482 10438 0 _0437_
rlabel metal1 22310 11186 22310 11186 0 _0438_
rlabel metal1 23184 15674 23184 15674 0 _0439_
rlabel metal2 26450 18326 26450 18326 0 _0440_
rlabel metal2 26266 21811 26266 21811 0 _0441_
rlabel via1 20470 21301 20470 21301 0 _0442_
rlabel metal2 18170 19108 18170 19108 0 _0443_
rlabel metal1 16560 18938 16560 18938 0 _0444_
rlabel metal2 17434 19890 17434 19890 0 _0445_
rlabel metal1 17848 22066 17848 22066 0 _0446_
rlabel metal1 16560 20434 16560 20434 0 _0447_
rlabel metal1 18078 19380 18078 19380 0 _0448_
rlabel metal1 18216 18938 18216 18938 0 _0449_
rlabel metal1 19228 20434 19228 20434 0 _0450_
rlabel metal1 18952 19278 18952 19278 0 _0451_
rlabel metal1 17802 17306 17802 17306 0 _0452_
rlabel metal2 17250 17782 17250 17782 0 _0453_
rlabel metal1 21390 21862 21390 21862 0 _0454_
rlabel metal1 17710 21556 17710 21556 0 _0455_
rlabel metal1 19596 21998 19596 21998 0 _0456_
rlabel metal1 19136 22202 19136 22202 0 _0457_
rlabel metal1 20102 21624 20102 21624 0 _0458_
rlabel metal1 18331 21590 18331 21590 0 _0459_
rlabel metal1 17618 21658 17618 21658 0 _0460_
rlabel metal1 17204 21998 17204 21998 0 _0461_
rlabel metal1 21666 22032 21666 22032 0 _0462_
rlabel metal1 23368 21114 23368 21114 0 _0463_
rlabel metal1 22816 21658 22816 21658 0 _0464_
rlabel metal1 21344 22202 21344 22202 0 _0465_
rlabel metal1 20792 22746 20792 22746 0 _0466_
rlabel metal1 27048 21114 27048 21114 0 _0467_
rlabel metal1 26174 21930 26174 21930 0 _0468_
rlabel metal1 28612 18870 28612 18870 0 _0469_
rlabel metal1 28612 20570 28612 20570 0 _0470_
rlabel metal1 29302 22066 29302 22066 0 _0471_
rlabel metal1 27255 21930 27255 21930 0 _0472_
rlabel metal1 25530 22202 25530 22202 0 _0473_
rlabel metal1 23414 22610 23414 22610 0 _0474_
rlabel metal1 28106 20910 28106 20910 0 _0475_
rlabel metal1 27148 20774 27148 20774 0 _0476_
rlabel metal1 27646 21012 27646 21012 0 _0477_
rlabel metal1 27830 21114 27830 21114 0 _0478_
rlabel metal2 25162 22916 25162 22916 0 _0479_
rlabel metal1 27968 17646 27968 17646 0 _0480_
rlabel metal1 27508 17850 27508 17850 0 _0481_
rlabel metal2 26358 19142 26358 19142 0 _0482_
rlabel metal1 30084 19278 30084 19278 0 _0483_
rlabel metal1 28796 19482 28796 19482 0 _0484_
rlabel metal1 25714 19482 25714 19482 0 _0485_
rlabel metal1 24748 19822 24748 19822 0 _0486_
rlabel metal1 28336 18802 28336 18802 0 _0487_
rlabel metal1 28152 17850 28152 17850 0 _0488_
rlabel metal2 28474 18564 28474 18564 0 _0489_
rlabel metal2 26266 18496 26266 18496 0 _0490_
rlabel metal1 25208 18394 25208 18394 0 _0491_
rlabel metal1 25438 12852 25438 12852 0 _0492_
rlabel metal1 24472 12818 24472 12818 0 _0493_
rlabel metal2 24058 13838 24058 13838 0 _0494_
rlabel metal1 24380 14586 24380 14586 0 _0495_
rlabel metal1 25944 14858 25944 14858 0 _0496_
rlabel metal1 26404 15130 26404 15130 0 _0497_
rlabel metal1 27370 15504 27370 15504 0 _0498_
rlabel metal1 26818 15538 26818 15538 0 _0499_
rlabel metal1 26220 15674 26220 15674 0 _0500_
rlabel metal1 25254 16116 25254 16116 0 _0501_
rlabel metal1 23460 14042 23460 14042 0 _0502_
rlabel metal1 23736 14518 23736 14518 0 _0503_
rlabel metal1 21436 14586 21436 14586 0 _0504_
rlabel metal1 21298 14892 21298 14892 0 _0505_
rlabel metal1 23284 15402 23284 15402 0 _0506_
rlabel metal1 23552 15470 23552 15470 0 _0507_
rlabel metal1 24058 15674 24058 15674 0 _0508_
rlabel metal1 23276 16082 23276 16082 0 _0509_
rlabel metal1 21114 14926 21114 14926 0 _0510_
rlabel metal1 24518 13226 24518 13226 0 _0511_
rlabel metal1 24196 13498 24196 13498 0 _0512_
rlabel metal1 20562 14994 20562 14994 0 _0513_
rlabel metal2 19734 15232 19734 15232 0 _0514_
rlabel metal1 23782 12954 23782 12954 0 _0515_
rlabel viali 21521 14348 21521 14348 0 _0516_
rlabel metal2 22218 13804 22218 13804 0 _0517_
rlabel metal1 22218 13158 22218 13158 0 _0518_
rlabel metal1 20976 13158 20976 13158 0 _0519_
rlabel metal1 22310 10778 22310 10778 0 _0520_
rlabel metal1 25254 10234 25254 10234 0 _0521_
rlabel metal1 23253 11050 23253 11050 0 _0522_
rlabel metal1 21620 11322 21620 11322 0 _0523_
rlabel metal1 21712 11866 21712 11866 0 _0524_
rlabel metal1 15134 21522 15134 21522 0 _0525_
rlabel metal1 19780 19346 19780 19346 0 _0526_
rlabel metal1 12650 9554 12650 9554 0 _0527_
rlabel metal1 11592 15402 11592 15402 0 _0528_
rlabel metal1 4830 8976 4830 8976 0 _0529_
rlabel metal2 5152 9554 5152 9554 0 _0530_
rlabel metal1 18630 13974 18630 13974 0 _0531_
rlabel metal2 19182 14110 19182 14110 0 _0532_
rlabel metal2 19274 14178 19274 14178 0 _0533_
rlabel metal1 18676 13294 18676 13294 0 _0534_
rlabel metal1 19826 17170 19826 17170 0 _0535_
rlabel metal1 20838 18224 20838 18224 0 _0536_
rlabel metal2 20930 17714 20930 17714 0 _0537_
rlabel metal1 20930 19822 20930 19822 0 _0538_
rlabel metal2 15226 25738 15226 25738 0 _0539_
rlabel metal1 14444 23834 14444 23834 0 _0540_
rlabel metal1 15272 21658 15272 21658 0 _0541_
rlabel metal2 15686 22644 15686 22644 0 _0542_
rlabel metal1 19044 24378 19044 24378 0 _0543_
rlabel metal1 16422 23698 16422 23698 0 _0544_
rlabel metal2 12558 20944 12558 20944 0 _0545_
rlabel metal2 12742 20026 12742 20026 0 _0546_
rlabel metal1 16882 8500 16882 8500 0 _0547_
rlabel metal1 21666 12784 21666 12784 0 _0548_
rlabel metal1 16744 21522 16744 21522 0 _0549_
rlabel metal1 15916 20434 15916 20434 0 _0550_
rlabel metal1 19228 25806 19228 25806 0 _0551_
rlabel metal1 16974 26928 16974 26928 0 _0552_
rlabel metal2 14582 26486 14582 26486 0 _0553_
rlabel metal1 15410 25466 15410 25466 0 _0554_
rlabel metal1 11086 16592 11086 16592 0 _0555_
rlabel metal1 12144 16490 12144 16490 0 _0556_
rlabel metal1 9752 14926 9752 14926 0 _0557_
rlabel metal1 6762 15368 6762 15368 0 _0558_
rlabel metal1 5152 14586 5152 14586 0 _0559_
rlabel metal1 4094 13770 4094 13770 0 _0560_
rlabel metal1 5014 12274 5014 12274 0 _0561_
rlabel metal1 4922 10642 4922 10642 0 _0562_
rlabel metal1 6256 9622 6256 9622 0 _0563_
rlabel metal2 5382 8126 5382 8126 0 _0564_
rlabel metal2 7682 7548 7682 7548 0 _0565_
rlabel metal2 12742 9231 12742 9231 0 _0566_
rlabel metal1 17710 6834 17710 6834 0 _0567_
rlabel metal1 17664 8534 17664 8534 0 _0568_
rlabel metal1 18354 11594 18354 11594 0 _0569_
rlabel metal1 16882 14008 16882 14008 0 _0570_
rlabel metal1 15502 14314 15502 14314 0 _0571_
rlabel metal1 19826 8058 19826 8058 0 _0572_
rlabel metal1 20102 6868 20102 6868 0 _0573_
rlabel metal1 19918 7378 19918 7378 0 _0574_
rlabel metal1 19918 10642 19918 10642 0 _0575_
rlabel metal1 19504 13362 19504 13362 0 _0576_
rlabel metal2 20654 17272 20654 17272 0 _0577_
rlabel metal1 23046 18054 23046 18054 0 _0578_
rlabel metal2 26542 17646 26542 17646 0 _0579_
rlabel metal1 24610 17714 24610 17714 0 _0580_
rlabel metal1 23644 19278 23644 19278 0 _0581_
rlabel metal1 23782 20026 23782 20026 0 _0582_
rlabel metal1 23644 20298 23644 20298 0 _0583_
rlabel metal2 21206 19584 21206 19584 0 _0584_
rlabel metal1 20010 20808 20010 20808 0 _0585_
rlabel metal1 19688 17578 19688 17578 0 _0586_
rlabel metal2 14490 18802 14490 18802 0 _0587_
rlabel metal1 18446 12886 18446 12886 0 clknet_0_clock
rlabel metal1 2346 9418 2346 9418 0 clknet_2_0__leaf_clock
rlabel metal1 2622 18258 2622 18258 0 clknet_2_1__leaf_clock
rlabel metal1 15732 7922 15732 7922 0 clknet_2_2__leaf_clock
rlabel metal1 16192 20978 16192 20978 0 clknet_2_3__leaf_clock
rlabel metal1 5520 16150 5520 16150 0 clock
rlabel metal1 18216 29274 18216 29274 0 logisim_clock_tree_0_out
rlabel metal1 13018 25398 13018 25398 0 manchester_baby_instance.BASE_0.s_countReg\[0\]
rlabel metal1 13616 26010 13616 26010 0 manchester_baby_instance.BASE_0.s_countReg\[1\]
rlabel metal2 16238 26180 16238 26180 0 manchester_baby_instance.BASE_0.s_countReg\[2\]
rlabel metal1 15870 26418 15870 26418 0 manchester_baby_instance.BASE_0.s_tickNext
rlabel metal1 18906 26010 18906 26010 0 manchester_baby_instance.BASE_0.s_tickReg
rlabel metal1 18722 24684 18722 24684 0 manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
rlabel metal1 18952 26418 18952 26418 0 manchester_baby_instance.BASE_1.s_counterValue
rlabel metal1 19044 25330 19044 25330 0 manchester_baby_instance.BASE_1.s_derivedClock
rlabel metal2 12006 23562 12006 23562 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
rlabel metal1 12328 24786 12328 24786 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
rlabel metal1 9706 22066 9706 22066 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
rlabel metal1 5750 21556 5750 21556 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
rlabel metal1 4094 22644 4094 22644 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
rlabel metal2 19458 21012 19458 21012 0 manchester_baby_instance.CIRCUIT_0.Acc.tick
rlabel metal1 14490 24242 14490 24242 0 manchester_baby_instance.CIRCUIT_0.GATES_13.result
rlabel metal1 13984 19278 13984 19278 0 manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
rlabel metal1 17894 16150 17894 16150 0 manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
rlabel metal1 15870 16014 15870 16014 0 manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
rlabel metal1 15410 17170 15410 17170 0 manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
rlabel metal1 9476 19890 9476 19890 0 manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
rlabel metal1 7452 19890 7452 19890 0 manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
rlabel metal2 5014 18836 5014 18836 0 manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
rlabel metal1 4692 20910 4692 20910 0 manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
rlabel metal1 13570 23766 13570 23766 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
rlabel metal1 14858 23732 14858 23732 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
rlabel metal1 15410 21454 15410 21454 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
rlabel metal1 12834 21964 12834 21964 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
rlabel metal1 14858 24072 14858 24072 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
rlabel metal1 14766 22712 14766 22712 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
rlabel metal2 13478 16320 13478 16320 0 manchester_baby_instance.ram_data_i_0
rlabel metal1 9154 18190 9154 18190 0 manchester_baby_instance.ram_data_i_1
rlabel metal1 13340 5610 13340 5610 0 manchester_baby_instance.ram_data_i_10
rlabel metal1 15686 6256 15686 6256 0 manchester_baby_instance.ram_data_i_11
rlabel metal1 16330 7378 16330 7378 0 manchester_baby_instance.ram_data_i_12
rlabel metal1 15686 15538 15686 15538 0 manchester_baby_instance.ram_data_i_13
rlabel metal1 14398 13838 14398 13838 0 manchester_baby_instance.ram_data_i_14
rlabel metal1 14352 13702 14352 13702 0 manchester_baby_instance.ram_data_i_15
rlabel metal1 21574 10064 21574 10064 0 manchester_baby_instance.ram_data_i_16
rlabel metal1 24978 7208 24978 7208 0 manchester_baby_instance.ram_data_i_17
rlabel metal1 22471 10574 22471 10574 0 manchester_baby_instance.ram_data_i_18
rlabel metal1 21735 10778 21735 10778 0 manchester_baby_instance.ram_data_i_19
rlabel metal1 8740 15674 8740 15674 0 manchester_baby_instance.ram_data_i_2
rlabel metal1 23276 13362 23276 13362 0 manchester_baby_instance.ram_data_i_20
rlabel metal1 21574 15504 21574 15504 0 manchester_baby_instance.ram_data_i_21
rlabel metal1 24978 15640 24978 15640 0 manchester_baby_instance.ram_data_i_22
rlabel metal1 27922 15946 27922 15946 0 manchester_baby_instance.ram_data_i_23
rlabel metal1 27922 17578 27922 17578 0 manchester_baby_instance.ram_data_i_24
rlabel metal1 27646 18700 27646 18700 0 manchester_baby_instance.ram_data_i_25
rlabel metal2 27968 22202 27968 22202 0 manchester_baby_instance.ram_data_i_26
rlabel metal1 27186 22542 27186 22542 0 manchester_baby_instance.ram_data_i_27
rlabel metal1 21344 21454 21344 21454 0 manchester_baby_instance.ram_data_i_28
rlabel metal1 19826 22508 19826 22508 0 manchester_baby_instance.ram_data_i_29
rlabel metal1 8510 16592 8510 16592 0 manchester_baby_instance.ram_data_i_3
rlabel metal2 18998 18360 18998 18360 0 manchester_baby_instance.ram_data_i_30
rlabel metal2 16238 19584 16238 19584 0 manchester_baby_instance.ram_data_i_31
rlabel metal1 4738 21964 4738 21964 0 manchester_baby_instance.ram_data_i_4
rlabel metal2 6118 12551 6118 12551 0 manchester_baby_instance.ram_data_i_5
rlabel metal1 8234 11322 8234 11322 0 manchester_baby_instance.ram_data_i_6
rlabel metal2 8602 9656 8602 9656 0 manchester_baby_instance.ram_data_i_7
rlabel metal2 7222 8262 7222 8262 0 manchester_baby_instance.ram_data_i_8
rlabel metal1 9430 7888 9430 7888 0 manchester_baby_instance.ram_data_i_9
rlabel metal1 13478 14416 13478 14416 0 manchester_baby_instance.ram_data_o_0
rlabel metal1 9660 17170 9660 17170 0 manchester_baby_instance.ram_data_o_1
rlabel metal1 13570 5814 13570 5814 0 manchester_baby_instance.ram_data_o_10
rlabel metal1 17250 6732 17250 6732 0 manchester_baby_instance.ram_data_o_11
rlabel metal2 17158 8228 17158 8228 0 manchester_baby_instance.ram_data_o_12
rlabel metal1 17986 9894 17986 9894 0 manchester_baby_instance.ram_data_o_13
rlabel metal1 14030 13974 14030 13974 0 manchester_baby_instance.ram_data_o_14
rlabel metal1 13478 12308 13478 12308 0 manchester_baby_instance.ram_data_o_15
rlabel metal1 21804 8466 21804 8466 0 manchester_baby_instance.ram_data_o_16
rlabel metal1 24886 7378 24886 7378 0 manchester_baby_instance.ram_data_o_17
rlabel metal1 24610 8330 24610 8330 0 manchester_baby_instance.ram_data_o_18
rlabel metal1 21298 11628 21298 11628 0 manchester_baby_instance.ram_data_o_19
rlabel metal1 5934 15028 5934 15028 0 manchester_baby_instance.ram_data_o_2
rlabel metal1 20516 13226 20516 13226 0 manchester_baby_instance.ram_data_o_20
rlabel metal2 21022 16150 21022 16150 0 manchester_baby_instance.ram_data_o_21
rlabel metal1 23690 17238 23690 17238 0 manchester_baby_instance.ram_data_o_22
rlabel metal1 27554 14994 27554 14994 0 manchester_baby_instance.ram_data_o_23
rlabel metal1 28750 17612 28750 17612 0 manchester_baby_instance.ram_data_o_24
rlabel metal1 28014 19822 28014 19822 0 manchester_baby_instance.ram_data_o_25
rlabel metal1 25208 20978 25208 20978 0 manchester_baby_instance.ram_data_o_26
rlabel metal1 23966 21590 23966 21590 0 manchester_baby_instance.ram_data_o_27
rlabel metal1 21482 20842 21482 20842 0 manchester_baby_instance.ram_data_o_28
rlabel metal1 19734 20978 19734 20978 0 manchester_baby_instance.ram_data_o_29
rlabel metal2 4186 16320 4186 16320 0 manchester_baby_instance.ram_data_o_3
rlabel metal1 18998 18802 18998 18802 0 manchester_baby_instance.ram_data_o_30
rlabel metal1 14306 19414 14306 19414 0 manchester_baby_instance.ram_data_o_31
rlabel metal1 3588 14586 3588 14586 0 manchester_baby_instance.ram_data_o_4
rlabel metal1 6118 12886 6118 12886 0 manchester_baby_instance.ram_data_o_5
rlabel metal1 6670 11050 6670 11050 0 manchester_baby_instance.ram_data_o_6
rlabel metal1 8510 9486 8510 9486 0 manchester_baby_instance.ram_data_o_7
rlabel metal1 7130 7888 7130 7888 0 manchester_baby_instance.ram_data_o_8
rlabel metal1 9108 5678 9108 5678 0 manchester_baby_instance.ram_data_o_9
rlabel metal2 1702 14076 1702 14076 0 net1
rlabel metal1 7360 14926 7360 14926 0 net10
rlabel metal1 20608 16082 20608 16082 0 net11
rlabel metal1 19826 13940 19826 13940 0 net12
rlabel metal1 14122 17646 14122 17646 0 net13
rlabel via1 18174 24106 18174 24106 0 net14
rlabel metal1 18492 25126 18492 25126 0 net15
rlabel metal1 14490 25874 14490 25874 0 net16
rlabel metal2 15594 25738 15594 25738 0 net17
rlabel via1 16969 25942 16969 25942 0 net18
rlabel metal1 14812 26282 14812 26282 0 net19
rlabel metal1 17572 24378 17572 24378 0 net2
rlabel metal2 19918 26690 19918 26690 0 net20
rlabel metal1 17894 25330 17894 25330 0 net21
rlabel metal1 14812 20910 14812 20910 0 net22
rlabel metal1 14352 20502 14352 20502 0 net23
rlabel metal1 18032 26894 18032 26894 0 net24
rlabel metal1 12420 14926 12420 14926 0 net25
rlabel metal1 6854 24072 6854 24072 0 net26
rlabel metal1 6808 19482 6808 19482 0 net27
rlabel metal1 10028 19482 10028 19482 0 net28
rlabel metal1 4370 18666 4370 18666 0 net29
rlabel metal1 13248 20026 13248 20026 0 net3
rlabel metal1 4646 20570 4646 20570 0 net30
rlabel metal1 13064 18394 13064 18394 0 net31
rlabel metal1 1702 19788 1702 19788 0 net4
rlabel metal1 1702 18836 1702 18836 0 net5
rlabel metal1 2231 19346 2231 19346 0 net6
rlabel metal1 4692 20298 4692 20298 0 net7
rlabel metal2 12650 17442 12650 17442 0 net8
rlabel metal1 15594 21046 15594 21046 0 net9
rlabel metal1 13156 29274 13156 29274 0 ram_addr_o[0]
rlabel metal3 820 19788 820 19788 0 ram_addr_o[1]
rlabel metal3 820 18428 820 18428 0 ram_addr_o[2]
rlabel metal3 1096 19108 1096 19108 0 ram_addr_o[3]
rlabel metal3 751 20468 751 20468 0 ram_addr_o[4]
rlabel metal2 12650 16898 12650 16898 0 ram_data_io[0]
rlabel metal2 12282 823 12282 823 0 ram_data_io[10]
rlabel metal2 18078 6562 18078 6562 0 ram_data_io[11]
rlabel metal2 18170 6256 18170 6256 0 ram_data_io[12]
rlabel metal1 18768 12206 18768 12206 0 ram_data_io[13]
rlabel metal1 17020 13838 17020 13838 0 ram_data_io[14]
rlabel metal1 15502 4114 15502 4114 0 ram_data_io[15]
rlabel metal1 20654 7820 20654 7820 0 ram_data_io[16]
rlabel metal2 21390 6783 21390 6783 0 ram_data_io[17]
rlabel metal2 22586 1761 22586 1761 0 ram_data_io[18]
rlabel metal3 30161 10948 30161 10948 0 ram_data_io[19]
rlabel metal1 9982 14892 9982 14892 0 ram_data_io[1]
rlabel metal1 21666 13294 21666 13294 0 ram_data_io[20]
rlabel metal2 21942 16286 21942 16286 0 ram_data_io[21]
rlabel metal1 23138 17034 23138 17034 0 ram_data_io[22]
rlabel metal1 29302 16558 29302 16558 0 ram_data_io[23]
rlabel metal1 27278 18292 27278 18292 0 ram_data_io[24]
rlabel metal1 28060 19890 28060 19890 0 ram_data_io[25]
rlabel metal3 30161 21148 30161 21148 0 ram_data_io[26]
rlabel metal1 25530 21386 25530 21386 0 ram_data_io[27]
rlabel metal1 23046 19822 23046 19822 0 ram_data_io[28]
rlabel metal1 20792 20434 20792 20434 0 ram_data_io[29]
rlabel metal1 7038 15572 7038 15572 0 ram_data_io[2]
rlabel metal1 19458 17714 19458 17714 0 ram_data_io[30]
rlabel metal1 15042 18734 15042 18734 0 ram_data_io[31]
rlabel metal2 4462 15810 4462 15810 0 ram_data_io[3]
rlabel metal1 4830 13804 4830 13804 0 ram_data_io[4]
rlabel metal1 5198 12308 5198 12308 0 ram_data_io[5]
rlabel metal1 5474 10676 5474 10676 0 ram_data_io[6]
rlabel metal1 7452 9622 7452 9622 0 ram_data_io[7]
rlabel metal1 5658 7956 5658 7956 0 ram_data_io[8]
rlabel metal1 9752 6290 9752 6290 0 ram_data_io[9]
rlabel metal3 820 21148 820 21148 0 ram_rw_en_o
rlabel metal3 820 14348 820 14348 0 reset_i
rlabel metal1 15594 29274 15594 29274 0 stop_lamp_o
<< properties >>
string FIXED_BBOX 0 0 32000 32000
<< end >>
