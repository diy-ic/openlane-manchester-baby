* NGSPICE file created from openlane_manchester_baby.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt openlane_manchester_baby VGND VPWR clock logisim_clock_tree_0_out ram_addr_o[0]
+ ram_addr_o[1] ram_addr_o[2] ram_addr_o[3] ram_addr_o[4] ram_data_io[0] ram_data_io[10]
+ ram_data_io[11] ram_data_io[12] ram_data_io[13] ram_data_io[14] ram_data_io[15]
+ ram_data_io[16] ram_data_io[17] ram_data_io[18] ram_data_io[19] ram_data_io[1] ram_data_io[20]
+ ram_data_io[21] ram_data_io[22] ram_data_io[23] ram_data_io[24] ram_data_io[25]
+ ram_data_io[26] ram_data_io[27] ram_data_io[28] ram_data_io[29] ram_data_io[2] ram_data_io[30]
+ ram_data_io[31] ram_data_io[3] ram_data_io[4] ram_data_io[5] ram_data_io[6] ram_data_io[7]
+ ram_data_io[8] ram_data_io[9] ram_rw_en_o reset_i stop_lamp_o
XFILLER_0_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_247 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ clknet_2_2__leaf_clock _0094_ _0043_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_12
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0985_ _0461_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_14_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ _0196_ _0253_ _0266_ _0271_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a31o_1
X_1253_ clknet_2_1__leaf_clock _0077_ _0026_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1184_ _0547_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0968_ manchester_baby_instance.ram_data_o_31 _0445_ _0446_ VGND VGND VPWR VPWR _0447_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0899_ _0379_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ _0311_ _0315_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0753_ _0158_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__xnor2_1
X_0684_ _0106_ _0180_ _0183_ _0193_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a32o_1
X_1305_ manchester_baby_instance.ram_data_o_28 _0584_ VGND VGND VPWR VPWR ram_data_io[28]
+ sky130_fd_sc_hd__ebufn_8
X_1236_ ram_data_io[17] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_17
+ sky130_fd_sc_hd__dlxtn_1
X_1167_ net1 VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__buf_4
X_1098_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1021_ _0173_ _0400_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0805_ _0239_ _0294_ _0300_ _0301_ _0229_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a32o_1
X_0736_ _0140_ _0155_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__nor2_1
X_0667_ _0107_ _0108_ _0176_ _0177_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a311o_1
X_0598_ _0109_ _0110_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__nor2_1
X_1219_ ram_data_io[0] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_0
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_15_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1004_ _0204_ _0470_ _0475_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0719_ _0163_ _0216_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput7 net7 VGND VGND VPWR VPWR ram_addr_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_41_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_37_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ manchester_baby_instance.ram_data_o_29 _0460_ _0446_ VGND VGND VPWR VPWR _0461_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1252_ clknet_2_3__leaf_clock _0000_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.Acc.tick
+ sky130_fd_sc_hd__dfxtp_1
X_1183_ _0547_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0967_ _0198_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ net28 manchester_baby_instance.ram_data_i_1 _0372_ VGND VGND VPWR VPWR _0379_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0102_ VGND VGND
+ VPWR VPWR _0315_ sky130_fd_sc_hd__and2b_1
X_0752_ _0140_ _0155_ _0153_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_24_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1166_ _0550_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
X_1304_ manchester_baby_instance.ram_data_o_27 _0583_ VGND VGND VPWR VPWR ram_data_io[27]
+ sky130_fd_sc_hd__ebufn_8
X_1235_ ram_data_io[16] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_16
+ sky130_fd_sc_hd__dlxtn_1
X_1097_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__nand4b_2
XTAP_TAPCELL_ROW_22_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ _0491_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_44_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0735_ manchester_baby_instance.ram_data_o_10 manchester_baby_instance.ram_data_i_10
+ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0804_ _0124_ _0128_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__xor2_1
X_0666_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__inv_2
X_0597_ manchester_baby_instance.ram_data_o_7 manchester_baby_instance.ram_data_i_7
+ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__and2b_1
X_1149_ net20 manchester_baby_instance.BASE_0.s_tickReg VGND VGND VPWR VPWR _0551_
+ sky130_fd_sc_hd__or2b_1
X_1218_ clknet_2_3__leaf_clock net18 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_tickReg
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0194_ _0467_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0718_ manchester_baby_instance.ram_data_i_13 _0187_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nand2_1
X_0649_ manchester_baby_instance.ram_data_i_14 manchester_baby_instance.ram_data_o_14
+ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_11_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput8 net13 VGND VGND VPWR VPWR ram_rw_en_o sky130_fd_sc_hd__buf_2
XFILLER_0_41_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ _0239_ _0442_ _0455_ _0459_ _0229_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1251_ clknet_2_3__leaf_clock net14 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfxtp_1
X_1182_ _0547_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ _0106_ _0435_ _0436_ _0196_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a32o_1
X_0897_ _0378_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0820_ _0312_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0751_ manchester_baby_instance.ram_data_i_9 _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__nand2_1
X_1303_ manchester_baby_instance.ram_data_o_26 _0582_ VGND VGND VPWR VPWR ram_data_io[26]
+ sky130_fd_sc_hd__ebufn_8
X_0682_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_4
X_1165_ _0550_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1096_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nand4b_2
X_1234_ ram_data_io[15] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_15
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_22_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ manchester_baby_instance.ram_data_o_29 manchester_baby_instance.ram_data_i_29
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_30_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0734_ manchester_baby_instance.ram_data_i_11 _0232_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__nand2_1
X_0665_ manchester_baby_instance.ram_data_o_18 manchester_baby_instance.ram_data_i_18
+ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0803_ _0118_ _0293_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
X_0596_ manchester_baby_instance.ram_data_i_7 manchester_baby_instance.ram_data_o_7
+ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1217_ clknet_2_3__leaf_clock _0076_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1079_ _0331_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__buf_4
X_1148_ _0550_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold10 _0072_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ manchester_baby_instance.ram_data_i_26 _0440_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0648_ manchester_baby_instance.ram_data_o_15 manchester_baby_instance.ram_data_i_15
+ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and2b_1
X_0717_ _0225_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR stop_lamp_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0982_ _0457_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_14_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1250_ ram_data_io[31] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_31
+ sky130_fd_sc_hd__dlxtn_1
X_1181_ _0547_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0896_ net27 _0118_ _0372_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux2_1
X_0965_ manchester_baby_instance.ram_data_i_31 _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ manchester_baby_instance.ram_data_i_8 _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0681_ _0104_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0103_ _0101_ VGND VGND
+ VPWR VPWR _0194_ sky130_fd_sc_hd__and4bb_2
X_1302_ manchester_baby_instance.ram_data_o_25 _0581_ VGND VGND VPWR VPWR ram_data_io[25]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1233_ ram_data_io[14] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_14
+ sky130_fd_sc_hd__dlxtn_1
X_1164_ _0550_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
X_1095_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__nand4b_2
X_0948_ manchester_baby_instance.ram_data_i_29 manchester_baby_instance.ram_data_o_29
+ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0879_ _0332_ _0321_ _0368_ _0343_ manchester_baby_instance.ram_data_i_0 VGND VGND
+ VPWR VPWR _0369_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_30_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0802_ _0299_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_0664_ manchester_baby_instance.ram_data_o_17 manchester_baby_instance.ram_data_i_17
+ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__and2b_1
X_0733_ _0195_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1216_ clknet_2_3__leaf_clock _0075_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_0595_ manchester_baby_instance.ram_data_i_16 manchester_baby_instance.ram_data_o_16
+ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1078_ _0101_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__buf_4
X_1147_ net1 VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 manchester_baby_instance.BASE_0.s_tickReg VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ _0469_ _0412_ _0418_ _0421_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0647_ _0152_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0716_ manchester_baby_instance.ram_data_o_14 _0224_ _0199_ VGND VGND VPWR VPWR _0225_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ _0456_ _0382_ _0426_ _0427_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clock clock VGND VGND VPWR VPWR clknet_0_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0547_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0964_ manchester_baby_instance.ram_data_i_30 _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or2_1
X_0895_ _0377_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0680_ manchester_baby_instance.ram_data_i_18 _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__xor2_1
X_1232_ ram_data_io[13] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_13
+ sky130_fd_sc_hd__dlxtn_1
X_1301_ manchester_baby_instance.ram_data_o_24 _0580_ VGND VGND VPWR VPWR ram_data_io[24]
+ sky130_fd_sc_hd__ebufn_8
X_1163_ _0550_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1094_ _0526_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__buf_4
X_0947_ _0420_ _0423_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_30_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0878_ _0337_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ manchester_baby_instance.ram_data_o_3 _0298_ _0251_ VGND VGND VPWR VPWR _0299_
+ sky130_fd_sc_hd__mux2_1
X_0594_ manchester_baby_instance.ram_data_i_17 manchester_baby_instance.ram_data_o_17
+ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__or2b_1
X_0732_ _0238_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_0663_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1215_ clknet_2_1__leaf_clock _0074_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ _0549_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1077_ _0104_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold12 manchester_baby_instance.ram_data_o_0 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ _0474_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0715_ _0196_ _0211_ _0222_ _0223_ _0204_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a32o_1
X_0646_ _0155_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1129_ _0548_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ manchester_baby_instance.ram_data_o_14 manchester_baby_instance.ram_data_i_14
+ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0382_ _0426_ _0427_ _0456_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0963_ manchester_baby_instance.ram_data_i_28 manchester_baby_instance.ram_data_i_29
+ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or3_1
X_0894_ net29 manchester_baby_instance.ram_data_i_3 _0372_ VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1162_ _0550_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
X_1231_ ram_data_io[12] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_12
+ sky130_fd_sc_hd__dlxtn_1
X_1300_ manchester_baby_instance.ram_data_o_23 _0579_ VGND VGND VPWR VPWR ram_data_io[23]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_47_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ _0331_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0877_ manchester_baby_instance.ram_data_o_31 _0334_ _0337_ VGND VGND VPWR VPWR _0367_
+ sky130_fd_sc_hd__and3b_1
X_0946_ _0382_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0731_ manchester_baby_instance.ram_data_o_12 _0237_ _0199_ VGND VGND VPWR VPWR _0238_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ _0239_ _0184_ _0295_ _0297_ _0229_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a32o_1
X_0662_ _0173_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__and2b_1
X_0593_ _0105_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ clknet_2_3__leaf_clock _0073_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_counterValue
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1145_ _0549_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0929_ _0407_ _0395_ _0392_ _0394_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_45_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold13 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] VGND VGND VPWR VPWR
+ net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0645_ _0156_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__nand2_1
X_0714_ _0142_ _0217_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__xnor2_1
X_1059_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1128_ _0548_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ manchester_baby_instance.ram_data_o_15 manchester_baby_instance.ram_data_i_15
+ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0962_ manchester_baby_instance.ram_data_i_26 manchester_baby_instance.ram_data_i_27
+ _0440_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or3_1
X_0893_ _0376_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1161_ _0554_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ _0101_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__buf_4
X_1230_ ram_data_io[11] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_11
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_47_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0876_ _0337_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__inv_2
X_0945_ manchester_baby_instance.ram_data_o_28 manchester_baby_instance.ram_data_i_28
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0730_ _0196_ _0187_ _0234_ _0236_ _0229_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a32o_1
X_0661_ manchester_baby_instance.ram_data_o_16 manchester_baby_instance.ram_data_i_16
+ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ clknet_2_3__leaf_clock net15 VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0592_ _0101_ _0103_ _0104_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1144_ _0549_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
X_1075_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0859_ _0317_ _0339_ _0341_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or3_1
X_0928_ _0387_ _0401_ _0406_ _0386_ _0391_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__a311o_1
Xhold14 manchester_baby_instance.CIRCUIT_0.IR.q\[2\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0644_ manchester_baby_instance.ram_data_o_9 manchester_baby_instance.ram_data_i_9
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2b_1
X_0713_ manchester_baby_instance.ram_data_i_14 _0188_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__nand2_1
X_1058_ _0524_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
X_1127_ _0548_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0627_ _0113_ _0116_ _0133_ _0139_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0961_ manchester_baby_instance.ram_data_i_23 manchester_baby_instance.ram_data_i_24
+ manchester_baby_instance.ram_data_i_25 _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or4_1
X_0892_ net30 manchester_baby_instance.ram_data_i_4 _0372_ VGND VGND VPWR VPWR _0376_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1160_ net17 _0539_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2_1
X_1091_ _0104_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_2
X_0944_ _0419_ _0421_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0319_ _0317_ _0365_ _0316_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1289_ manchester_baby_instance.ram_data_o_12 _0568_ VGND VGND VPWR VPWR ram_data_io[12]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_21_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0660_ _0140_ _0149_ _0160_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__o31a_2
X_0591_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1212_ clknet_2_3__leaf_clock net23 _0025_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ _0549_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ _0405_ _0389_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__nand2_1
X_0858_ _0335_ _0340_ _0344_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0789_ _0132_ _0282_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
Xhold15 manchester_baby_instance.CIRCUIT_0.IR.q\[1\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0643_ manchester_baby_instance.ram_data_i_9 manchester_baby_instance.ram_data_o_9
+ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0712_ _0221_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ _0548_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_2
X_1057_ manchester_baby_instance.ram_data_o_19 _0523_ _0198_ VGND VGND VPWR VPWR _0524_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0626_ _0113_ _0135_ _0138_ _0109_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0540_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0609_ _0118_ manchester_baby_instance.ram_data_o_2 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0960_ manchester_baby_instance.ram_data_i_20 manchester_baby_instance.ram_data_i_21
+ manchester_baby_instance.ram_data_i_22 _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0891_ _0375_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nand4b_2
X_0943_ _0414_ _0416_ _0413_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o21ba_1
X_0874_ manchester_baby_instance.ram_data_i_1 _0343_ _0361_ _0334_ _0364_ VGND VGND
+ VPWR VPWR _0365_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1288_ manchester_baby_instance.ram_data_o_11 _0567_ VGND VGND VPWR VPWR ram_data_io[11]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_21_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0590_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0102_ VGND VGND
+ VPWR VPWR _0103_ sky130_fd_sc_hd__and2_2
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1211_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
+ _0024_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_1142_ _0549_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1073_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__nand4b_2
X_0857_ manchester_baby_instance.ram_data_i_3 _0343_ _0349_ _0332_ VGND VGND VPWR
+ VPWR _0350_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ manchester_baby_instance.ram_data_o_19 _0402_ _0182_ _0399_ _0404_ VGND VGND
+ VPWR VPWR _0405_ sky130_fd_sc_hd__a221o_1
Xhold16 manchester_baby_instance.CIRCUIT_0.IR.q\[3\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
X_0788_ _0287_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_2__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0711_ manchester_baby_instance.ram_data_o_15 _0220_ _0199_ VGND VGND VPWR VPWR _0221_
+ sky130_fd_sc_hd__mux2_1
X_0642_ _0153_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1125_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_49_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1056_ _0195_ _0438_ _0520_ _0522_ _0106_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a32o_1
XFILLER_0_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0909_ _0386_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0625_ _0137_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1108_ _0102_ _0525_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1039_ manchester_baby_instance.ram_data_o_22 _0508_ _0446_ VGND VGND VPWR VPWR _0509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0608_ _0117_ _0118_ _0119_ _0120_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__o31a_1
XFILLER_0_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0890_ _0331_ manchester_baby_instance.ram_data_i_13 _0372_ VGND VGND VPWR VPWR _0375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ _0383_ _0411_ _0410_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__a21o_1
X_0873_ _0332_ _0322_ _0362_ _0363_ _0315_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ manchester_baby_instance.ram_data_o_10 _0566_ VGND VGND VPWR VPWR ram_data_io[10]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_21_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
+ _0023_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1141_ _0549_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1072_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nand4b_2
XPHY_EDGE_ROW_23_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0856_ _0325_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0925_ manchester_baby_instance.ram_data_o_19 _0402_ _0403_ VGND VGND VPWR VPWR _0404_
+ sky130_fd_sc_hd__o21a_1
X_0787_ manchester_baby_instance.ram_data_o_5 _0286_ _0251_ VGND VGND VPWR VPWR _0287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 manchester_baby_instance.CIRCUIT_0.IR.q\[4\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0641_ manchester_baby_instance.ram_data_o_8 manchester_baby_instance.ram_data_i_8
+ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0710_ _0196_ _0190_ _0212_ _0219_ _0204_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1055_ _0398_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1124_ net1 VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__buf_4
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0839_ _0329_ _0330_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__o21a_1
X_0908_ manchester_baby_instance.ram_data_i_21 manchester_baby_instance.ram_data_o_21
+ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0624_ _0110_ _0136_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__or2_1
X_1107_ net17 _0539_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_tickNext
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ _0204_ _0495_ _0503_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0607_ manchester_baby_instance.ram_data_i_3 manchester_baby_instance.ram_data_o_3
+ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0941_ _0385_ _0409_ _0412_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or4_1
X_0872_ _0319_ _0337_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_38_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ manchester_baby_instance.ram_data_o_9 _0565_ VGND VGND VPWR VPWR ram_data_io[9]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ _0549_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ manchester_baby_instance.ram_data_i_18 manchester_baby_instance.ram_data_o_18
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__and2b_1
X_0855_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__xnor2_1
X_0786_ _0239_ _0276_ _0281_ _0285_ _0229_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold18 manchester_baby_instance.CIRCUIT_0.IR.q\[0\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
X_1269_ clknet_2_2__leaf_clock _0093_ _0042_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_11
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_40_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0640_ manchester_baby_instance.ram_data_i_8 manchester_baby_instance.ram_data_o_8
+ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1123_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0545_ _0546_ manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__a22o_1
X_1054_ _0403_ _0180_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0907_ manchester_baby_instance.ram_data_o_21 manchester_baby_instance.ram_data_i_21
+ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0838_ _0331_ _0311_ _0312_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and3_1
X_0769_ _0261_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0623_ manchester_baby_instance.ram_data_i_6 manchester_baby_instance.ram_data_o_6
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__or2b_1
X_1106_ net16 net19 VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ _0194_ _0439_ _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0606_ manchester_baby_instance.ram_data_o_3 manchester_baby_instance.ram_data_i_3
+ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout10 net13 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0940_ _0415_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0871_ _0320_ _0321_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nand2_1
X_1285_ manchester_baby_instance.ram_data_o_8 _0564_ VGND VGND VPWR VPWR ram_data_io[8]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_38_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__nand4b_2
X_0854_ net26 _0317_ _0347_ _0316_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0923_ manchester_baby_instance.ram_data_i_19 VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0785_ _0116_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__xor2_1
X_1268_ clknet_2_0__leaf_clock _0092_ _0041_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_10
+ sky130_fd_sc_hd__dfrtp_1
X_1199_ clknet_2_3__leaf_clock _0062_ _0013_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_31
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1122_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0545_ _0546_ manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__a22o_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1053_ manchester_baby_instance.ram_data_i_17 manchester_baby_instance.ram_data_i_18
+ _0191_ manchester_baby_instance.ram_data_i_19 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ _0383_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0837_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0699_ manchester_baby_instance.ram_data_o_16 _0209_ _0199_ VGND VGND VPWR VPWR _0210_
+ sky130_fd_sc_hd__mux2_1
X_0768_ _0111_ _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0622_ _0115_ _0134_ _0114_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__a21oi_1
X_1105_ _0104_ _0101_ _0331_ _0526_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__nand4b_2
X_1036_ manchester_baby_instance.ram_data_i_22 _0505_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ manchester_baby_instance.ram_data_i_2 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__buf_2
X_1019_ manchester_baby_instance.ram_data_o_24 _0490_ _0446_ VGND VGND VPWR VPWR _0491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout11 net12 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_0_36_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ _0338_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1284_ manchester_baby_instance.ram_data_o_7 _0563_ VGND VGND VPWR VPWR ram_data_io[7]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_46_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0999_ manchester_baby_instance.ram_data_o_27 _0473_ _0446_ VGND VGND VPWR VPWR _0474_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0853_ _0333_ _0342_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or3b_1
X_0922_ manchester_baby_instance.ram_data_i_20 manchester_baby_instance.ram_data_o_20
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or2b_1
X_0784_ _0134_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nand2_1
X_1267_ clknet_2_0__leaf_clock _0091_ _0040_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_9
+ sky130_fd_sc_hd__dfrtp_1
Xinput1 reset_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
X_1198_ clknet_2_3__leaf_clock _0061_ _0012_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_30
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_27_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0545_ _0546_ manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__a22o_1
X_1052_ _0519_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0836_ manchester_baby_instance.ram_data_i_4 _0328_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0767_ _0267_ _0268_ _0136_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o21ai_1
X_0905_ manchester_baby_instance.ram_data_o_24 manchester_baby_instance.ram_data_i_24
+ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0698_ _0196_ _0191_ _0207_ _0208_ _0204_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0621_ manchester_baby_instance.ram_data_i_4 manchester_baby_instance.ram_data_o_4
+ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1035_ manchester_baby_instance.ram_data_i_21 _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__or2_1
X_1104_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__nand4b_2
XTAP_TAPCELL_ROW_16_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0819_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0604_ manchester_baby_instance.ram_data_o_2 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ _0204_ _0469_ _0487_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_14_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout12 net13 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_0_19_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1283_ manchester_baby_instance.ram_data_o_6 _0562_ VGND VGND VPWR VPWR ram_data_io[6]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_46_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ _0195_ _0441_ _0468_ _0472_ _0106_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0181_ _0174_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nand3_1
X_0852_ manchester_baby_instance.ram_data_i_4 _0343_ _0345_ VGND VGND VPWR VPWR _0346_
+ sky130_fd_sc_hd__a21oi_1
X_0783_ _0132_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1197_ clknet_2_3__leaf_clock _0060_ _0011_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_29
+ sky130_fd_sc_hd__dfrtp_1
X_1266_ clknet_2_0__leaf_clock _0090_ _0039_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_8
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1120_ _0319_ _0545_ _0546_ manchester_baby_instance.CIRCUIT_0.IR.q\[1\] VGND VGND
+ VPWR VPWR net4 sky130_fd_sc_hd__a22o_1
X_1051_ manchester_baby_instance.ram_data_o_20 _0518_ _0198_ VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0904_ manchester_baby_instance.ram_data_i_24 manchester_baby_instance.ram_data_o_24
+ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or2b_1
X_0835_ manchester_baby_instance.ram_data_i_4 _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0697_ _0174_ _0173_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__xnor2_1
X_0766_ _0116_ _0133_ _0135_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1249_ ram_data_io[30] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_30
+ sky130_fd_sc_hd__dlxtn_1
XPHY_EDGE_ROW_44_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0620_ _0121_ _0131_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1103_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nand4b_2
X_1034_ manchester_baby_instance.ram_data_i_20 _0438_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0818_ _0104_ _0101_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__nor2_1
X_0749_ manchester_baby_instance.ram_data_i_7 _0185_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0603_ _0114_ _0115_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ _0194_ _0481_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 net8 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ manchester_baby_instance.ram_data_o_5 _0561_ VGND VGND VPWR VPWR ram_data_io[5]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_46_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0997_ _0415_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0178_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and2_1
X_0851_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ _0340_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__and4b_1
X_0782_ _0121_ _0131_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__nand2_1
X_1265_ clknet_2_0__leaf_clock _0089_ _0038_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_7
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1196_ clknet_2_3__leaf_clock _0059_ _0010_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_28
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1050_ _0204_ _0494_ _0515_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0834_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0327_ VGND VGND VPWR
+ VPWR _0328_ sky130_fd_sc_hd__xnor2_1
X_0903_ manchester_baby_instance.ram_data_i_28 manchester_baby_instance.ram_data_o_28
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0696_ manchester_baby_instance.ram_data_i_16 _0190_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nand2_1
X_0765_ _0112_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__inv_2
X_1248_ ram_data_io[29] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_29
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1179_ _0547_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_17_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1033_ _0502_ _0393_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or2b_1
X_0817_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0311_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_16_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0748_ _0252_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_0679_ manchester_baby_instance.ram_data_i_17 _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0602_ manchester_baby_instance.ram_data_i_5 manchester_baby_instance.ram_data_o_5
+ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1016_ manchester_baby_instance.ram_data_i_24 _0480_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1281_ manchester_baby_instance.ram_data_o_4 _0560_ VGND VGND VPWR VPWR ram_data_io[4]
+ sky130_fd_sc_hd__ebufn_8
XTAP_TAPCELL_ROW_46_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ _0416_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_107 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ manchester_baby_instance.ram_data_o_31 _0334_ _0315_ VGND VGND VPWR VPWR _0344_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0781_ manchester_baby_instance.ram_data_i_5 _0275_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__nand2_1
X_1264_ clknet_2_0__leaf_clock _0088_ _0037_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_6
+ sky130_fd_sc_hd__dfrtp_2
X_1195_ clknet_2_3__leaf_clock _0058_ _0009_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_27
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0979_ manchester_baby_instance.ram_data_o_29 manchester_baby_instance.ram_data_i_29
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_40_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21o_1
X_0902_ manchester_baby_instance.ram_data_i_30 manchester_baby_instance.ram_data_o_30
+ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and2b_1
X_0695_ _0206_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0764_ manchester_baby_instance.ram_data_i_7 _0185_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1247_ ram_data_io[28] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_28
+ sky130_fd_sc_hd__dlxtn_1
X_1178_ _0547_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ _0387_ _0401_ _0494_ _0386_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_33_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0747_ manchester_baby_instance.ram_data_o_10 _0250_ _0251_ VGND VGND VPWR VPWR _0252_
+ sky130_fd_sc_hd__mux2_1
X_0816_ manchester_baby_instance.ram_data_i_0 _0199_ _0309_ _0310_ net25 VGND VGND
+ VPWR VPWR _0082_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0678_ manchester_baby_instance.ram_data_i_16 _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0601_ manchester_baby_instance.ram_data_o_5 manchester_baby_instance.ram_data_i_5
+ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0385_ _0409_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1280_ manchester_baby_instance.ram_data_o_3 _0559_ VGND VGND VPWR VPWR ram_data_io[3]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0995_ _0383_ _0469_ _0411_ _0418_ _0410_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a311o_1
XFILLER_0_18_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ _0280_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1194_ clknet_2_3__leaf_clock _0057_ _0008_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_26
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1263_ clknet_2_0__leaf_clock _0087_ _0036_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_5
+ sky130_fd_sc_hd__dfrtp_1
X_0978_ manchester_baby_instance.ram_data_i_29 _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0832_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o21a_1
X_0901_ _0380_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_0763_ _0265_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0694_ manchester_baby_instance.ram_data_o_17 _0205_ _0199_ VGND VGND VPWR VPWR _0206_
+ sky130_fd_sc_hd__mux2_1
X_1246_ ram_data_io[27] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_27
+ sky130_fd_sc_hd__dlxtn_1
X_1177_ _0555_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1100_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1031_ _0501_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0746_ _0198_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__buf_4
X_0815_ manchester_baby_instance.ram_data_i_0 _0261_ _0199_ VGND VGND VPWR VPWR _0310_
+ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_48_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0677_ _0188_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__or2_1
X_1229_ ram_data_io[10] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_10
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0600_ _0111_ _0112_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_242 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0486_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0729_ _0144_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0994_ _0385_ _0409_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1193_ clknet_2_3__leaf_clock _0056_ _0007_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_25
+ sky130_fd_sc_hd__dfrtp_1
X_1262_ clknet_2_0__leaf_clock _0086_ _0035_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_4
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ manchester_baby_instance.ram_data_i_28 _0441_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ net31 manchester_baby_instance.ram_data_i_0 _0372_ VGND VGND VPWR VPWR _0380_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0831_ _0318_ _0323_ _0324_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__o21ai_1
X_0762_ manchester_baby_instance.ram_data_o_8 _0264_ _0251_ VGND VGND VPWR VPWR _0265_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0693_ _0196_ _0192_ _0201_ _0203_ _0204_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ ram_data_io[26] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_26
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1176_ _0555_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ manchester_baby_instance.ram_data_o_23 _0500_ _0446_ VGND VGND VPWR VPWR _0501_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0814_ _0196_ manchester_baby_instance.ram_data_o_0 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0745_ _0239_ _0232_ _0248_ _0249_ _0229_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__a32o_1
X_0676_ manchester_baby_instance.ram_data_i_15 manchester_baby_instance.ram_data_i_14
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1228_ ram_data_io[9] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_9
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ _0539_ _0553_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ manchester_baby_instance.ram_data_o_25 _0485_ _0446_ VGND VGND VPWR VPWR _0486_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0728_ _0169_ _0214_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__nor2_1
X_0659_ _0161_ _0162_ _0164_ _0170_ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ manchester_baby_instance.ram_data_i_27 _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1261_ clknet_2_0__leaf_clock _0085_ _0034_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_3
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1192_ clknet_2_3__leaf_clock _0055_ _0006_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_24
+ sky130_fd_sc_hd__dfrtp_1
X_0976_ _0453_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0830_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0118_ VGND VGND VPWR
+ VPWR _0324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0761_ _0239_ _0254_ _0260_ _0262_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0692_ _0106_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_4
X_1244_ ram_data_io[25] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_25
+ sky130_fd_sc_hd__dlxtn_1
X_1175_ _0555_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
X_0959_ manchester_baby_instance.ram_data_i_13 _0187_ _0189_ _0437_ VGND VGND VPWR
+ VPWR _0438_ sky130_fd_sc_hd__or4_2
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ _0308_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_0744_ _0151_ _0243_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__xnor2_1
X_0675_ manchester_baby_instance.ram_data_i_13 _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__or2_1
X_1158_ net16 net19 VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
X_1227_ ram_data_io[8] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_8
+ sky130_fd_sc_hd__dlxtn_1
X_1089_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__nand4b_2
XTAP_TAPCELL_ROW_7_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1012_ _0195_ _0440_ _0482_ _0484_ _0106_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ manchester_baby_instance.ram_data_i_12 _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__nand2_1
X_0589_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ manchester_baby_instance.ram_data_i_15 manchester_baby_instance.ram_data_o_15
+ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ manchester_baby_instance.ram_data_i_26 _0440_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__or2_1
Xclkbuf_2_1__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_1__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1191_ clknet_2_2__leaf_clock _0054_ _0005_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_23
+ sky130_fd_sc_hd__dfrtp_1
X_1260_ clknet_2_1__leaf_clock _0084_ _0033_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ manchester_baby_instance.ram_data_o_30 _0452_ _0446_ VGND VGND VPWR VPWR _0453_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0760_ _0140_ _0155_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nand2_1
X_0691_ _0181_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ ram_data_io[24] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_24
+ sky130_fd_sc_hd__dlxtn_1
X_1174_ _0555_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0958_ manchester_baby_instance.ram_data_i_16 manchester_baby_instance.ram_data_i_17
+ manchester_baby_instance.ram_data_i_18 manchester_baby_instance.ram_data_i_19 VGND
+ VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
X_0889_ _0374_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_25 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ manchester_baby_instance.ram_data_i_10 _0186_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0812_ manchester_baby_instance.ram_data_o_1 _0307_ _0251_ VGND VGND VPWR VPWR _0308_
+ sky130_fd_sc_hd__mux2_1
X_0674_ manchester_baby_instance.ram_data_i_10 manchester_baby_instance.ram_data_i_11
+ manchester_baby_instance.ram_data_i_12 _0186_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__or4_2
X_1157_ net16 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
X_1226_ ram_data_io[7] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_7
+ sky130_fd_sc_hd__dlxtn_1
X_1088_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ _0412_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0726_ manchester_baby_instance.ram_data_i_11 _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0657_ _0149_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or2b_1
X_0588_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_4
X_1209_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
+ _0022_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0141_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_23_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0991_ _0466_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ clknet_2_2__leaf_clock _0053_ _0004_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_22
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ _0239_ _0443_ _0448_ _0449_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0690_ _0108_ _0176_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0555_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
X_1242_ ram_data_io[23] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_23
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ _0381_ _0432_ _0433_ _0434_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0888_ _0101_ manchester_baby_instance.ram_data_i_14 _0372_ VGND VGND VPWR VPWR _0374_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0742_ _0247_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ manchester_baby_instance.ram_data_i_7 manchester_baby_instance.ram_data_i_8
+ manchester_baby_instance.ram_data_i_9 _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0811_ _0239_ _0293_ _0304_ _0306_ _0229_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1156_ _0552_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_1087_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__nand4b_2
X_1225_ ram_data_io[6] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_6
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_15_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _0383_ _0469_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0656_ manchester_baby_instance.ram_data_o_11 _0165_ _0152_ _0166_ _0168_ VGND VGND
+ VPWR VPWR _0169_ sky130_fd_sc_hd__a221o_1
X_0725_ manchester_baby_instance.ram_data_i_10 _0186_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__or2_1
X_1208_ clknet_2_3__leaf_clock _0071_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_derivedClock
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1139_ _0549_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 manchester_baby_instance.BASE_1.s_bufferRegs\[0\] VGND VGND VPWR VPWR net14
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_49_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_13_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0708_ _0213_ _0217_ _0162_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0990_ manchester_baby_instance.ram_data_o_28 _0465_ _0446_ VGND VGND VPWR VPWR _0466_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0431_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1241_ ram_data_io[22] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_22
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0555_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
X_0956_ _0381_ _0432_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or4_1
XFILLER_0_42_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ _0373_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0810_ _0305_ _0126_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0741_ manchester_baby_instance.ram_data_o_11 _0246_ _0199_ VGND VGND VPWR VPWR _0247_
+ sky130_fd_sc_hd__mux2_1
X_0672_ manchester_baby_instance.ram_data_i_4 manchester_baby_instance.ram_data_i_5
+ manchester_baby_instance.ram_data_i_6 _0184_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__or4_1
X_1224_ ram_data_io[5] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_5
+ sky130_fd_sc_hd__dlxtn_1
X_1155_ net24 net20 VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__and2b_1
X_1086_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__nand4b_2
X_0939_ _0416_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0655_ manchester_baby_instance.ram_data_o_11 _0165_ _0167_ VGND VGND VPWR VPWR _0168_
+ sky130_fd_sc_hd__o21a_1
X_0724_ _0231_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1207_ clknet_2_2__leaf_clock _0070_ _0021_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1069_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nand4b_2
X_1138_ _0549_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 manchester_baby_instance.BASE_1.s_derivedClock VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ _0163_ _0147_ _0216_ _0146_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a31o_1
X_0638_ manchester_baby_instance.ram_data_o_10 manchester_baby_instance.ram_data_i_10
+ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ _0382_ _0426_ _0427_ _0428_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1171_ _0555_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
X_1240_ ram_data_io[21] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_21
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ manchester_baby_instance.ram_data_o_31 manchester_baby_instance.ram_data_i_31
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ _0104_ manchester_baby_instance.ram_data_i_15 _0372_ VGND VGND VPWR VPWR _0373_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ _0239_ _0233_ _0240_ _0245_ _0229_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0671_ manchester_baby_instance.ram_data_i_3 manchester_baby_instance.ram_data_i_2
+ manchester_baby_instance.ram_data_i_1 manchester_baby_instance.ram_data_i_0 VGND
+ VGND VPWR VPWR _0184_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1154_ _0550_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
X_1223_ ram_data_io[4] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_4
+ sky130_fd_sc_hd__dlxtn_2
X_1085_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__nand4b_2
X_0938_ manchester_baby_instance.ram_data_o_26 manchester_baby_instance.ram_data_i_26
+ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or2b_1
X_0869_ _0337_ manchester_baby_instance.ram_data_o_31 _0319_ VGND VGND VPWR VPWR _0360_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ manchester_baby_instance.ram_data_o_13 _0230_ _0199_ VGND VGND VPWR VPWR _0231_
+ sky130_fd_sc_hd__mux2_1
X_0654_ manchester_baby_instance.ram_data_i_10 manchester_baby_instance.ram_data_o_10
+ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1137_ _0549_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1206_ clknet_2_2__leaf_clock _0069_ _0020_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1068_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 manchester_baby_instance.BASE_0.s_countReg\[0\] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0706_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__inv_2
X_0637_ manchester_baby_instance.ram_data_o_11 manchester_baby_instance.ram_data_i_11
+ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_159 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0971_ _0261_ _0432_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0555_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__buf_2
X_0954_ manchester_baby_instance.ram_data_o_31 manchester_baby_instance.ram_data_i_31
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1299_ manchester_baby_instance.ram_data_o_22 _0578_ VGND VGND VPWR VPWR ram_data_io[22]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ _0181_ _0175_ _0178_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a211o_1
X_1153_ _0550_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
X_1084_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__nand4b_2
X_1222_ ram_data_io[3] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_3
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0868_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0317_ _0359_ _0316_
+ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a22o_1
X_0937_ manchester_baby_instance.ram_data_i_26 manchester_baby_instance.ram_data_o_26
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0799_ _0296_ _0130_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0653_ _0153_ _0156_ _0157_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0722_ _0196_ _0188_ _0226_ _0228_ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1067_ _0527_ _0528_ _0529_ _0530_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nand4b_2
X_1205_ clknet_2_2__leaf_clock _0068_ _0019_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1136_ net1 VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 manchester_baby_instance.BASE_0.s_countReg\[2\] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0705_ _0169_ _0214_ _0144_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o21a_1
X_0636_ _0143_ _0145_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ _0337_ _0545_ _0546_ manchester_baby_instance.CIRCUIT_0.IR.q\[0\] VGND VGND
+ VPWR VPWR net3 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ manchester_baby_instance.ram_data_o_4 manchester_baby_instance.ram_data_i_4
+ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0970_ manchester_baby_instance.ram_data_i_30 _0442_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.Acc.tick manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
+ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__and4b_1
X_0953_ _0382_ _0426_ _0427_ _0428_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1298_ manchester_baby_instance.ram_data_o_21 _0577_ VGND VGND VPWR VPWR ram_data_io[21]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_18_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ ram_data_io[2] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_2
+ sky130_fd_sc_hd__dlxtn_1
X_1152_ _0550_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
X_1083_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0936_ _0413_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0867_ _0118_ _0343_ _0353_ _0341_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ _0124_ _0128_ _0122_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0652_ manchester_baby_instance.ram_data_i_11 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0721_ _0106_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_4
X_1204_ clknet_2_1__leaf_clock _0067_ _0018_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1135_ _0548_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
X_1066_ _0526_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0919_ manchester_baby_instance.ram_data_o_19 manchester_baby_instance.ram_data_i_19
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 manchester_baby_instance.BASE_0.s_tickNext VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0704_ _0140_ _0160_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__nor2_1
X_0635_ _0146_ _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1118_ _0103_ _0312_ _0314_ _0526_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a22o_1
X_1049_ _0194_ _0504_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0618_ _0124_ _0128_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_34_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0883_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR
+ VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1297_ manchester_baby_instance.ram_data_o_20 _0576_ VGND VGND VPWR VPWR ram_data_io[20]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_18_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1151_ _0550_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
X_1220_ ram_data_io[1] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_1
+ sky130_fd_sc_hd__dlxtn_2
X_1082_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nand4b_2
X_0935_ manchester_baby_instance.ram_data_o_27 manchester_baby_instance.ram_data_i_27
+ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__and2b_1
X_0866_ _0332_ _0356_ _0357_ _0339_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0797_ manchester_baby_instance.ram_data_i_3 _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ _0148_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__xnor2_1
X_0651_ _0163_ _0147_ _0146_ _0143_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1134_ _0548_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1203_ clknet_2_1__leaf_clock _0066_ _0017_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0331_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__buf_4
X_0849_ _0331_ _0311_ _0312_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__and3b_1
X_0918_ _0390_ _0393_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 manchester_baby_instance.BASE_0.s_countReg\[1\] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0703_ manchester_baby_instance.ram_data_o_14 manchester_baby_instance.ram_data_i_14
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__and2b_1
X_0634_ manchester_baby_instance.ram_data_i_13 manchester_baby_instance.ram_data_o_13
+ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_48_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0545_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ manchester_baby_instance.ram_data_i_20 _0438_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0617_ _0120_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0882_ manchester_baby_instance.CIRCUIT_0.Acc.tick _0331_ _0103_ _0313_ net22 VGND
+ VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a41o_1
X_0951_ _0381_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1296_ manchester_baby_instance.ram_data_o_19 _0575_ VGND VGND VPWR VPWR ram_data_io[19]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1150_ net15 net21 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__xnor2_1
X_1081_ _0531_ _0532_ _0533_ _0534_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_23_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0934_ manchester_baby_instance.ram_data_i_27 manchester_baby_instance.ram_data_o_27
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and2b_1
X_0865_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0338_ VGND VGND VPWR
+ VPWR _0357_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ _0118_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__or2_1
X_1279_ manchester_baby_instance.ram_data_o_2 _0558_ VGND VGND VPWR VPWR ram_data_io[2]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_271 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0650_ manchester_baby_instance.ram_data_i_12 manchester_baby_instance.ram_data_o_12
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or2b_1
X_1133_ _0548_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
X_1202_ clknet_2_1__leaf_clock _0065_ _0016_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1064_ _0101_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0848_ _0336_ _0339_ _0341_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o31a_1
X_0779_ manchester_baby_instance.ram_data_o_6 _0279_ _0251_ VGND VGND VPWR VPWR _0280_
+ sky130_fd_sc_hd__mux2_1
X_0917_ _0394_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_3_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold7 manchester_baby_instance.BASE_1.s_counterValue VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0633_ manchester_baby_instance.ram_data_o_13 manchester_baby_instance.ram_data_i_13
+ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2b_1
X_0702_ manchester_baby_instance.ram_data_i_15 _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1116_ _0544_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.GATES_13.result
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ _0405_ _0389_ _0492_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0616_ manchester_baby_instance.ram_data_o_3 manchester_baby_instance.ram_data_i_3
+ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ _0337_ _0317_ _0370_ _0316_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ manchester_baby_instance.ram_data_o_30 manchester_baby_instance.ram_data_i_30
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and2b_1
XFILLER_0_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1295_ manchester_baby_instance.ram_data_o_18 _0574_ VGND VGND VPWR VPWR ram_data_io[18]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_41_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1080_ _0526_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0933_ _0410_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or2b_1
X_0864_ _0323_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ manchester_baby_instance.ram_data_i_1 manchester_baby_instance.ram_data_i_0
+ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1278_ manchester_baby_instance.ram_data_o_1 _0557_ VGND VGND VPWR VPWR ram_data_io[1]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_283 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1201_ clknet_2_1__leaf_clock _0064_ _0015_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1132_ _0548_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
X_1063_ _0104_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__clkbuf_2
X_0916_ manchester_baby_instance.ram_data_i_23 manchester_baby_instance.ram_data_o_23
+ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or2b_1
X_0847_ _0340_ _0315_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and2b_1
X_0778_ _0204_ _0274_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 _0551_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0632_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
X_0701_ manchester_baby_instance.ram_data_i_14 _0188_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ net9 net2 VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ _0514_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0615_ _0125_ _0126_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ _0496_ _0497_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0366_ _0344_ _0367_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1294_ manchester_baby_instance.ram_data_o_17 _0573_ VGND VGND VPWR VPWR ram_data_io[17]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_33_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0932_ manchester_baby_instance.ram_data_i_25 manchester_baby_instance.ram_data_o_25
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ _0324_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ _0292_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1277_ manchester_baby_instance.ram_data_o_0 _0556_ VGND VGND VPWR VPWR ram_data_io[0]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_14_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ clknet_2_1__leaf_clock _0063_ _0014_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1062_ _0556_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__inv_2
X_1131_ _0548_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
X_0915_ manchester_baby_instance.ram_data_o_23 manchester_baby_instance.ram_data_i_23
+ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__and2b_1
X_0846_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0319_ _0337_ VGND
+ VGND VPWR VPWR _0340_ sky130_fd_sc_hd__and3_1
X_0777_ _0195_ _0185_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 net9 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
X_0700_ _0210_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_0631_ manchester_baby_instance.ram_data_o_12 manchester_baby_instance.ram_data_i_12
+ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__xnor2_2
X_1114_ _0543_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ manchester_baby_instance.ram_data_o_21 _0513_ _0198_ VGND VGND VPWR VPWR _0514_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0829_ _0319_ manchester_baby_instance.ram_data_i_1 _0322_ VGND VGND VPWR VPWR _0323_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0614_ manchester_baby_instance.ram_data_i_1 manchester_baby_instance.ram_data_o_1
+ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__and2b_1
X_1028_ manchester_baby_instance.ram_data_i_23 _0439_ _0498_ VGND VGND VPWR VPWR _0499_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1293_ manchester_baby_instance.ram_data_o_16 _0572_ VGND VGND VPWR VPWR ram_data_io[16]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0862_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0118_ VGND VGND VPWR
+ VPWR _0354_ sky130_fd_sc_hd__or2_1
X_0931_ manchester_baby_instance.ram_data_o_25 manchester_baby_instance.ram_data_i_25
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_15_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0793_ manchester_baby_instance.ram_data_o_4 _0291_ _0251_ VGND VGND VPWR VPWR _0292_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ clknet_2_2__leaf_clock _0100_ _0049_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_18
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1130_ _0548_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
X_1061_ _0104_ _0101_ _0331_ _0526_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nand4b_4
X_0845_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0338_ _0334_ VGND
+ VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21boi_1
X_0914_ _0391_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or2b_1
X_0776_ manchester_baby_instance.ram_data_i_6 _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_0__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_0__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1259_ clknet_2_1__leaf_clock _0083_ _0032_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0630_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1113_ manchester_baby_instance.BASE_1.s_bufferRegs\[0\] net15 VGND VGND VPWR VPWR
+ _0543_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1044_ _0195_ _0505_ _0510_ _0512_ _0106_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0828_ _0320_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0759_ _0261_ _0242_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0613_ manchester_baby_instance.ram_data_o_0 manchester_baby_instance.ram_data_i_0
+ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ _0195_ _0480_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ manchester_baby_instance.ram_data_o_15 _0571_ VGND VGND VPWR VPWR ram_data_io[15]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0861_ _0319_ _0337_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] VGND
+ VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ _0173_ _0397_ _0400_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__o31a_1
X_0792_ _0204_ _0283_ _0288_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1275_ clknet_2_2__leaf_clock _0099_ _0048_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_17
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0525_ VGND VGND
+ VPWR VPWR _0526_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0844_ _0319_ _0337_ manchester_baby_instance.ram_data_o_31 VGND VGND VPWR VPWR _0338_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0775_ manchester_baby_instance.ram_data_i_5 _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__or2_1
X_0913_ manchester_baby_instance.ram_data_i_22 manchester_baby_instance.ram_data_o_22
+ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1258_ clknet_2_0__leaf_clock _0082_ _0031_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_0
+ sky130_fd_sc_hd__dfrtp_1
X_1189_ clknet_2_2__leaf_clock _0052_ _0003_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_21
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1112_ _0542_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1043_ _0388_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_31_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0827_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] manchester_baby_instance.ram_data_i_0
+ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0758_ _0101_ _0103_ _0104_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nand3b_4
XTAP_TAPCELL_ROW_39_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0689_ manchester_baby_instance.ram_data_i_17 _0191_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0612_ manchester_baby_instance.ram_data_o_1 manchester_baby_instance.ram_data_i_1
+ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__or2b_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1026_ _0392_ _0396_ _0495_ _0261_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1009_ manchester_baby_instance.ram_data_i_25 _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput2 net2 VGND VGND VPWR VPWR logisim_clock_tree_0_out sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ manchester_baby_instance.ram_data_o_14 _0570_ VGND VGND VPWR VPWR ram_data_io[14]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0860_ _0316_ _0351_ _0352_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a22o_1
X_0791_ _0195_ _0275_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1274_ clknet_2_2__leaf_clock _0098_ _0047_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_16
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0195_ _0454_ _0462_ _0464_ _0106_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ manchester_baby_instance.ram_data_o_22 manchester_baby_instance.ram_data_i_22
+ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_28_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0843_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] VGND VGND VPWR VPWR
+ _0337_ sky130_fd_sc_hd__buf_2
X_0774_ manchester_baby_instance.ram_data_i_4 _0184_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__or2_1
X_1257_ clknet_2_1__leaf_clock _0081_ _0030_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1188_ clknet_2_2__leaf_clock _0051_ _0002_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_20
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1111_ _0526_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1042_ _0401_ _0494_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0826_ _0319_ manchester_baby_instance.ram_data_i_1 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__xnor2_1
X_0688_ _0200_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_0757_ manchester_baby_instance.ram_data_i_8 _0253_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0611_ _0122_ _0123_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ _0392_ _0495_ _0396_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a21oi_1
X_0809_ _0127_ _0125_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1008_ manchester_baby_instance.ram_data_i_24 _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput3 net3 VGND VGND VPWR VPWR ram_addr_o[0] sky130_fd_sc_hd__clkbuf_4
X_1290_ manchester_baby_instance.ram_data_o_13 _0569_ VGND VGND VPWR VPWR ram_data_io[13]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0790_ manchester_baby_instance.ram_data_i_4 _0184_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1273_ clknet_2_0__leaf_clock _0097_ _0046_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_15
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ _0426_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0842_ _0315_ _0334_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__o21a_1
X_0911_ _0388_ _0389_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__nand2_1
X_0773_ _0112_ _0268_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__xnor2_1
X_1256_ clknet_2_1__leaf_clock _0080_ _0029_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1187_ clknet_2_2__leaf_clock _0050_ _0001_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_19
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0525_ VGND VGND
+ VPWR VPWR _0541_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ manchester_baby_instance.ram_data_i_21 _0504_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nand2_1
X_0825_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] VGND VGND VPWR VPWR
+ _0319_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0756_ _0259_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_0687_ manchester_baby_instance.ram_data_o_18 _0197_ _0199_ VGND VGND VPWR VPWR _0200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_46_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1308_ manchester_baby_instance.ram_data_o_31 _0587_ VGND VGND VPWR VPWR ram_data_io[31]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1239_ ram_data_io[20] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_20
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0610_ manchester_baby_instance.ram_data_o_2 _0118_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_36_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1024_ _0387_ _0401_ _0494_ _0393_ _0386_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a311o_1
XFILLER_0_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0808_ manchester_baby_instance.ram_data_i_1 manchester_baby_instance.ram_data_i_0
+ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nand2_1
X_0739_ _0150_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1007_ manchester_baby_instance.ram_data_i_23 _0439_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput4 net4 VGND VGND VPWR VPWR ram_addr_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_3__leaf_clock sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_9_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ clknet_2_0__leaf_clock _0096_ _0045_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_14
+ sky130_fd_sc_hd__dfrtp_1
X_0987_ _0425_ _0420_ _0423_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0841_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] VGND VGND VPWR VPWR
+ _0335_ sky130_fd_sc_hd__inv_2
X_0772_ _0273_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_0910_ manchester_baby_instance.ram_data_o_20 manchester_baby_instance.ram_data_i_20
+ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1255_ clknet_2_1__leaf_clock _0079_ _0028_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ _0547_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_20_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0509_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0824_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0118_ VGND VGND VPWR
+ VPWR _0318_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ manchester_baby_instance.ram_data_o_9 _0258_ _0251_ VGND VGND VPWR VPWR _0259_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0686_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_39_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1238_ ram_data_io[19] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_19
+ sky130_fd_sc_hd__dlxtn_1
X_1169_ _0555_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
X_1307_ manchester_baby_instance.ram_data_o_30 _0586_ VGND VGND VPWR VPWR ram_data_io[30]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0738_ _0241_ _0243_ _0167_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o21ba_1
X_0807_ _0303_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0669_ _0107_ _0108_ _0177_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ _0479_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput5 net5 VGND VGND VPWR VPWR ram_addr_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_37_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ clknet_2_2__leaf_clock _0095_ _0044_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_13
+ sky130_fd_sc_hd__dfrtp_1
X_0986_ manchester_baby_instance.ram_data_i_28 _0441_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ _0331_ _0311_ _0313_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__and3b_1
X_0771_ manchester_baby_instance.ram_data_o_7 _0272_ _0251_ VGND VGND VPWR VPWR _0273_
+ sky130_fd_sc_hd__mux2_1
X_1254_ clknet_2_1__leaf_clock _0078_ _0027_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1185_ _0547_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ _0447_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0823_ _0311_ _0314_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0754_ _0239_ _0186_ _0255_ _0257_ _0229_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a32o_1
X_0685_ _0106_ _0194_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0198_ sky130_fd_sc_hd__o21a_2
X_1306_ manchester_baby_instance.ram_data_o_29 _0585_ VGND VGND VPWR VPWR ram_data_io[29]
+ sky130_fd_sc_hd__ebufn_8
XFILLER_0_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1099_ _0535_ _0536_ _0537_ _0538_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nand4b_2
X_1237_ ram_data_io[18] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_18
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1168_ _0555_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1022_ _0405_ _0492_ _0389_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_44_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0737_ _0156_ _0157_ _0242_ _0166_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a31oi_2
X_0668_ _0177_ _0107_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0806_ manchester_baby_instance.ram_data_o_2 _0302_ _0251_ VGND VGND VPWR VPWR _0303_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0599_ manchester_baby_instance.ram_data_o_6 manchester_baby_instance.ram_data_i_6
+ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1005_ manchester_baby_instance.ram_data_o_26 _0478_ _0446_ VGND VGND VPWR VPWR _0479_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR ram_addr_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

