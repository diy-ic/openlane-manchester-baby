VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openlane_manchester_baby
  CLASS BLOCK ;
  FOREIGN openlane_manchester_baby ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 160.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.590 10.640 28.190 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.730 10.640 65.330 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.870 10.640 102.470 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.010 10.640 139.610 147.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.380 154.340 31.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 64.380 154.340 65.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 98.380 154.340 99.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 132.380 154.340 133.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.290 10.640 24.890 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.430 10.640 62.030 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.570 10.640 99.170 147.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.710 10.640 136.310 147.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.080 154.340 28.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 61.080 154.340 62.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 95.080 154.340 96.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 129.080 154.340 130.680 ;
    END
  END VPWR
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END clock
  PIN logisim_clock_tree_0_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 156.000 90.530 160.000 ;
    END
  END logisim_clock_tree_0_out
  PIN ram_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 156.000 64.770 160.000 ;
    END
  END ram_addr_o[0]
  PIN ram_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END ram_addr_o[1]
  PIN ram_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END ram_addr_o[2]
  PIN ram_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END ram_addr_o[3]
  PIN ram_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END ram_addr_o[4]
  PIN ram_data_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END ram_data_io[0]
  PIN ram_data_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END ram_data_io[10]
  PIN ram_data_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END ram_data_io[11]
  PIN ram_data_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END ram_data_io[12]
  PIN ram_data_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END ram_data_io[13]
  PIN ram_data_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END ram_data_io[14]
  PIN ram_data_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END ram_data_io[15]
  PIN ram_data_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END ram_data_io[16]
  PIN ram_data_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END ram_data_io[17]
  PIN ram_data_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END ram_data_io[18]
  PIN ram_data_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 54.440 160.000 55.040 ;
    END
  END ram_data_io[19]
  PIN ram_data_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END ram_data_io[1]
  PIN ram_data_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 68.040 160.000 68.640 ;
    END
  END ram_data_io[20]
  PIN ram_data_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 78.240 160.000 78.840 ;
    END
  END ram_data_io[21]
  PIN ram_data_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 85.040 160.000 85.640 ;
    END
  END ram_data_io[22]
  PIN ram_data_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 81.640 160.000 82.240 ;
    END
  END ram_data_io[23]
  PIN ram_data_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 91.840 160.000 92.440 ;
    END
  END ram_data_io[24]
  PIN ram_data_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 98.640 160.000 99.240 ;
    END
  END ram_data_io[25]
  PIN ram_data_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 105.440 160.000 106.040 ;
    END
  END ram_data_io[26]
  PIN ram_data_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 108.840 160.000 109.440 ;
    END
  END ram_data_io[27]
  PIN ram_data_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 102.040 160.000 102.640 ;
    END
  END ram_data_io[28]
  PIN ram_data_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 156.000 103.410 160.000 ;
    END
  END ram_data_io[29]
  PIN ram_data_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END ram_data_io[2]
  PIN ram_data_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 156.000 88.440 160.000 89.040 ;
    END
  END ram_data_io[30]
  PIN ram_data_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 156.000 74.430 160.000 ;
    END
  END ram_data_io[31]
  PIN ram_data_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ram_data_io[3]
  PIN ram_data_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END ram_data_io[4]
  PIN ram_data_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ram_data_io[5]
  PIN ram_data_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END ram_data_io[6]
  PIN ram_data_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END ram_data_io[7]
  PIN ram_data_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END ram_data_io[8]
  PIN ram_data_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END ram_data_io[9]
  PIN ram_rw_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END ram_rw_en_o
  PIN reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END reset_i
  PIN stop_lamp_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 156.000 77.650 160.000 ;
    END
  END stop_lamp_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 154.100 146.965 ;
      LAYER met1 ;
        RECT 4.670 10.640 154.100 147.120 ;
      LAYER met2 ;
        RECT 4.690 155.720 64.210 156.810 ;
        RECT 65.050 155.720 73.870 156.810 ;
        RECT 74.710 155.720 77.090 156.810 ;
        RECT 77.930 155.720 89.970 156.810 ;
        RECT 90.810 155.720 102.850 156.810 ;
        RECT 103.690 155.720 152.170 156.810 ;
        RECT 4.690 4.280 152.170 155.720 ;
        RECT 4.690 3.670 41.670 4.280 ;
        RECT 42.510 3.670 60.990 4.280 ;
        RECT 61.830 3.670 73.870 4.280 ;
        RECT 74.710 3.670 83.530 4.280 ;
        RECT 84.370 3.670 86.750 4.280 ;
        RECT 87.590 3.670 89.970 4.280 ;
        RECT 90.810 3.670 93.190 4.280 ;
        RECT 94.030 3.670 99.630 4.280 ;
        RECT 100.470 3.670 106.070 4.280 ;
        RECT 106.910 3.670 112.510 4.280 ;
        RECT 113.350 3.670 152.170 4.280 ;
      LAYER met3 ;
        RECT 3.990 130.240 156.000 147.045 ;
        RECT 4.400 128.840 156.000 130.240 ;
        RECT 3.990 109.840 156.000 128.840 ;
        RECT 3.990 108.440 155.600 109.840 ;
        RECT 3.990 106.440 156.000 108.440 ;
        RECT 4.400 105.040 155.600 106.440 ;
        RECT 3.990 103.040 156.000 105.040 ;
        RECT 4.400 101.640 155.600 103.040 ;
        RECT 3.990 99.640 156.000 101.640 ;
        RECT 4.400 98.240 155.600 99.640 ;
        RECT 3.990 96.240 156.000 98.240 ;
        RECT 4.400 94.840 156.000 96.240 ;
        RECT 3.990 92.840 156.000 94.840 ;
        RECT 4.400 91.440 155.600 92.840 ;
        RECT 3.990 89.440 156.000 91.440 ;
        RECT 3.990 88.040 155.600 89.440 ;
        RECT 3.990 86.040 156.000 88.040 ;
        RECT 4.400 84.640 155.600 86.040 ;
        RECT 3.990 82.640 156.000 84.640 ;
        RECT 4.400 81.240 155.600 82.640 ;
        RECT 3.990 79.240 156.000 81.240 ;
        RECT 4.400 77.840 155.600 79.240 ;
        RECT 3.990 75.840 156.000 77.840 ;
        RECT 4.400 74.440 156.000 75.840 ;
        RECT 3.990 72.440 156.000 74.440 ;
        RECT 4.400 71.040 156.000 72.440 ;
        RECT 3.990 69.040 156.000 71.040 ;
        RECT 4.400 67.640 155.600 69.040 ;
        RECT 3.990 62.240 156.000 67.640 ;
        RECT 4.400 60.840 156.000 62.240 ;
        RECT 3.990 55.440 156.000 60.840 ;
        RECT 4.400 54.040 155.600 55.440 ;
        RECT 3.990 48.640 156.000 54.040 ;
        RECT 4.400 47.240 156.000 48.640 ;
        RECT 3.990 41.840 156.000 47.240 ;
        RECT 4.400 40.440 156.000 41.840 ;
        RECT 3.990 10.715 156.000 40.440 ;
  END
END openlane_manchester_baby
END LIBRARY

