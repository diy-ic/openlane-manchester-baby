magic
tech sky130A
magscale 1 2
timestamp 1700924124
<< obsli1 >>
rect 1104 2159 30820 29393
<< obsm1 >>
rect 934 2128 30820 29424
<< metal2 >>
rect 12898 31200 12954 32000
rect 14830 31200 14886 32000
rect 15474 31200 15530 32000
rect 18050 31200 18106 32000
rect 20626 31200 20682 32000
rect 8390 0 8446 800
rect 12254 0 12310 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
<< obsm2 >>
rect 938 31144 12842 31362
rect 13010 31144 14774 31362
rect 14942 31144 15418 31362
rect 15586 31144 17994 31362
rect 18162 31144 20570 31362
rect 20738 31144 30434 31362
rect 938 856 30434 31144
rect 938 734 8334 856
rect 8502 734 12198 856
rect 12366 734 14774 856
rect 14942 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18638 856
rect 18806 734 19926 856
rect 20094 734 21214 856
rect 21382 734 22502 856
rect 22670 734 30434 856
<< metal3 >>
rect 0 25848 800 25968
rect 31200 21768 32000 21888
rect 0 21088 800 21208
rect 31200 21088 32000 21208
rect 0 20408 800 20528
rect 31200 20408 32000 20528
rect 0 19728 800 19848
rect 31200 19728 32000 19848
rect 0 19048 800 19168
rect 0 18368 800 18488
rect 31200 18368 32000 18488
rect 31200 17688 32000 17808
rect 0 17008 800 17128
rect 31200 17008 32000 17128
rect 0 16328 800 16448
rect 31200 16328 32000 16448
rect 0 15648 800 15768
rect 31200 15648 32000 15768
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 31200 13608 32000 13728
rect 0 12248 800 12368
rect 0 10888 800 11008
rect 31200 10888 32000 11008
rect 0 9528 800 9648
rect 0 8168 800 8288
<< obsm3 >>
rect 798 26048 31200 29409
rect 880 25768 31200 26048
rect 798 21968 31200 25768
rect 798 21688 31120 21968
rect 798 21288 31200 21688
rect 880 21008 31120 21288
rect 798 20608 31200 21008
rect 880 20328 31120 20608
rect 798 19928 31200 20328
rect 880 19648 31120 19928
rect 798 19248 31200 19648
rect 880 18968 31200 19248
rect 798 18568 31200 18968
rect 880 18288 31120 18568
rect 798 17888 31200 18288
rect 798 17608 31120 17888
rect 798 17208 31200 17608
rect 880 16928 31120 17208
rect 798 16528 31200 16928
rect 880 16248 31120 16528
rect 798 15848 31200 16248
rect 880 15568 31120 15848
rect 798 15168 31200 15568
rect 880 14888 31200 15168
rect 798 14488 31200 14888
rect 880 14208 31200 14488
rect 798 13808 31200 14208
rect 880 13528 31120 13808
rect 798 12448 31200 13528
rect 880 12168 31200 12448
rect 798 11088 31200 12168
rect 880 10808 31120 11088
rect 798 9728 31200 10808
rect 880 9448 31200 9728
rect 798 8368 31200 9448
rect 880 8088 31200 8368
rect 798 2143 31200 8088
<< metal4 >>
rect 4658 2128 4978 29424
rect 5318 2128 5638 29424
rect 12086 2128 12406 29424
rect 12746 2128 13066 29424
rect 19514 2128 19834 29424
rect 20174 2128 20494 29424
rect 26942 2128 27262 29424
rect 27602 2128 27922 29424
<< metal5 >>
rect 1056 26476 30868 26796
rect 1056 25816 30868 26136
rect 1056 19676 30868 19996
rect 1056 19016 30868 19336
rect 1056 12876 30868 13196
rect 1056 12216 30868 12536
rect 1056 6076 30868 6396
rect 1056 5416 30868 5736
<< labels >>
rlabel metal4 s 5318 2128 5638 29424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12746 2128 13066 29424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 20174 2128 20494 29424 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27602 2128 27922 29424 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6076 30868 6396 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12876 30868 13196 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 19676 30868 19996 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 26476 30868 26796 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4658 2128 4978 29424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12086 2128 12406 29424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19514 2128 19834 29424 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26942 2128 27262 29424 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5416 30868 5736 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 12216 30868 12536 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 19016 30868 19336 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 25816 30868 26136 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 25848 800 25968 6 clock
port 3 nsew signal input
rlabel metal2 s 18050 31200 18106 32000 6 logisim_clock_tree_0_out
port 4 nsew signal output
rlabel metal2 s 12898 31200 12954 32000 6 ram_addr_o[0]
port 5 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 ram_addr_o[1]
port 6 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 ram_addr_o[2]
port 7 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 ram_addr_o[3]
port 8 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 ram_addr_o[4]
port 9 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 ram_data_io[0]
port 10 nsew signal bidirectional
rlabel metal2 s 12254 0 12310 800 6 ram_data_io[10]
port 11 nsew signal bidirectional
rlabel metal2 s 18050 0 18106 800 6 ram_data_io[11]
port 12 nsew signal bidirectional
rlabel metal2 s 17406 0 17462 800 6 ram_data_io[12]
port 13 nsew signal bidirectional
rlabel metal2 s 18694 0 18750 800 6 ram_data_io[13]
port 14 nsew signal bidirectional
rlabel metal2 s 16762 0 16818 800 6 ram_data_io[14]
port 15 nsew signal bidirectional
rlabel metal2 s 14830 0 14886 800 6 ram_data_io[15]
port 16 nsew signal bidirectional
rlabel metal2 s 19982 0 20038 800 6 ram_data_io[16]
port 17 nsew signal bidirectional
rlabel metal2 s 21270 0 21326 800 6 ram_data_io[17]
port 18 nsew signal bidirectional
rlabel metal2 s 22558 0 22614 800 6 ram_data_io[18]
port 19 nsew signal bidirectional
rlabel metal3 s 31200 10888 32000 11008 6 ram_data_io[19]
port 20 nsew signal bidirectional
rlabel metal3 s 0 14968 800 15088 6 ram_data_io[1]
port 21 nsew signal bidirectional
rlabel metal3 s 31200 13608 32000 13728 6 ram_data_io[20]
port 22 nsew signal bidirectional
rlabel metal3 s 31200 15648 32000 15768 6 ram_data_io[21]
port 23 nsew signal bidirectional
rlabel metal3 s 31200 17008 32000 17128 6 ram_data_io[22]
port 24 nsew signal bidirectional
rlabel metal3 s 31200 16328 32000 16448 6 ram_data_io[23]
port 25 nsew signal bidirectional
rlabel metal3 s 31200 18368 32000 18488 6 ram_data_io[24]
port 26 nsew signal bidirectional
rlabel metal3 s 31200 19728 32000 19848 6 ram_data_io[25]
port 27 nsew signal bidirectional
rlabel metal3 s 31200 21088 32000 21208 6 ram_data_io[26]
port 28 nsew signal bidirectional
rlabel metal3 s 31200 21768 32000 21888 6 ram_data_io[27]
port 29 nsew signal bidirectional
rlabel metal3 s 31200 20408 32000 20528 6 ram_data_io[28]
port 30 nsew signal bidirectional
rlabel metal2 s 20626 31200 20682 32000 6 ram_data_io[29]
port 31 nsew signal bidirectional
rlabel metal3 s 0 15648 800 15768 6 ram_data_io[2]
port 32 nsew signal bidirectional
rlabel metal3 s 31200 17688 32000 17808 6 ram_data_io[30]
port 33 nsew signal bidirectional
rlabel metal2 s 14830 31200 14886 32000 6 ram_data_io[31]
port 34 nsew signal bidirectional
rlabel metal3 s 0 16328 800 16448 6 ram_data_io[3]
port 35 nsew signal bidirectional
rlabel metal3 s 0 13608 800 13728 6 ram_data_io[4]
port 36 nsew signal bidirectional
rlabel metal3 s 0 12248 800 12368 6 ram_data_io[5]
port 37 nsew signal bidirectional
rlabel metal3 s 0 10888 800 11008 6 ram_data_io[6]
port 38 nsew signal bidirectional
rlabel metal3 s 0 9528 800 9648 6 ram_data_io[7]
port 39 nsew signal bidirectional
rlabel metal3 s 0 8168 800 8288 6 ram_data_io[8]
port 40 nsew signal bidirectional
rlabel metal2 s 8390 0 8446 800 6 ram_data_io[9]
port 41 nsew signal bidirectional
rlabel metal3 s 0 21088 800 21208 6 ram_rw_en_o
port 42 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 reset_i
port 43 nsew signal input
rlabel metal2 s 15474 31200 15530 32000 6 stop_lamp_o
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32000 32000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2401382
string GDS_FILE /openlane/designs/openlane-manchester-baby/runs/RUN_2023.11.25_14.53.08/results/signoff/openlane_manchester_baby.magic.gds
string GDS_START 535932
<< end >>

