* NGSPICE file created from openlane_manchester_baby.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt openlane_manchester_baby VGND VPWR clock ram_addr_o[0] ram_addr_o[1] ram_addr_o[2]
+ ram_addr_o[3] ram_addr_o[4] ram_data_io[0] ram_data_io[10] ram_data_io[11] ram_data_io[12]
+ ram_data_io[13] ram_data_io[14] ram_data_io[15] ram_data_io[16] ram_data_io[17]
+ ram_data_io[18] ram_data_io[19] ram_data_io[1] ram_data_io[20] ram_data_io[21] ram_data_io[22]
+ ram_data_io[23] ram_data_io[24] ram_data_io[25] ram_data_io[26] ram_data_io[27]
+ ram_data_io[28] ram_data_io[29] ram_data_io[2] ram_data_io[30] ram_data_io[31] ram_data_io[3]
+ ram_data_io[4] ram_data_io[5] ram_data_io[6] ram_data_io[7] ram_data_io[8] ram_data_io[9]
+ ram_rw_en_o reset_i stop_lamp_o
XTAP_TAPCELL_ROW_37_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ _0639_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ _0207_ _0210_ _0377_ _0378_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o31a_1
X_1468_ manchester_baby_instance.ram_data_o_2 net11 VGND VGND VPWR VPWR ram_data_io[2]
+ sky130_fd_sc_hd__dlxtp_1
X_1399_ clknet_3_6__leaf_clock _0086_ _0040_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ _0199_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1322_ manchester_baby_instance.BASE_0.s_countReg\[10\] _0619_ VGND VGND VPWR VPWR
+ _0659_ sky130_fd_sc_hd__and2_1
X_1253_ _0640_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1184_ _0590_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_62_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0968_ manchester_baby_instance.ram_data_i_20 manchester_baby_instance.ram_data_i_21
+ _0399_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0899_ _0324_ _0331_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ _0253_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0753_ _0192_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
X_0684_ manchester_baby_instance.ram_data_i_2 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1236_ _0634_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
X_1305_ _0648_ net45 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1098_ _0515_ manchester_baby_instance.ram_data_o_16 _0470_ VGND VGND VPWR VPWR _0516_
+ sky130_fd_sc_hd__mux2_1
X_1167_ _0572_ _0573_ _0575_ _0484_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_356 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1021_ _0448_ manchester_baby_instance.ram_data_o_26 _0414_ VGND VGND VPWR VPWR _0449_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0805_ _0132_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0736_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0131_ _0180_ _0130_
+ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1219_ manchester_baby_instance.BASE_0.s_countReg\[10\] manchester_baby_instance.BASE_0.s_countReg\[11\]
+ net29 _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__or4_4
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold52 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] VGND VGND VPWR VPWR
+ net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 _0095_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1004_ _0376_ _0371_ _0374_ _0377_ _0386_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_32_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0719_ _0151_ _0155_ _0159_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput7 net15 VGND VGND VPWR VPWR ram_rw_en_o sky130_fd_sc_hd__buf_2
XFILLER_0_53_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1484_ manchester_baby_instance.ram_data_o_18 net13 VGND VGND VPWR VPWR ram_data_io[18]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ _0412_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_4
X_1398_ clknet_3_6__leaf_clock _0085_ _0039_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1467_ manchester_baby_instance.ram_data_o_1 net11 VGND VGND VPWR VPWR ram_data_io[1]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_19_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1321_ manchester_baby_instance.BASE_0.s_countReg\[10\] _0619_ VGND VGND VPWR VPWR
+ _0658_ sky130_fd_sc_hd__nor2_1
X_1252_ _0640_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
X_1183_ _0589_ manchester_baby_instance.ram_data_o_5 _0538_ VGND VGND VPWR VPWR _0590_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0967_ manchester_baby_instance.ram_data_i_16 manchester_baby_instance.ram_data_i_17
+ manchester_baby_instance.ram_data_i_18 manchester_baby_instance.ram_data_i_19 VGND
+ VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ manchester_baby_instance.ram_data_i_16 manchester_baby_instance.ram_data_o_16
+ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0752_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] manchester_baby_instance.ram_data_i_14
+ _0190_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ manchester_baby_instance.ram_data_o_8 manchester_baby_instance.ram_data_i_8
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__and2b_1
X_0683_ _0124_ _0127_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1235_ net18 net19 VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__and2b_1
X_1304_ net20 manchester_baby_instance.BASE_0.s_countReg\[1\] net44 VGND VGND VPWR
+ VPWR _0649_ sky130_fd_sc_hd__o21ai_1
X_1166_ _0395_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1097_ _0484_ _0513_ _0514_ _0424_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1020_ _0416_ _0439_ _0446_ _0447_ _0421_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0735_ _0134_ _0158_ _0175_ _0129_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a221o_1
X_0804_ _0236_ _0233_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1218_ manchester_baby_instance.BASE_0.s_countReg\[7\] manchester_baby_instance.BASE_0.s_countReg\[8\]
+ net49 _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or4_4
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1149_ _0544_ _0262_ _0261_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_47_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold20 manchester_baby_instance.BASE_0.s_countReg\[17\] VGND VGND VPWR VPWR net36
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _0107_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 manchester_baby_instance.ram_data_o_0 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0406_ _0432_ _0421_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0718_ manchester_baby_instance.ram_data_i_3 _0158_ _0164_ _0148_ VGND VGND VPWR
+ VPWR _0165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR stop_lamp_o sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_33_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1483_ manchester_baby_instance.ram_data_o_17 net13 VGND VGND VPWR VPWR ram_data_io[17]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ _0415_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1397_ clknet_3_6__leaf_clock _0084_ _0038_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1466_ manchester_baby_instance.ram_data_o_0 net12 VGND VGND VPWR VPWR ram_data_io[0]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1320_ _0619_ net50 manchester_baby_instance.BASE_0.s_tickNext VGND VGND VPWR VPWR
+ _0102_ sky130_fd_sc_hd__a21oi_1
X_1251_ _0640_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
X_1182_ _0416_ _0586_ _0588_ _0429_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_20_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0966_ _0395_ _0396_ _0397_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__and4_1
X_0897_ manchester_baby_instance.ram_data_i_15 _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1449_ ram_data_io[15] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_15
+ sky130_fd_sc_hd__dlxtn_2
XTAP_TAPCELL_ROW_53_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0751_ _0191_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ manchester_baby_instance.ram_data_o_9 manchester_baby_instance.ram_data_i_9
+ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0682_ _0124_ _0129_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0130_ sky130_fd_sc_hd__o21a_1
X_1303_ manchester_baby_instance.BASE_0.s_countReg\[0\] manchester_baby_instance.BASE_0.s_countReg\[1\]
+ net44 VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1234_ _0633_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_1165_ manchester_baby_instance.ram_data_i_6 _0392_ _0393_ manchester_baby_instance.ram_data_i_7
+ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a31o_1
X_1096_ _0461_ _0333_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0949_ manchester_baby_instance.ram_data_o_31 manchester_baby_instance.ram_data_i_31
+ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_325 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0734_ _0148_ _0139_ _0176_ _0178_ _0150_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__a32o_1
X_0803_ _0132_ manchester_baby_instance.ram_data_o_2 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__xor2_2
Xfanout9 net16 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1217_ manchester_baby_instance.BASE_0.s_countReg\[4\] manchester_baby_instance.BASE_0.s_countReg\[5\]
+ manchester_baby_instance.BASE_0.s_countReg\[6\] _0617_ VGND VGND VPWR VPWR _0618_
+ sky130_fd_sc_hd__or4_4
X_1148_ _0559_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_1079_ _0499_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold21 _0110_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 manchester_baby_instance.BASE_0.s_countReg\[24\] VGND VGND VPWR VPWR net59
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 manchester_baby_instance.CIRCUIT_0.IR.q\[0\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 _0663_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1002_ manchester_baby_instance.ram_data_i_28 _0404_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ _0142_ _0163_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1482_ manchester_baby_instance.ram_data_o_16 net10 VGND VGND VPWR VPWR ram_data_io[16]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ _0410_ manchester_baby_instance.ram_data_o_31 _0414_ VGND VGND VPWR VPWR _0415_
+ sky130_fd_sc_hd__mux2_1
X_1465_ ram_data_io[31] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_31
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1396_ clknet_3_1__leaf_clock _0083_ _0037_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_250 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ _0640_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
X_1181_ _0578_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_334 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_364 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ manchester_baby_instance.ram_data_i_15 manchester_baby_instance.ram_data_i_14
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__and2_1
X_0896_ manchester_baby_instance.ram_data_o_15 VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__inv_2
X_1448_ ram_data_io[14] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_14
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ clknet_3_5__leaf_clock _0066_ _0020_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_19
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0681_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0128_ VGND VGND
+ VPWR VPWR _0129_ sky130_fd_sc_hd__nor2_2
X_0750_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.ram_data_i_15
+ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1233_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0632_ VGND VGND VPWR VPWR _0633_
+ sky130_fd_sc_hd__and4b_1
X_1302_ net17 net61 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1095_ manchester_baby_instance.ram_data_i_16 _0399_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__xnor2_1
X_1164_ _0213_ _0225_ _0571_ _0386_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0948_ _0207_ _0210_ _0377_ _0378_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0879_ _0306_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0802_ _0232_ manchester_baby_instance.ram_data_o_0 _0233_ _0234_ VGND VGND VPWR
+ VPWR _0235_ sky130_fd_sc_hd__o22a_2
XFILLER_0_8_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0733_ _0153_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1216_ manchester_baby_instance.BASE_0.s_countReg\[0\] manchester_baby_instance.BASE_0.s_countReg\[1\]
+ manchester_baby_instance.BASE_0.s_countReg\[2\] manchester_baby_instance.BASE_0.s_countReg\[3\]
+ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or4_4
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1147_ _0558_ manchester_baby_instance.ram_data_o_10 _0538_ VGND VGND VPWR VPWR _0559_
+ sky130_fd_sc_hd__mux2_1
X_1078_ _0498_ manchester_baby_instance.ram_data_o_19 _0470_ VGND VGND VPWR VPWR _0499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold22 manchester_baby_instance.BASE_0.s_countReg\[19\] VGND VGND VPWR VPWR net38
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 _0653_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold44 net8 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 manchester_baby_instance.BASE_0.s_countReg\[9\] VGND VGND VPWR VPWR net49
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 manchester_baby_instance.CIRCUIT_0.IR.q\[1\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ _0431_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0716_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1481_ manchester_baby_instance.ram_data_o_15 net10 VGND VGND VPWR VPWR ram_data_io[15]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_270 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0981_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1395_ clknet_3_1__leaf_clock _0082_ _0036_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1464_ ram_data_io[30] net12 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_30
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clock clock VGND VGND VPWR VPWR clknet_0_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1180_ manchester_baby_instance.ram_data_i_4 _0392_ manchester_baby_instance.ram_data_i_5
+ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ manchester_baby_instance.ram_data_i_13 manchester_baby_instance.ram_data_i_12
+ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0895_ _0326_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__and2_1
X_1447_ ram_data_io[13] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_13
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1378_ clknet_3_5__leaf_clock _0065_ _0019_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_18
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0680_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__or2_1
X_1232_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0631_ VGND VGND
+ VPWR VPWR _0632_ sky130_fd_sc_hd__nor2_1
X_1301_ net20 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1094_ _0512_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_1163_ _0225_ _0571_ _0213_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0947_ _0203_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ _0308_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_21_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0801_ _0134_ manchester_baby_instance.ram_data_o_1 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0732_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] manchester_baby_instance.ram_data_o_31
+ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] VGND VGND VPWR VPWR _0177_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1215_ net59 VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__inv_2
X_1146_ _0484_ _0555_ _0557_ _0424_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1077_ _0412_ _0494_ _0495_ _0497_ _0429_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__a32o_1
Xhold23 _0669_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 _0657_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 manchester_baby_instance.CIRCUIT_0.IR.q\[4\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 manchester_baby_instance.BASE_0.s_countReg\[1\] VGND VGND VPWR VPWR net61
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0099_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1000_ _0430_ manchester_baby_instance.ram_data_o_29 _0414_ VGND VGND VPWR VPWR _0431_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0715_ net68 _0131_ _0162_ _0130_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1129_ _0542_ manchester_baby_instance.ram_data_o_12 _0538_ VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ manchester_baby_instance.ram_data_o_14 net12 VGND VGND VPWR VPWR ram_data_io[14]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0412_ _0388_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0413_ sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_57_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1394_ clknet_3_1__leaf_clock _0081_ _0035_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1463_ ram_data_io[29] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_29
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_54_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0963_ manchester_baby_instance.ram_data_i_8 manchester_baby_instance.ram_data_i_9
+ manchester_baby_instance.ram_data_i_10 manchester_baby_instance.ram_data_i_11 VGND
+ VGND VPWR VPWR _0396_ sky130_fd_sc_hd__and4_1
X_0894_ _0324_ _0325_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1377_ clknet_3_4__leaf_clock _0064_ _0018_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_17
+ sky130_fd_sc_hd__dfrtp_1
X_1446_ ram_data_io[12] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_12
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_61_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1300_ _0647_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_1231_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_2__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_2__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1162_ _0216_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2b_1
X_1093_ _0511_ manchester_baby_instance.ram_data_o_17 _0470_ VGND VGND VPWR VPWR _0512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0946_ _0199_ _0202_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__nand2_1
X_0877_ manchester_baby_instance.ram_data_o_19 _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ clknet_3_2__leaf_clock net33 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0731_ _0135_ _0137_ _0136_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a21bo_1
X_0800_ manchester_baby_instance.ram_data_o_1 _0134_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1214_ net69 _0614_ _0615_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR VPWR
+ _0047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1145_ _0546_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1076_ _0309_ _0496_ _0482_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a21o_1
X_0929_ _0209_ _0360_ manchester_baby_instance.ram_data_o_26 _0361_ VGND VGND VPWR
+ VPWR _0362_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_15_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 manchester_baby_instance.BASE_0.s_countReg\[18\] VGND VGND VPWR VPWR net62
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 manchester_baby_instance.BASE_0.s_countReg\[25\] VGND VGND VPWR VPWR net40
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 manchester_baby_instance.CIRCUIT_0.IR.q\[2\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 manchester_baby_instance.BASE_0.s_countReg\[12\] VGND VGND VPWR VPWR net29
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0714_ _0149_ _0157_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1128_ _0484_ _0540_ _0541_ _0424_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__a22o_1
X_1059_ manchester_baby_instance.ram_data_i_18 manchester_baby_instance.ram_data_i_19
+ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1462_ ram_data_io[28] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_28
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1393_ clknet_3_6__leaf_clock _0080_ _0034_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ _0324_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2_1
X_0962_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_2
X_1445_ ram_data_io[11] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_11
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ clknet_3_4__leaf_clock _0063_ _0017_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_16
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1230_ _0630_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_tickNext sky130_fd_sc_hd__inv_4
X_1092_ _0416_ _0508_ _0510_ _0429_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1161_ _0231_ _0242_ _0244_ _0224_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0945_ manchester_baby_instance.ram_data_o_28 _0204_ _0206_ VGND VGND VPWR VPWR _0378_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ manchester_baby_instance.ram_data_i_19 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__inv_2
X_1428_ clknet_3_3__leaf_clock _0114_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1359_ _0639_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0730_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_12_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1213_ manchester_baby_instance.ram_data_o_0 _0389_ _0414_ VGND VGND VPWR VPWR _0615_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1144_ _0252_ _0281_ _0545_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and3_1
X_1075_ manchester_baby_instance.ram_data_i_18 _0481_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0928_ manchester_baby_instance.ram_data_i_26 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0859_ manchester_baby_instance.ram_data_o_23 manchester_baby_instance.ram_data_i_23
+ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold47 manchester_baby_instance.BASE_0.s_tickReg VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _0113_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 manchester_baby_instance.BASE_0.s_countReg\[16\] VGND VGND VPWR VPWR net74
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0661_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0713_ manchester_baby_instance.ram_data_i_4 _0158_ _0160_ VGND VGND VPWR VPWR _0161_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1058_ manchester_baby_instance.ram_data_i_15 manchester_baby_instance.ram_data_i_16
+ manchester_baby_instance.ram_data_i_17 _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__and4_1
X_1127_ _0277_ _0518_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1461_ ram_data_io[27] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_27
+ sky130_fd_sc_hd__dlxtn_1
X_1392_ clknet_3_6__leaf_clock _0079_ _0033_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ manchester_baby_instance.ram_data_i_6 manchester_baby_instance.ram_data_i_7
+ _0392_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0892_ manchester_baby_instance.ram_data_o_17 manchester_baby_instance.ram_data_i_17
+ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__xnor2_1
X_1444_ ram_data_io[10] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_10
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_10_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1375_ clknet_3_5__leaf_clock _0062_ _0016_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_15
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1160_ _0569_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
X_1091_ _0502_ _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0944_ _0371_ _0374_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0305_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1427_ clknet_3_2__leaf_clock net52 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_1358_ _0639_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
X_1289_ _0643_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1212_ _0232_ _0424_ _0414_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ _0550_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nand2_1
X_1074_ _0316_ _0317_ _0320_ _0493_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_55_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0927_ manchester_baby_instance.ram_data_i_27 manchester_baby_instance.ram_data_o_27
+ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0789_ _0220_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__nand2_1
X_0858_ manchester_baby_instance.ram_data_o_22 manchester_baby_instance.ram_data_i_22
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold59 manchester_baby_instance.CIRCUIT_0.IR.q\[3\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 manchester_baby_instance.BASE_0.s_countReg\[4\] VGND VGND VPWR VPWR net42
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_34_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0712_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ _0155_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__and4b_1
XFILLER_0_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1126_ manchester_baby_instance.ram_data_i_12 _0479_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__xnor2_1
X_1057_ manchester_baby_instance.ram_data_i_14 manchester_baby_instance.ram_data_i_13
+ manchester_baby_instance.ram_data_i_12 _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ _0525_ manchester_baby_instance.ram_data_o_15 _0470_ VGND VGND VPWR VPWR _0526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1460_ ram_data_io[26] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_26
+ sky130_fd_sc_hd__dlxtn_2
X_1391_ clknet_3_7__leaf_clock _0078_ _0032_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_31
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_35_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0960_ manchester_baby_instance.ram_data_i_4 manchester_baby_instance.ram_data_i_5
+ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0891_ manchester_baby_instance.ram_data_o_16 manchester_baby_instance.ram_data_i_16
+ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ clknet_3_4__leaf_clock _0061_ _0015_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_14
+ sky130_fd_sc_hd__dfrtp_1
X_1443_ ram_data_io[9] net9 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_9
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1090_ manchester_baby_instance.ram_data_i_17 _0501_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0943_ _0210_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0874_ manchester_baby_instance.ram_data_i_20 manchester_baby_instance.ram_data_o_20
+ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1357_ _0639_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
X_1426_ clknet_3_2__leaf_clock _0112_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_1288_ _0643_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1211_ _0613_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_1142_ manchester_baby_instance.ram_data_i_10 _0549_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1073_ _0320_ _0493_ _0316_ _0317_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ _0353_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0857_ _0279_ _0284_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold38 _0098_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 _0652_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ clknet_3_2__leaf_clock net46 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_0788_ manchester_baby_instance.ram_data_o_3 manchester_baby_instance.ram_data_i_3
+ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2b_2
Xhold49 _0660_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ manchester_baby_instance.ram_data_o_31 _0150_ _0129_ VGND VGND VPWR VPWR _0159_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1125_ _0539_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1056_ _0395_ _0396_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0909_ _0326_ _0341_ _0327_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1108_ _0424_ _0521_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a21o_1
X_1039_ _0339_ _0463_ _0301_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ clknet_3_7__leaf_clock _0077_ _0031_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_30
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_5__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0316_ _0317_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1442_ ram_data_io[8] net9 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_8
+ sky130_fd_sc_hd__dlxtn_1
X_1373_ clknet_3_4__leaf_clock _0060_ _0014_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_13
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_18_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ _0208_ _0209_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0873_ _0304_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__xor2_1
X_1425_ clknet_3_2__leaf_clock _0111_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1356_ _0639_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
X_1287_ _0643_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1210_ _0612_ manchester_baby_instance.ram_data_o_1 _0413_ VGND VGND VPWR VPWR _0613_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1141_ _0553_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
X_1072_ _0342_ _0492_ _0322_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0925_ _0356_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__nand2_1
X_0787_ manchester_baby_instance.ram_data_i_4 manchester_baby_instance.ram_data_o_4
+ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__xor2_2
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0856_ _0266_ _0271_ _0286_ _0287_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o311a_1
Xhold39 manchester_baby_instance.BASE_1.s_counterValue VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 _0115_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1408_ clknet_3_2__leaf_clock _0094_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold28 manchester_baby_instance.BASE_0.s_countReg\[2\] VGND VGND VPWR VPWR net44
+ sky130_fd_sc_hd__dlygate4sd3_1
X_1339_ _0622_ _0623_ net62 VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0710_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0124_ _0125_ VGND VGND VPWR
+ VPWR _0158_ sky130_fd_sc_hd__and3b_1
XFILLER_0_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1124_ _0537_ manchester_baby_instance.ram_data_o_13 _0538_ VGND VGND VPWR VPWR _0539_
+ sky130_fd_sc_hd__mux2_1
X_1055_ _0306_ _0477_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0839_ manchester_baby_instance.ram_data_i_13 manchester_baby_instance.ram_data_o_13
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0908_ manchester_baby_instance.ram_data_i_15 _0329_ _0332_ VGND VGND VPWR VPWR _0341_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1107_ _0399_ _0523_ _0484_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__o21a_1
X_1038_ _0312_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1441_ ram_data_io[7] net9 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_7
+ sky130_fd_sc_hd__dlxtn_1
X_1372_ clknet_3_1__leaf_clock _0059_ _0013_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_12
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0941_ _0363_ _0367_ _0370_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0872_ manchester_baby_instance.ram_data_o_20 manchester_baby_instance.ram_data_i_20
+ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and2b_1
X_1355_ _0639_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
X_1424_ clknet_3_2__leaf_clock net37 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1286_ _0643_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1140_ _0552_ manchester_baby_instance.ram_data_o_11 _0538_ VGND VGND VPWR VPWR _0553_
+ sky130_fd_sc_hd__mux2_1
X_1071_ _0461_ _0334_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__or2_1
X_0924_ _0292_ _0355_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0786_ _0217_ manchester_baby_instance.ram_data_o_4 _0218_ VGND VGND VPWR VPWR _0219_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0855_ _0264_ _0265_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__or2_1
X_1338_ net62 _0622_ _0623_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__or3_1
Xhold18 manchester_baby_instance.BASE_0.s_countReg\[15\] VGND VGND VPWR VPWR net34
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold29 _0649_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ clknet_3_2__leaf_clock _0093_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_1269_ _0641_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1123_ _0413_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__clkbuf_4
X_1054_ _0337_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0907_ _0294_ _0299_ _0302_ _0339_ _0295_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0769_ _0200_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nor2_1
X_0838_ _0269_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1106_ manchester_baby_instance.ram_data_i_14 _0522_ manchester_baby_instance.ram_data_i_15
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1037_ _0461_ _0335_ _0344_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ clknet_3_4__leaf_clock _0058_ _0012_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_11
+ sky130_fd_sc_hd__dfrtp_1
X_1440_ ram_data_io[6] net9 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_6
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_61_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout10 net16 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0940_ _0362_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0871_ _0298_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nor2_1
X_1354_ _0630_ _0675_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__nand2_1
X_1423_ clknet_3_2__leaf_clock _0109_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_1285_ _0643_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0491_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
X_0923_ _0292_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0854_ _0264_ _0265_ _0269_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0785_ manchester_baby_instance.ram_data_o_5 manchester_baby_instance.ram_data_i_5
+ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1406_ clknet_3_3__leaf_clock _0092_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_counterValue
+ sky130_fd_sc_hd__dfxtp_1
X_1337_ net36 _0665_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__xor2_1
Xhold19 _0664_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
X_1268_ _0641_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1199_ _0235_ _0237_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1122_ _0533_ _0534_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_48_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1053_ _0311_ _0462_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0837_ _0267_ _0268_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ _0304_ _0305_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0699_ manchester_baby_instance.ram_data_i_4 _0145_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__nor2_1
X_0768_ manchester_baby_instance.ram_data_i_30 manchester_baby_instance.ram_data_o_30
+ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_39_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1105_ _0395_ _0396_ _0397_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1036_ _0280_ _0290_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1019_ manchester_baby_instance.ram_data_i_26 _0403_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1370_ clknet_3_1__leaf_clock _0057_ _0011_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_10
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1499_ clknet_3_6__leaf_clock _0000_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.Acc.tick
+ sky130_fd_sc_hd__dfxtp_1
Xfanout11 net16 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ manchester_baby_instance.ram_data_i_21 manchester_baby_instance.ram_data_o_21
+ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ clknet_3_2__leaf_clock _0108_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_50_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ net40 _0628_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__nand2_1
X_1284_ _0643_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0999_ _0424_ _0427_ _0428_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0922_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0853_ _0272_ _0273_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a21bo_1
X_1405_ clknet_3_6__leaf_clock net19 VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_0784_ manchester_baby_instance.ram_data_i_4 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1336_ _0665_ _0666_ _0630_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o21a_1
X_1198_ _0602_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
Xinput1 reset_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_26_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1267_ _0641_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1052_ _0475_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_1121_ _0522_ _0535_ _0421_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0767_ manchester_baby_instance.ram_data_o_30 manchester_baby_instance.ram_data_i_30
+ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_31_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0836_ _0267_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__or2_1
X_0905_ _0304_ _0305_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o21a_1
X_0698_ manchester_baby_instance.ram_data_i_4 _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1319_ manchester_baby_instance.BASE_0.s_countReg\[7\] manchester_baby_instance.BASE_0.s_countReg\[8\]
+ _0618_ net49 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_39_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ _0460_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1104_ _0266_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__xnor2_1
X_0819_ _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _0369_ _0438_ _0372_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1498_ clknet_3_6__leaf_clock net18 VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.GATES_13.input1
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout12 net16 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421_ clknet_3_2__leaf_clock net58 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_1352_ _0616_ _0627_ _0674_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__o21ai_1
X_1283_ _0643_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0998_ _0388_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0921_ manchester_baby_instance.ram_data_o_24 manchester_baby_instance.ram_data_i_24
+ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_23_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0783_ _0214_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__xnor2_2
X_0852_ _0272_ _0273_ _0275_ _0276_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1404_ manchester_baby_instance.CIRCUIT_0.GATES_13.result _0091_ VGND VGND VPWR VPWR
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] sky130_fd_sc_hd__dfxtp_1
X_1335_ net74 _0622_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ _0601_ manchester_baby_instance.ram_data_o_3 _0413_ VGND VGND VPWR VPWR _0602_
+ sky130_fd_sc_hd__mux2_1
X_1266_ _0641_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1051_ _0474_ manchester_baby_instance.ram_data_o_22 _0470_ VGND VGND VPWR VPWR _0475_
+ sky130_fd_sc_hd__mux2_1
X_1120_ manchester_baby_instance.ram_data_i_12 _0479_ manchester_baby_instance.ram_data_i_13
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0904_ _0308_ _0310_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0697_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0144_ VGND VGND VPWR
+ VPWR _0145_ sky130_fd_sc_hd__xnor2_1
X_0766_ manchester_baby_instance.ram_data_o_29 manchester_baby_instance.ram_data_i_29
+ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__and2b_1
X_0835_ manchester_baby_instance.ram_data_o_13 manchester_baby_instance.ram_data_i_13
+ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1318_ manchester_baby_instance.BASE_0.s_tickNext net67 VGND VGND VPWR VPWR _0101_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1249_ _0640_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1034_ _0459_ manchester_baby_instance.ram_data_o_24 _0414_ VGND VGND VPWR VPWR _0460_
+ sky130_fd_sc_hd__mux2_1
X_1103_ _0271_ _0519_ _0269_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_26_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0749_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_10_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0818_ manchester_baby_instance.ram_data_o_9 manchester_baby_instance.ram_data_i_9
+ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _0445_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1497_ manchester_baby_instance.ram_data_o_31 net12 VGND VGND VPWR VPWR ram_data_io[31]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout13 net15 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_0_32_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1351_ net77 _0626_ net59 manchester_baby_instance.BASE_0.s_countReg\[25\] VGND VGND
+ VPWR VPWR _0674_ sky130_fd_sc_hd__or4b_4
X_1420_ clknet_3_2__leaf_clock _0106_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_1282_ _0643_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0997_ manchester_baby_instance.ram_data_i_29 _0406_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0920_ _0350_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0851_ _0248_ _0252_ _0281_ _0282_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__o311a_1
X_0782_ manchester_baby_instance.ram_data_o_6 manchester_baby_instance.ram_data_i_6
+ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__xnor2_1
X_1334_ manchester_baby_instance.BASE_0.s_countReg\[16\] _0622_ VGND VGND VPWR VPWR
+ _0665_ sky130_fd_sc_hd__nor2_1
X_1403_ manchester_baby_instance.CIRCUIT_0.GATES_13.result _0090_ VGND VGND VPWR VPWR
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1265_ _0641_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
X_1196_ _0386_ _0597_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _0416_ _0464_ _0472_ _0473_ _0421_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_31_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0834_ manchester_baby_instance.ram_data_i_14 manchester_baby_instance.ram_data_o_14
+ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0903_ _0280_ _0290_ _0313_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0696_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ _0143_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a21o_1
X_0765_ _0198_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1317_ manchester_baby_instance.BASE_0.s_countReg\[8\] _0654_ VGND VGND VPWR VPWR
+ _0656_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1248_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _0583_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1102_ _0278_ _0518_ _0286_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1033_ _0416_ _0450_ _0457_ _0458_ _0421_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__a32o_1
XFILLER_0_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0817_ _0247_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0679_ _0125_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nor2_1
X_0748_ manchester_baby_instance.CIRCUIT_0.Acc.tick _0089_ _0187_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1016_ _0444_ manchester_baby_instance.ram_data_o_27 _0414_ VGND VGND VPWR VPWR _0445_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1496_ manchester_baby_instance.ram_data_o_30 net12 VGND VGND VPWR VPWR ram_data_io[30]
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout14 net15 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XFILLER_0_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1350_ _0673_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_1281_ _0639_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0996_ _0425_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1479_ manchester_baby_instance.ram_data_o_13 net12 VGND VGND VPWR VPWR ram_data_io[13]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0850_ _0246_ _0247_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__or2_1
X_1402_ manchester_baby_instance.CIRCUIT_0.GATES_13.result _0089_ VGND VGND VPWR VPWR
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0781_ manchester_baby_instance.ram_data_o_5 manchester_baby_instance.ram_data_i_5
+ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and2b_1
X_1333_ _0622_ net35 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__nand2_1
X_1264_ _0641_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
X_1195_ _0392_ _0599_ _0421_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0979_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_34_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0902_ _0323_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ _0264_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0695_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] manchester_baby_instance.ram_data_i_3
+ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__o21a_1
X_0764_ net70 manchester_baby_instance.ram_data_i_0 _0190_ VGND VGND VPWR VPWR _0198_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1316_ _0654_ _0655_ _0630_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__o21a_1
X_1247_ net1 VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__buf_4
X_1178_ _0584_ _0243_ _0222_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1032_ manchester_baby_instance.ram_data_i_24 _0402_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__xnor2_1
X_1101_ _0517_ _0284_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0747_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR
+ VPWR _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0816_ manchester_baby_instance.ram_data_i_10 manchester_baby_instance.ram_data_o_10
+ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0678_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ _0440_ _0441_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_64_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_1__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1495_ manchester_baby_instance.ram_data_o_29 net14 VGND VGND VPWR VPWR ram_data_io[29]
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_52_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout15 net16 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _0642_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0995_ _0210_ _0377_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1478_ manchester_baby_instance.ram_data_o_12 net10 VGND VGND VPWR VPWR ram_data_io[12]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ _0211_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1401_ clknet_3_6__leaf_clock _0088_ _0041_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1332_ manchester_baby_instance.BASE_0.s_countReg\[14\] _0662_ net34 VGND VGND VPWR
+ VPWR _0664_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1194_ manchester_baby_instance.ram_data_i_3 _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__nor2_1
X_1263_ _0641_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0978_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] _0188_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__and3b_1
XFILLER_0_6_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0763_ _0197_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0832_ manchester_baby_instance.ram_data_o_14 manchester_baby_instance.ram_data_i_14
+ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__and2b_1
X_0901_ _0328_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0694_ _0133_ _0140_ _0141_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__o21ai_1
X_1315_ manchester_baby_instance.BASE_0.s_countReg\[7\] _0618_ VGND VGND VPWR VPWR
+ _0655_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1246_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0637_ _0638_ manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1177_ _0231_ _0242_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1031_ _0437_ _0358_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _0228_ _0245_ _0263_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_44_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0746_ manchester_baby_instance.CIRCUIT_0.Acc.tick manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ _0126_ _0188_ net60 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__a41o_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0815_ _0246_ _0247_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0677_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1229_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__buf_6
XFILLER_0_62_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ _0404_ _0442_ _0421_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_14_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0729_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0131_ _0174_ _0130_
+ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1494_ manchester_baby_instance.ram_data_o_28 net14 VGND VGND VPWR VPWR ram_data_io[28]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout16 net7 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0207_ _0378_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1477_ manchester_baby_instance.ram_data_o_11 net10 VGND VGND VPWR VPWR ram_data_io[11]
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1400_ clknet_3_3__leaf_clock _0087_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_derivedClock
+ sky130_fd_sc_hd__dfxtp_1
X_1331_ manchester_baby_instance.BASE_0.s_countReg\[14\] _0662_ VGND VGND VPWR VPWR
+ _0107_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1193_ _0132_ _0134_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR VPWR _0598_
+ sky130_fd_sc_hd__and3_1
X_1262_ _0641_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ _0384_ _0387_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0330_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0693_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0132_ VGND VGND VPWR
+ VPWR _0141_ sky130_fd_sc_hd__nand2_1
X_0762_ net71 _0134_ _0190_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0831_ manchester_baby_instance.ram_data_i_15 manchester_baby_instance.ram_data_o_15
+ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1314_ manchester_baby_instance.BASE_0.s_countReg\[7\] _0618_ VGND VGND VPWR VPWR
+ _0654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1245_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0637_ _0638_ manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__a22o_1
X_1176_ _0219_ _0223_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _0456_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ manchester_baby_instance.ram_data_o_10 manchester_baby_instance.ram_data_i_10
+ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0676_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR VPWR
+ _0124_ sky130_fd_sc_hd__and3b_1
X_0745_ _0187_ _0128_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1228_ manchester_baby_instance.BASE_0.s_countReg\[25\] _0628_ VGND VGND VPWR VPWR
+ _0629_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1159_ _0568_ manchester_baby_instance.ram_data_o_8 _0538_ VGND VGND VPWR VPWR _0569_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1013_ manchester_baby_instance.ram_data_i_26 _0403_ manchester_baby_instance.ram_data_i_27
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ _0132_ _0158_ _0168_ _0156_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1493_ manchester_baby_instance.ram_data_o_27 net14 VGND VGND VPWR VPWR ram_data_io[27]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0412_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_14_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1476_ manchester_baby_instance.ram_data_o_10 net10 VGND VGND VPWR VPWR ram_data_io[10]
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_37_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1330_ _0662_ net48 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__nand2_1
X_1261_ _0641_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
X_1192_ _0595_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__xnor2_1
X_0976_ _0389_ _0407_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1459_ ram_data_io[25] net15 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_25
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_25_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0830_ _0248_ _0252_ _0257_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or4b_1
X_0692_ _0135_ _0139_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__and2_1
X_0761_ _0196_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1244_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0637_ _0638_ manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__a22o_1
X_1313_ _0618_ net27 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1175_ _0582_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_0959_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0813_ manchester_baby_instance.ram_data_o_11 manchester_baby_instance.ram_data_i_11
+ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR
+ VPWR _0187_ sky130_fd_sc_hd__inv_2
X_1227_ _0616_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__nand2_2
X_1158_ _0484_ _0566_ _0567_ _0424_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1089_ _0328_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_50_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1012_ _0364_ _0367_ _0439_ _0386_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0727_ _0148_ _0171_ _0172_ _0154_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1492_ manchester_baby_instance.ram_data_o_26 net14 VGND VGND VPWR VPWR ram_data_io[26]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0992_ _0423_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1475_ manchester_baby_instance.ram_data_o_9 net9 VGND VGND VPWR VPWR ram_data_io[9]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1191_ _0231_ _0239_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nor2_1
X_1260_ _0641_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0975_ manchester_baby_instance.ram_data_i_29 manchester_baby_instance.ram_data_i_30
+ _0406_ _0390_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1458_ ram_data_io[24] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_24
+ sky130_fd_sc_hd__dlxtn_1
X_1389_ clknet_3_5__leaf_clock _0076_ _0030_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_29
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0760_ net73 _0132_ _0190_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0691_ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1243_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0637_ _0638_ manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
+ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__a22o_1
X_1312_ manchester_baby_instance.BASE_0.s_countReg\[5\] _0651_ manchester_baby_instance.BASE_0.s_countReg\[6\]
+ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__o21ai_1
X_1174_ _0581_ manchester_baby_instance.ram_data_o_6 _0538_ VGND VGND VPWR VPWR _0582_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0958_ manchester_baby_instance.ram_data_i_3 manchester_baby_instance.ram_data_i_2
+ manchester_baby_instance.ram_data_i_1 manchester_baby_instance.ram_data_i_0 VGND
+ VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_30_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0889_ _0320_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__nand2_1
Xclkbuf_3_4__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_4__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0743_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] _0131_ _0186_ _0130_
+ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0812_ _0229_ _0231_ _0242_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1226_ net76 _0626_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nor2_4
X_1157_ _0544_ _0262_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1088_ _0506_ _0333_ _0341_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_58_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1011_ _0367_ _0439_ _0364_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0726_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0153_ VGND VGND VPWR
+ VPWR _0172_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1209_ _0412_ _0609_ _0610_ _0611_ _0429_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1491_ manchester_baby_instance.ram_data_o_25 net15 VGND VGND VPWR VPWR ram_data_io[25]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0152_ _0154_ _0156_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__o31a_1
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0991_ _0422_ manchester_baby_instance.ram_data_o_30 _0414_ VGND VGND VPWR VPWR _0423_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1474_ manchester_baby_instance.ram_data_o_8 net9 VGND VGND VPWR VPWR ram_data_io[8]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1190_ _0235_ _0237_ _0241_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ manchester_baby_instance.ram_data_i_29 manchester_baby_instance.ram_data_i_30
+ _0390_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__and4_1
X_1457_ ram_data_io[23] net14 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_23
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1388_ clknet_3_7__leaf_clock _0075_ _0029_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_28
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0690_ _0136_ _0137_ _0135_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1311_ manchester_baby_instance.BASE_0.s_countReg\[5\] _0651_ VGND VGND VPWR VPWR
+ _0098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1242_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] _0637_ _0638_ manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
+ VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0484_ _0579_ _0580_ _0424_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0957_ manchester_baby_instance.ram_data_i_31 VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0888_ _0318_ _0319_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0742_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] _0182_ _0185_ VGND
+ VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a21o_1
X_0811_ _0219_ _0223_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1225_ _0625_ manchester_baby_instance.BASE_0.s_countReg\[22\] VGND VGND VPWR VPWR
+ _0626_ sky130_fd_sc_hd__or2_4
X_1156_ manchester_baby_instance.ram_data_i_8 _0395_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__xnor2_1
X_1087_ _0280_ _0290_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _0438_ _0372_ _0369_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_6_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0725_ _0140_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__xor2_1
X_1208_ _0134_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1139_ _0416_ _0548_ _0551_ _0429_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1490_ manchester_baby_instance.ram_data_o_24 net15 VGND VGND VPWR VPWR ram_data_io[24]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0708_ _0155_ _0129_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ _0416_ _0381_ _0418_ _0420_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1473_ manchester_baby_instance.ram_data_o_7 net9 VGND VGND VPWR VPWR ram_data_io[7]
+ sky130_fd_sc_hd__dlxtp_1
XPHY_EDGE_ROW_59_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0973_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1387_ clknet_3_7__leaf_clock _0074_ _0028_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_27
+ sky130_fd_sc_hd__dfrtp_1
X_1456_ ram_data_io[22] net15 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_22
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_10_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1241_ _0125_ _0188_ _0632_ _0127_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a22o_1
X_1310_ _0651_ net43 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0216_ _0570_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0956_ _0388_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0887_ _0318_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or2_1
X_1439_ ram_data_io[5] net9 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_5
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_18_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0810_ _0220_ _0221_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__xor2_2
X_0741_ _0183_ _0159_ _0184_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR
+ VPWR _0185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1224_ manchester_baby_instance.BASE_0.s_countReg\[20\] net21 _0624_ VGND VGND VPWR
+ VPWR _0625_ sky130_fd_sc_hd__or3_4
X_1155_ _0565_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
X_1086_ _0505_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0939_ _0350_ _0356_ _0351_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0724_ _0141_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1207_ _0232_ manchester_baby_instance.ram_data_o_0 _0233_ _0234_ VGND VGND VPWR
+ VPWR _0610_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1138_ manchester_baby_instance.ram_data_i_11 _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__xor2_1
X_1069_ _0490_ manchester_baby_instance.ram_data_o_20 _0470_ VGND VGND VPWR VPWR _0491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 manchester_baby_instance.BASE_1.s_bufferRegs\[0\] VGND VGND VPWR VPWR net18
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0707_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
+ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] VGND VGND VPWR VPWR _0155_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ manchester_baby_instance.ram_data_o_6 net9 VGND VGND VPWR VPWR ram_data_io[6]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0972_ manchester_baby_instance.ram_data_i_28 _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1386_ clknet_3_7__leaf_clock _0073_ _0027_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_26
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1455_ ram_data_io[21] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_21
+ sky130_fd_sc_hd__dlxtn_1
XTAP_TAPCELL_ROW_25_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1240_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__dlymetal6s2s_1
X_1171_ manchester_baby_instance.ram_data_i_6 _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0955_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ _0188_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] VGND VGND VPWR VPWR _0388_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0886_ manchester_baby_instance.ram_data_o_17 manchester_baby_instance.ram_data_i_17
+ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1438_ ram_data_io[4] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_4
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1369_ clknet_3_1__leaf_clock _0056_ _0010_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_9
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_90 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0740_ _0148_ _0136_ _0158_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a21o_1
X_1223_ manchester_baby_instance.BASE_0.s_countReg\[18\] net38 _0622_ _0623_ VGND
+ VGND VPWR VPWR _0624_ sky130_fd_sc_hd__or4_4
X_1154_ _0564_ manchester_baby_instance.ram_data_o_9 _0538_ VGND VGND VPWR VPWR _0565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1085_ _0504_ manchester_baby_instance.ram_data_o_18 _0470_ VGND VGND VPWR VPWR _0505_
+ sky130_fd_sc_hd__mux2_1
X_0938_ _0336_ _0340_ _0345_ _0359_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__a311o_1
X_0869_ _0296_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0723_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0132_ VGND VGND VPWR
+ VPWR _0169_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1206_ _0235_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__inv_2
X_1137_ manchester_baby_instance.ram_data_i_10 _0549_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ _0416_ _0476_ _0488_ _0489_ _0429_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 manchester_baby_instance.BASE_1.s_derivedClock VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0706_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0153_ _0150_ VGND
+ VGND VPWR VPWR _0154_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_40_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ manchester_baby_instance.ram_data_o_5 net9 VGND VGND VPWR VPWR ram_data_io[5]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_7__leaf_clock sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_28_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0971_ manchester_baby_instance.ram_data_i_26 manchester_baby_instance.ram_data_i_27
+ _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1454_ ram_data_io[20] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_20
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ clknet_3_7__leaf_clock _0072_ _0026_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_25
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0392_ _0393_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0954_ _0203_ _0381_ _0383_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ manchester_baby_instance.ram_data_o_18 manchester_baby_instance.ram_data_i_18
+ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1437_ ram_data_io[3] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_3
+ sky130_fd_sc_hd__dlxtn_2
XFILLER_0_2_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1299_ net63 net55 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__and2b_1
X_1368_ clknet_3_0__leaf_clock _0055_ _0009_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_8
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1222_ manchester_baby_instance.BASE_0.s_countReg\[16\] manchester_baby_instance.BASE_0.s_countReg\[17\]
+ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or2_1
X_1153_ _0416_ _0561_ _0563_ _0429_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__a22o_1
X_1084_ _0412_ _0493_ _0500_ _0503_ _0429_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0937_ _0364_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0799_ manchester_baby_instance.ram_data_i_0 VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0868_ _0299_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0722_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] VGND VGND VPWR VPWR _0168_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1205_ _0608_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1136_ manchester_baby_instance.ram_data_i_8 manchester_baby_instance.ram_data_i_9
+ _0395_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__and3_1
X_1067_ manchester_baby_instance.ram_data_i_20 _0482_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 manchester_baby_instance.BASE_0.s_countReg\[0\] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0705_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ manchester_baby_instance.ram_data_o_31 VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _0274_ _0531_ _0532_ _0386_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1470_ manchester_baby_instance.ram_data_o_4 net11 VGND VGND VPWR VPWR ram_data_io[4]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ manchester_baby_instance.ram_data_i_24 manchester_baby_instance.ram_data_i_25
+ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__and3_1
X_1453_ ram_data_io[19] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_19
+ sky130_fd_sc_hd__dlxtn_1
X_1384_ clknet_3_5__leaf_clock _0071_ _0025_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_24
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0953_ _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0884_ _0310_ _0314_ _0315_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ ram_data_io[2] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_2
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_2_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1367_ clknet_3_0__leaf_clock _0054_ _0008_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_7
+ sky130_fd_sc_hd__dfrtp_2
X_1298_ _0646_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__buf_6
XFILLER_0_32_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1152_ _0549_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or2_1
X_1083_ manchester_baby_instance.ram_data_i_18 _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0936_ _0367_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0798_ manchester_baby_instance.ram_data_o_2 _0221_ _0230_ _0132_ VGND VGND VPWR
+ VPWR _0231_ sky130_fd_sc_hd__and4b_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0867_ _0297_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1419_ clknet_3_2__leaf_clock _0105_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0721_ _0130_ _0166_ _0167_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1204_ _0607_ manchester_baby_instance.ram_data_o_2 _0413_ VGND VGND VPWR VPWR _0608_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1135_ _0248_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__xor2_1
X_1066_ _0311_ _0462_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0919_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 manchester_baby_instance.BASE_0.s_countReg\[21\] VGND VGND VPWR VPWR net21
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0704_ _0129_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1049_ manchester_baby_instance.ram_data_i_22 _0401_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__xnor2_1
X_1118_ _0531_ _0532_ _0274_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1383_ clknet_3_5__leaf_clock _0070_ _0024_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_23
+ sky130_fd_sc_hd__dfrtp_1
X_1452_ ram_data_io[18] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_18
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0952_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] _0187_ _0128_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or4b_1
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1504_ clknet_3_3__leaf_clock _0123_ _0046_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0883_ _0310_ _0314_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__and3_1
X_1435_ ram_data_io[1] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_1
+ sky130_fd_sc_hd__dlxtn_1
X_1366_ clknet_3_0__leaf_clock _0053_ _0007_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_6
+ sky130_fd_sc_hd__dfrtp_1
X_1297_ _0129_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1220_ manchester_baby_instance.BASE_0.s_countReg\[13\] manchester_baby_instance.BASE_0.s_countReg\[14\]
+ manchester_baby_instance.BASE_0.s_countReg\[15\] _0620_ VGND VGND VPWR VPWR _0621_
+ sky130_fd_sc_hd__or4_4
X_1151_ manchester_baby_instance.ram_data_i_8 _0395_ manchester_baby_instance.ram_data_i_9
+ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1082_ manchester_baby_instance.ram_data_i_17 _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0935_ _0365_ _0347_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0866_ _0297_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__or2_1
X_0797_ manchester_baby_instance.ram_data_i_3 manchester_baby_instance.ram_data_o_3
+ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1349_ _0627_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or2_1
X_1418_ clknet_3_2__leaf_clock _0104_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0720_ _0131_ _0154_ _0156_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1203_ _0412_ _0603_ _0604_ _0606_ _0429_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__a32o_1
X_1134_ _0250_ _0251_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _0487_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0918_ _0346_ manchester_baby_instance.ram_data_i_24 _0349_ VGND VGND VPWR VPWR _0351_
+ sky130_fd_sc_hd__and3_1
X_0849_ _0246_ _0247_ _0250_ _0251_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold6 _0670_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0703_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] VGND VGND VPWR VPWR
+ _0151_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ _0517_ _0284_ _0277_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_332 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ _0301_ _0339_ _0463_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand3_1
XFILLER_0_43_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1382_ clknet_3_5__leaf_clock _0069_ _0023_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_22
+ sky130_fd_sc_hd__dfrtp_1
X_1451_ ram_data_io[17] net13 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_17
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0951_ _0203_ _0381_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_30_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ manchester_baby_instance.ram_data_o_18 manchester_baby_instance.ram_data_i_18
+ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__and2b_1
X_1503_ clknet_3_3__leaf_clock _0122_ _0045_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1296_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] _0128_ VGND VGND
+ VPWR VPWR _0645_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1434_ ram_data_io[0] net11 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_0
+ sky130_fd_sc_hd__dlxtn_2
X_1365_ clknet_3_0__leaf_clock _0052_ _0006_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_5
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_0__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1150_ _0257_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1081_ manchester_baby_instance.ram_data_i_16 _0399_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0934_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ manchester_baby_instance.ram_data_o_21 manchester_baby_instance.ram_data_i_21
+ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and2b_1
X_1417_ clknet_3_2__leaf_clock _0103_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ _0213_ _0216_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__or2_1
X_1348_ manchester_baby_instance.BASE_0.s_countReg\[23\] _0626_ VGND VGND VPWR VPWR
+ _0672_ sky130_fd_sc_hd__and2_1
X_1279_ _0642_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1202_ _0598_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or2_1
X_1133_ _0281_ _0545_ _0252_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1064_ _0486_ manchester_baby_instance.ram_data_o_21 _0470_ VGND VGND VPWR VPWR _0487_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0917_ _0346_ manchester_baby_instance.ram_data_i_24 _0349_ VGND VGND VPWR VPWR _0350_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0848_ _0255_ _0261_ _0256_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a21bo_1
X_0779_ manchester_baby_instance.ram_data_o_7 manchester_baby_instance.ram_data_i_7
+ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0702_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0124_ _0126_ VGND VGND VPWR
+ VPWR _0150_ sky130_fd_sc_hd__and3b_1
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1047_ _0471_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ _0275_ _0276_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450_ ram_data_io[16] net10 VGND VGND VPWR VPWR manchester_baby_instance.ram_data_i_16
+ sky130_fd_sc_hd__dlxtn_1
XFILLER_0_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1381_ clknet_3_5__leaf_clock _0068_ _0022_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_21
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ _0200_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0881_ manchester_baby_instance.ram_data_o_19 _0309_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1502_ clknet_3_3__leaf_clock _0121_ _0044_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_1433_ clknet_3_3__leaf_clock manchester_baby_instance.BASE_0.s_tickNext VGND VGND
+ VPWR VPWR manchester_baby_instance.BASE_0.s_tickReg sky130_fd_sc_hd__dfxtp_1
X_1295_ _0128_ _0631_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1364_ clknet_3_0__leaf_clock _0051_ _0005_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_4
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ _0322_ _0342_ _0492_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__nand3_1
XFILLER_0_59_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0933_ _0365_ _0347_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nor2_1
X_0864_ manchester_baby_instance.ram_data_o_22 manchester_baby_instance.ram_data_i_22
+ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0795_ _0213_ _0216_ _0224_ _0226_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__o311a_1
XFILLER_0_23_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1347_ _0626_ _0671_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1416_ clknet_3_1__leaf_clock _0102_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0642_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1201_ _0134_ manchester_baby_instance.ram_data_i_0 _0132_ VGND VGND VPWR VPWR _0605_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1132_ _0257_ _0262_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1063_ _0424_ _0478_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_63_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0916_ _0347_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ manchester_baby_instance.ram_data_o_6 manchester_baby_instance.ram_data_i_6
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__and2b_1
X_0847_ _0228_ _0245_ _0263_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_342 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 _0650_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0701_ _0146_ _0147_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1046_ _0469_ manchester_baby_instance.ram_data_o_23 _0470_ VGND VGND VPWR VPWR _0471_
+ sky130_fd_sc_hd__mux2_1
X_1115_ _0530_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1029_ _0455_ manchester_baby_instance.ram_data_o_25 _0414_ VGND VGND VPWR VPWR _0456_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ clknet_3_5__leaf_clock _0067_ _0021_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_20
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ _0302_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or2b_1
X_1501_ clknet_3_3__leaf_clock _0120_ _0043_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_1432_ clknet_3_2__leaf_clock _0118_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_1363_ clknet_3_0__leaf_clock _0050_ _0004_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_3
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1294_ _0639_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_43_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ manchester_baby_instance.ram_data_o_26 manchester_baby_instance.ram_data_i_26
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0863_ _0294_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ _0211_ _0212_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or2_1
X_1346_ manchester_baby_instance.BASE_0.s_countReg\[22\] _0625_ VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1415_ clknet_3_1__leaf_clock _0101_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_1277_ _0642_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1200_ _0235_ _0237_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1131_ _0228_ _0245_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_1
X_1062_ _0401_ _0483_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__o21a_1
X_0915_ manchester_baby_instance.ram_data_i_25 manchester_baby_instance.ram_data_o_25
+ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0777_ _0208_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0846_ _0266_ _0271_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1329_ manchester_baby_instance.BASE_0.s_countReg\[13\] _0620_ VGND VGND VPWR VPWR
+ _0663_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 _0096_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0700_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0124_ _0125_ VGND VGND VPWR
+ VPWR _0148_ sky130_fd_sc_hd__and3_2
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1114_ _0529_ manchester_baby_instance.ram_data_o_14 _0470_ VGND VGND VPWR VPWR _0530_
+ sky130_fd_sc_hd__mux2_1
X_1045_ _0413_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0829_ manchester_baby_instance.ram_data_o_7 _0259_ _0261_ VGND VGND VPWR VPWR _0262_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1028_ _0451_ _0452_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_230 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1500_ clknet_3_6__leaf_clock _0119_ _0042_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1293_ net19 net56 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__xnor2_1
X_1431_ clknet_3_3__leaf_clock _0117_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_1362_ clknet_3_1__leaf_clock _0049_ _0003_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_2
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0931_ _0362_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__or2_1
X_0862_ _0292_ _0293_ _0291_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a21o_1
Xrebuffer1 manchester_baby_instance.BASE_0.s_countReg\[0\] VGND VGND VPWR VPWR net17
+ sky130_fd_sc_hd__dlygate4sd1_1
X_0793_ _0211_ _0212_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_21_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1345_ _0625_ net22 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__nand2_1
X_1276_ _0642_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
X_1414_ clknet_3_2__leaf_clock _0100_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1130_ _0543_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_1061_ _0388_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ manchester_baby_instance.ram_data_o_25 manchester_baby_instance.ram_data_i_25
+ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0845_ _0274_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0776_ manchester_baby_instance.ram_data_o_27 manchester_baby_instance.ram_data_i_27
+ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1328_ manchester_baby_instance.BASE_0.s_countReg\[13\] _0620_ VGND VGND VPWR VPWR
+ _0662_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ _0639_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_3_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1044_ _0465_ _0466_ _0468_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__o21ai_1
X_1113_ _0484_ _0527_ _0528_ _0424_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0759_ _0195_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_0828_ _0260_ manchester_baby_instance.ram_data_i_7 _0258_ VGND VGND VPWR VPWR _0261_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ _0403_ _0453_ _0421_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_3__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_3__leaf_clock sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_10_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1430_ clknet_3_3__leaf_clock _0116_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_1292_ net55 manchester_baby_instance.BASE_0.s_tickReg VGND VGND VPWR VPWR _0644_
+ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_38_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1361_ clknet_3_6__leaf_clock _0048_ _0002_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0930_ manchester_baby_instance.ram_data_o_26 manchester_baby_instance.ram_data_i_26
+ _0209_ _0360_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and4b_1
X_0861_ _0291_ _0292_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ _0214_ _0215_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or2_1
X_1413_ clknet_3_1__leaf_clock net28 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1344_ manchester_baby_instance.BASE_0.s_countReg\[20\] _0624_ net21 VGND VGND VPWR
+ VPWR _0670_ sky130_fd_sc_hd__o21ai_1
X_1275_ _0642_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ manchester_baby_instance.ram_data_i_20 _0482_ manchester_baby_instance.ram_data_i_21
+ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0775_ manchester_baby_instance.ram_data_o_28 manchester_baby_instance.ram_data_i_28
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__xor2_1
X_0913_ manchester_baby_instance.ram_data_o_24 VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0844_ _0275_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_54_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1327_ _0620_ net30 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1189_ _0594_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
X_1258_ _0640_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1043_ _0402_ _0467_ _0421_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o21ai_1
X_1112_ _0271_ _0519_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0758_ net75 manchester_baby_instance.ram_data_i_3 _0190_ VGND VGND VPWR VPWR _0195_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ manchester_baby_instance.ram_data_o_7 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0689_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0134_ VGND VGND VPWR
+ VPWR _0137_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1026_ manchester_baby_instance.ram_data_i_24 _0402_ manchester_baby_instance.ram_data_i_25
+ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1009_ _0437_ _0359_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput2 net2 VGND VGND VPWR VPWR ram_addr_o[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1360_ clknet_3_4__leaf_clock _0047_ _0001_ VGND VGND VPWR VPWR manchester_baby_instance.ram_data_o_0
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1291_ _0643_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1489_ manchester_baby_instance.ram_data_o_23 net15 VGND VGND VPWR VPWR ram_data_io[23]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ manchester_baby_instance.ram_data_i_23 manchester_baby_instance.ram_data_o_23
+ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__or2b_1
X_0791_ _0219_ _0222_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a21bo_1
X_1343_ manchester_baby_instance.BASE_0.s_countReg\[20\] _0624_ VGND VGND VPWR VPWR
+ _0113_ sky130_fd_sc_hd__xnor2_1
X_1412_ clknet_3_1__leaf_clock net54 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1274_ _0642_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0388_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_57_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0912_ _0313_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0774_ manchester_baby_instance.ram_data_o_28 _0204_ _0206_ VGND VGND VPWR VPWR _0207_
+ sky130_fd_sc_hd__o21a_1
X_0843_ manchester_baby_instance.ram_data_o_11 manchester_baby_instance.ram_data_i_11
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nand2b_1
X_1326_ manchester_baby_instance.BASE_0.s_countReg\[10\] manchester_baby_instance.BASE_0.s_countReg\[11\]
+ _0619_ net29 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_54_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ _0593_ manchester_baby_instance.ram_data_o_4 _0538_ VGND VGND VPWR VPWR _0594_
+ sky130_fd_sc_hd__mux2_1
X_1257_ _0640_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1042_ manchester_baby_instance.ram_data_i_22 _0401_ manchester_baby_instance.ram_data_i_23
+ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a21oi_1
X_1111_ manchester_baby_instance.ram_data_i_14 _0522_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0688_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] manchester_baby_instance.ram_data_i_0
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__nand2_1
X_0757_ _0194_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
X_0826_ manchester_baby_instance.ram_data_i_7 _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1309_ net42 _0617_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1025_ _0353_ _0356_ _0450_ _0386_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__a31o_1
X_0809_ _0235_ _0237_ _0239_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1008_ _0336_ _0340_ _0345_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput3 net3 VGND VGND VPWR VPWR ram_addr_o[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1290_ _0643_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_78 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1488_ manchester_baby_instance.ram_data_o_22 net15 VGND VGND VPWR VPWR ram_data_io[22]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0790_ _0217_ manchester_baby_instance.ram_data_o_4 _0218_ VGND VGND VPWR VPWR _0223_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1342_ _0624_ net39 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nand2_1
X_1411_ clknet_3_0__leaf_clock _0097_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_1273_ _0642_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ manchester_baby_instance.ram_data_i_30 _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0911_ _0316_ _0320_ _0323_ _0342_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o221a_1
X_0842_ manchester_baby_instance.ram_data_o_12 manchester_baby_instance.ram_data_i_12
+ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ _0199_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1325_ manchester_baby_instance.BASE_0.s_tickNext net65 VGND VGND VPWR VPWR _0104_
+ sky130_fd_sc_hd__nor2_1
X_1256_ _0640_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1187_ _0416_ _0591_ _0592_ _0484_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1110_ _0526_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1041_ _0296_ _0299_ _0464_ _0386_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ manchester_baby_instance.ram_data_o_8 manchester_baby_instance.ram_data_i_8
+ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0687_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0134_ VGND VGND VPWR
+ VPWR _0135_ sky130_fd_sc_hd__nand2_1
X_0756_ net72 manchester_baby_instance.ram_data_i_4 _0190_ VGND VGND VPWR VPWR _0194_
+ sky130_fd_sc_hd__mux2_1
X_1239_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ _0187_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1308_ manchester_baby_instance.BASE_0.s_countReg\[4\] _0617_ VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1024_ _0356_ _0450_ _0353_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0808_ _0240_ manchester_baby_instance.ram_data_o_1 _0236_ VGND VGND VPWR VPWR _0241_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_12_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0739_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] VGND VGND VPWR VPWR
+ _0183_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold60 manchester_baby_instance.BASE_0.s_countReg\[23\] VGND VGND VPWR VPWR net76
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1007_ _0436_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput4 net4 VGND VGND VPWR VPWR ram_addr_o[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1487_ manchester_baby_instance.ram_data_o_21 net13 VGND VGND VPWR VPWR ram_data_io[21]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1410_ clknet_3_0__leaf_clock net25 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1341_ manchester_baby_instance.BASE_0.s_countReg\[18\] _0622_ _0623_ net38 VGND
+ VGND VPWR VPWR _0669_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1272_ _0642_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ manchester_baby_instance.ram_data_i_29 _0406_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0772_ manchester_baby_instance.ram_data_i_29 manchester_baby_instance.ram_data_o_29
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ _0317_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__inv_2
X_0841_ _0272_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1324_ manchester_baby_instance.BASE_0.s_countReg\[11\] _0658_ VGND VGND VPWR VPWR
+ _0660_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ manchester_baby_instance.ram_data_i_4 _0392_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__xnor2_1
X_1255_ _0640_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_6__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_3_6__leaf_clock sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_36_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ _0299_ _0464_ _0296_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0755_ _0193_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0824_ _0255_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nand2_1
X_0686_ manchester_baby_instance.ram_data_i_1 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1238_ _0635_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.GATES_13.result
+ sky130_fd_sc_hd__clkbuf_1
X_1307_ _0617_ net24 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1169_ _0577_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _0437_ _0358_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0738_ _0148_ _0136_ _0150_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0807_ _0134_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold61 manchester_baby_instance.BASE_0.s_countReg\[23\] VGND VGND VPWR VPWR net77
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _0435_ manchester_baby_instance.ram_data_o_28 _0414_ VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput5 net5 VGND VGND VPWR VPWR ram_addr_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1486_ manchester_baby_instance.ram_data_o_20 net15 VGND VGND VPWR VPWR ram_data_io[20]
+ sky130_fd_sc_hd__dlxtp_1
XFILLER_0_64_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1340_ _0667_ _0668_ manchester_baby_instance.BASE_0.s_tickNext VGND VGND VPWR VPWR
+ _0111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1271_ _0642_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ _0380_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1469_ manchester_baby_instance.ram_data_o_3 net11 VGND VGND VPWR VPWR ram_data_io[3]
+ sky130_fd_sc_hd__dlxtp_1
XTAP_TAPCELL_ROW_57_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0771_ manchester_baby_instance.ram_data_i_28 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0840_ manchester_baby_instance.ram_data_o_12 manchester_baby_instance.ram_data_i_12
+ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ _0658_ _0659_ _0630_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__o21a_1
X_1185_ _0584_ _0243_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_19_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1254_ _0640_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0969_ manchester_baby_instance.ram_data_i_22 manchester_baby_instance.ram_data_i_23
+ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0685_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0132_ VGND VGND VPWR
+ VPWR _0133_ sky130_fd_sc_hd__nor2_1
X_0754_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] manchester_baby_instance.ram_data_i_13
+ _0190_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ _0253_ _0254_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1306_ manchester_baby_instance.BASE_0.s_countReg\[3\] _0648_ VGND VGND VPWR VPWR
+ _0650_ sky130_fd_sc_hd__nand2_1
X_1237_ net8 manchester_baby_instance.CIRCUIT_0.GATES_13.input1 VGND VGND VPWR VPWR
+ _0635_ sky130_fd_sc_hd__and2b_1
X_1099_ _0516_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
X_1168_ _0576_ manchester_baby_instance.ram_data_o_7 _0538_ VGND VGND VPWR VPWR _0577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_344 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1022_ _0449_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0737_ manchester_baby_instance.ram_data_o_31 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__inv_2
X_0806_ _0221_ _0230_ _0238_ manchester_baby_instance.ram_data_o_2 VGND VGND VPWR
+ VPWR _0239_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_12_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_241 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold40 _0644_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold51 _0656_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1005_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR ram_addr_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_53_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1485_ manchester_baby_instance.ram_data_o_19 net13 VGND VGND VPWR VPWR ram_data_io[19]
+ sky130_fd_sc_hd__dlxtp_1
.ends

