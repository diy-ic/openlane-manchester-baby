// This is the unpowered netlist.
module openlane_manchester_baby (clock,
    logisim_clock_tree_0_out,
    ram_rw_en_o,
    reset_i,
    stop_lamp_o,
    ram_addr_o,
    ram_data_io);
 input clock;
 output logisim_clock_tree_0_out;
 output ram_rw_en_o;
 input reset_i;
 output stop_lamp_o;
 output [4:0] ram_addr_o;
 inout [31:0] ram_data_io;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire \manchester_baby_instance.BASE_0.s_countReg[0] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[1] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[2] ;
 wire \manchester_baby_instance.BASE_0.s_tickNext ;
 wire \manchester_baby_instance.BASE_0.s_tickReg ;
 wire \manchester_baby_instance.BASE_1.s_bufferRegs[0] ;
 wire \manchester_baby_instance.BASE_1.s_counterValue ;
 wire \manchester_baby_instance.BASE_1.s_derivedClock ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.Acc.tick ;
 wire \manchester_baby_instance.CIRCUIT_0.GATES_13.result ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[13] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[14] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[15] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ;
 wire \manchester_baby_instance.ram_data_i_0 ;
 wire \manchester_baby_instance.ram_data_i_1 ;
 wire \manchester_baby_instance.ram_data_i_10 ;
 wire \manchester_baby_instance.ram_data_i_11 ;
 wire \manchester_baby_instance.ram_data_i_12 ;
 wire \manchester_baby_instance.ram_data_i_13 ;
 wire \manchester_baby_instance.ram_data_i_14 ;
 wire \manchester_baby_instance.ram_data_i_15 ;
 wire \manchester_baby_instance.ram_data_i_16 ;
 wire \manchester_baby_instance.ram_data_i_17 ;
 wire \manchester_baby_instance.ram_data_i_18 ;
 wire \manchester_baby_instance.ram_data_i_19 ;
 wire \manchester_baby_instance.ram_data_i_2 ;
 wire \manchester_baby_instance.ram_data_i_20 ;
 wire \manchester_baby_instance.ram_data_i_21 ;
 wire \manchester_baby_instance.ram_data_i_22 ;
 wire \manchester_baby_instance.ram_data_i_23 ;
 wire \manchester_baby_instance.ram_data_i_24 ;
 wire \manchester_baby_instance.ram_data_i_25 ;
 wire \manchester_baby_instance.ram_data_i_26 ;
 wire \manchester_baby_instance.ram_data_i_27 ;
 wire \manchester_baby_instance.ram_data_i_28 ;
 wire \manchester_baby_instance.ram_data_i_29 ;
 wire \manchester_baby_instance.ram_data_i_3 ;
 wire \manchester_baby_instance.ram_data_i_30 ;
 wire \manchester_baby_instance.ram_data_i_31 ;
 wire \manchester_baby_instance.ram_data_i_4 ;
 wire \manchester_baby_instance.ram_data_i_5 ;
 wire \manchester_baby_instance.ram_data_i_6 ;
 wire \manchester_baby_instance.ram_data_i_7 ;
 wire \manchester_baby_instance.ram_data_i_8 ;
 wire \manchester_baby_instance.ram_data_i_9 ;
 wire \manchester_baby_instance.ram_data_o_0 ;
 wire \manchester_baby_instance.ram_data_o_1 ;
 wire \manchester_baby_instance.ram_data_o_10 ;
 wire \manchester_baby_instance.ram_data_o_11 ;
 wire \manchester_baby_instance.ram_data_o_12 ;
 wire \manchester_baby_instance.ram_data_o_13 ;
 wire \manchester_baby_instance.ram_data_o_14 ;
 wire \manchester_baby_instance.ram_data_o_15 ;
 wire \manchester_baby_instance.ram_data_o_16 ;
 wire \manchester_baby_instance.ram_data_o_17 ;
 wire \manchester_baby_instance.ram_data_o_18 ;
 wire \manchester_baby_instance.ram_data_o_19 ;
 wire \manchester_baby_instance.ram_data_o_2 ;
 wire \manchester_baby_instance.ram_data_o_20 ;
 wire \manchester_baby_instance.ram_data_o_21 ;
 wire \manchester_baby_instance.ram_data_o_22 ;
 wire \manchester_baby_instance.ram_data_o_23 ;
 wire \manchester_baby_instance.ram_data_o_24 ;
 wire \manchester_baby_instance.ram_data_o_25 ;
 wire \manchester_baby_instance.ram_data_o_26 ;
 wire \manchester_baby_instance.ram_data_o_27 ;
 wire \manchester_baby_instance.ram_data_o_28 ;
 wire \manchester_baby_instance.ram_data_o_29 ;
 wire \manchester_baby_instance.ram_data_o_3 ;
 wire \manchester_baby_instance.ram_data_o_30 ;
 wire \manchester_baby_instance.ram_data_o_31 ;
 wire \manchester_baby_instance.ram_data_o_4 ;
 wire \manchester_baby_instance.ram_data_o_5 ;
 wire \manchester_baby_instance.ram_data_o_6 ;
 wire \manchester_baby_instance.ram_data_o_7 ;
 wire \manchester_baby_instance.ram_data_o_8 ;
 wire \manchester_baby_instance.ram_data_o_9 ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_159 ();
 sky130_fd_sc_hd__clkbuf_4 _0588_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0101_));
 sky130_fd_sc_hd__nor2_1 _0589_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(_0102_));
 sky130_fd_sc_hd__and2_2 _0590_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__clkbuf_4 _0591_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .X(_0104_));
 sky130_fd_sc_hd__and3b_1 _0592_ (.A_N(_0101_),
    .B(_0103_),
    .C(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_4 _0593_ (.A(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__or2b_1 _0594_ (.A(\manchester_baby_instance.ram_data_i_17 ),
    .B_N(\manchester_baby_instance.ram_data_o_17 ),
    .X(_0107_));
 sky130_fd_sc_hd__or2b_1 _0595_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B_N(\manchester_baby_instance.ram_data_o_16 ),
    .X(_0108_));
 sky130_fd_sc_hd__and2b_1 _0596_ (.A_N(\manchester_baby_instance.ram_data_i_7 ),
    .B(\manchester_baby_instance.ram_data_o_7 ),
    .X(_0109_));
 sky130_fd_sc_hd__and2b_1 _0597_ (.A_N(\manchester_baby_instance.ram_data_o_7 ),
    .B(\manchester_baby_instance.ram_data_i_7 ),
    .X(_0110_));
 sky130_fd_sc_hd__nor2_1 _0598_ (.A(_0109_),
    .B(_0110_),
    .Y(_0111_));
 sky130_fd_sc_hd__xnor2_2 _0599_ (.A(\manchester_baby_instance.ram_data_o_6 ),
    .B(\manchester_baby_instance.ram_data_i_6 ),
    .Y(_0112_));
 sky130_fd_sc_hd__and2_1 _0600_ (.A(_0111_),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__and2b_1 _0601_ (.A_N(\manchester_baby_instance.ram_data_o_5 ),
    .B(\manchester_baby_instance.ram_data_i_5 ),
    .X(_0114_));
 sky130_fd_sc_hd__or2b_1 _0602_ (.A(\manchester_baby_instance.ram_data_i_5 ),
    .B_N(\manchester_baby_instance.ram_data_o_5 ),
    .X(_0115_));
 sky130_fd_sc_hd__nor2b_2 _0603_ (.A(_0114_),
    .B_N(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\manchester_baby_instance.ram_data_o_2 ),
    .Y(_0117_));
 sky130_fd_sc_hd__buf_2 _0605_ (.A(\manchester_baby_instance.ram_data_i_2 ),
    .X(_0118_));
 sky130_fd_sc_hd__and2b_1 _0606_ (.A_N(\manchester_baby_instance.ram_data_o_3 ),
    .B(\manchester_baby_instance.ram_data_i_3 ),
    .X(_0119_));
 sky130_fd_sc_hd__or2b_1 _0607_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B_N(\manchester_baby_instance.ram_data_o_3 ),
    .X(_0120_));
 sky130_fd_sc_hd__o31a_1 _0608_ (.A1(_0117_),
    .A2(_0118_),
    .A3(_0119_),
    .B1(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__or2b_1 _0609_ (.A(_0118_),
    .B_N(\manchester_baby_instance.ram_data_o_2 ),
    .X(_0122_));
 sky130_fd_sc_hd__or2b_1 _0610_ (.A(\manchester_baby_instance.ram_data_o_2 ),
    .B_N(_0118_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_1 _0611_ (.A(_0122_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__or2b_1 _0612_ (.A(\manchester_baby_instance.ram_data_o_1 ),
    .B_N(\manchester_baby_instance.ram_data_i_1 ),
    .X(_0125_));
 sky130_fd_sc_hd__or2b_1 _0613_ (.A(\manchester_baby_instance.ram_data_o_0 ),
    .B_N(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0126_));
 sky130_fd_sc_hd__and2b_1 _0614_ (.A_N(\manchester_baby_instance.ram_data_i_1 ),
    .B(\manchester_baby_instance.ram_data_o_1 ),
    .X(_0127_));
 sky130_fd_sc_hd__a21oi_1 _0615_ (.A1(_0125_),
    .A2(_0126_),
    .B1(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__or2b_1 _0616_ (.A(\manchester_baby_instance.ram_data_o_3 ),
    .B_N(\manchester_baby_instance.ram_data_i_3 ),
    .X(_0129_));
 sky130_fd_sc_hd__nand2_1 _0617_ (.A(_0120_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__or3_1 _0618_ (.A(_0124_),
    .B(_0128_),
    .C(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__xnor2_1 _0619_ (.A(\manchester_baby_instance.ram_data_o_4 ),
    .B(\manchester_baby_instance.ram_data_i_4 ),
    .Y(_0132_));
 sky130_fd_sc_hd__a21boi_2 _0620_ (.A1(_0121_),
    .A2(_0131_),
    .B1_N(_0132_),
    .Y(_0133_));
 sky130_fd_sc_hd__or2b_1 _0621_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B_N(\manchester_baby_instance.ram_data_o_4 ),
    .X(_0134_));
 sky130_fd_sc_hd__a21oi_1 _0622_ (.A1(_0115_),
    .A2(_0134_),
    .B1(_0114_),
    .Y(_0135_));
 sky130_fd_sc_hd__or2b_1 _0623_ (.A(\manchester_baby_instance.ram_data_i_6 ),
    .B_N(\manchester_baby_instance.ram_data_o_6 ),
    .X(_0136_));
 sky130_fd_sc_hd__or2_1 _0624_ (.A(_0110_),
    .B(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__inv_2 _0625_ (.A(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__a211o_1 _0626_ (.A1(_0113_),
    .A2(_0135_),
    .B1(_0138_),
    .C1(_0109_),
    .X(_0139_));
 sky130_fd_sc_hd__a31oi_4 _0627_ (.A1(_0113_),
    .A2(_0116_),
    .A3(_0133_),
    .B1(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__xnor2_1 _0628_ (.A(\manchester_baby_instance.ram_data_o_15 ),
    .B(\manchester_baby_instance.ram_data_i_15 ),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _0629_ (.A(\manchester_baby_instance.ram_data_o_14 ),
    .B(\manchester_baby_instance.ram_data_i_14 ),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _0630_ (.A(_0141_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__xnor2_2 _0631_ (.A(\manchester_baby_instance.ram_data_o_12 ),
    .B(\manchester_baby_instance.ram_data_i_12 ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _0632_ (.A(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__and2b_1 _0633_ (.A_N(\manchester_baby_instance.ram_data_o_13 ),
    .B(\manchester_baby_instance.ram_data_i_13 ),
    .X(_0146_));
 sky130_fd_sc_hd__or2b_1 _0634_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B_N(\manchester_baby_instance.ram_data_o_13 ),
    .X(_0147_));
 sky130_fd_sc_hd__or2b_1 _0635_ (.A(_0146_),
    .B_N(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__or3_1 _0636_ (.A(_0143_),
    .B(_0145_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__xnor2_1 _0637_ (.A(\manchester_baby_instance.ram_data_o_11 ),
    .B(\manchester_baby_instance.ram_data_i_11 ),
    .Y(_0150_));
 sky130_fd_sc_hd__xnor2_1 _0638_ (.A(\manchester_baby_instance.ram_data_o_10 ),
    .B(\manchester_baby_instance.ram_data_i_10 ),
    .Y(_0151_));
 sky130_fd_sc_hd__and2_1 _0639_ (.A(_0150_),
    .B(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__or2b_1 _0640_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B_N(\manchester_baby_instance.ram_data_o_8 ),
    .X(_0153_));
 sky130_fd_sc_hd__or2b_1 _0641_ (.A(\manchester_baby_instance.ram_data_o_8 ),
    .B_N(\manchester_baby_instance.ram_data_i_8 ),
    .X(_0154_));
 sky130_fd_sc_hd__nand2_1 _0642_ (.A(_0153_),
    .B(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__or2b_1 _0643_ (.A(\manchester_baby_instance.ram_data_i_9 ),
    .B_N(\manchester_baby_instance.ram_data_o_9 ),
    .X(_0156_));
 sky130_fd_sc_hd__or2b_1 _0644_ (.A(\manchester_baby_instance.ram_data_o_9 ),
    .B_N(\manchester_baby_instance.ram_data_i_9 ),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _0645_ (.A(_0156_),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2_1 _0646_ (.A(_0155_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _0647_ (.A(_0152_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__and2b_1 _0648_ (.A_N(\manchester_baby_instance.ram_data_o_15 ),
    .B(\manchester_baby_instance.ram_data_i_15 ),
    .X(_0161_));
 sky130_fd_sc_hd__or2b_1 _0649_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B_N(\manchester_baby_instance.ram_data_o_14 ),
    .X(_0162_));
 sky130_fd_sc_hd__or2b_1 _0650_ (.A(\manchester_baby_instance.ram_data_i_12 ),
    .B_N(\manchester_baby_instance.ram_data_o_12 ),
    .X(_0163_));
 sky130_fd_sc_hd__a211o_1 _0651_ (.A1(_0163_),
    .A2(_0147_),
    .B1(_0146_),
    .C1(_0143_),
    .X(_0164_));
 sky130_fd_sc_hd__inv_2 _0652_ (.A(\manchester_baby_instance.ram_data_i_11 ),
    .Y(_0165_));
 sky130_fd_sc_hd__a21boi_1 _0653_ (.A1(_0153_),
    .A2(_0156_),
    .B1_N(_0157_),
    .Y(_0166_));
 sky130_fd_sc_hd__and2b_1 _0654_ (.A_N(\manchester_baby_instance.ram_data_i_10 ),
    .B(\manchester_baby_instance.ram_data_o_10 ),
    .X(_0167_));
 sky130_fd_sc_hd__o21a_1 _0655_ (.A1(\manchester_baby_instance.ram_data_o_11 ),
    .A2(_0165_),
    .B1(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__a221o_1 _0656_ (.A1(\manchester_baby_instance.ram_data_o_11 ),
    .A2(_0165_),
    .B1(_0152_),
    .B2(_0166_),
    .C1(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__or2b_1 _0657_ (.A(_0149_),
    .B_N(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__or2b_1 _0658_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B_N(\manchester_baby_instance.ram_data_o_15 ),
    .X(_0171_));
 sky130_fd_sc_hd__o2111a_1 _0659_ (.A1(_0161_),
    .A2(_0162_),
    .B1(_0164_),
    .C1(_0170_),
    .D1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__o31a_2 _0660_ (.A1(_0140_),
    .A2(_0149_),
    .A3(_0160_),
    .B1(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__xnor2_2 _0661_ (.A(\manchester_baby_instance.ram_data_o_16 ),
    .B(\manchester_baby_instance.ram_data_i_16 ),
    .Y(_0174_));
 sky130_fd_sc_hd__and2b_1 _0662_ (.A_N(_0173_),
    .B(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _0663_ (.A(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__and2b_1 _0664_ (.A_N(\manchester_baby_instance.ram_data_o_17 ),
    .B(\manchester_baby_instance.ram_data_i_17 ),
    .X(_0177_));
 sky130_fd_sc_hd__xnor2_1 _0665_ (.A(\manchester_baby_instance.ram_data_o_18 ),
    .B(\manchester_baby_instance.ram_data_i_18 ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _0666_ (.A(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__a311o_1 _0667_ (.A1(_0107_),
    .A2(_0108_),
    .A3(_0176_),
    .B1(_0177_),
    .C1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__and2b_1 _0668_ (.A_N(_0177_),
    .B(_0107_),
    .X(_0181_));
 sky130_fd_sc_hd__a21oi_1 _0669_ (.A1(_0107_),
    .A2(_0108_),
    .B1(_0177_),
    .Y(_0182_));
 sky130_fd_sc_hd__a211o_1 _0670_ (.A1(_0181_),
    .A2(_0175_),
    .B1(_0178_),
    .C1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__or4_1 _0671_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B(\manchester_baby_instance.ram_data_i_2 ),
    .C(\manchester_baby_instance.ram_data_i_1 ),
    .D(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0184_));
 sky130_fd_sc_hd__or4_1 _0672_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(\manchester_baby_instance.ram_data_i_5 ),
    .C(\manchester_baby_instance.ram_data_i_6 ),
    .D(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or4_1 _0673_ (.A(\manchester_baby_instance.ram_data_i_7 ),
    .B(\manchester_baby_instance.ram_data_i_8 ),
    .C(\manchester_baby_instance.ram_data_i_9 ),
    .D(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__or4_2 _0674_ (.A(\manchester_baby_instance.ram_data_i_10 ),
    .B(\manchester_baby_instance.ram_data_i_11 ),
    .C(\manchester_baby_instance.ram_data_i_12 ),
    .D(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__or2_1 _0675_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__or2_1 _0676_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(\manchester_baby_instance.ram_data_i_14 ),
    .X(_0189_));
 sky130_fd_sc_hd__or2_1 _0677_ (.A(_0188_),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__or2_1 _0678_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _0679_ (.A(\manchester_baby_instance.ram_data_i_17 ),
    .B(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__xor2_1 _0680_ (.A(\manchester_baby_instance.ram_data_i_18 ),
    .B(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__and4bb_2 _0681_ (.A_N(_0104_),
    .B_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .C(_0103_),
    .D(_0101_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_4 _0682_ (.A(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_4 _0683_ (.A(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__a32o_1 _0684_ (.A1(_0106_),
    .A2(_0180_),
    .A3(_0183_),
    .B1(_0193_),
    .B2(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__o21a_2 _0685_ (.A1(_0106_),
    .A2(_0194_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_4 _0686_ (.A(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _0687_ (.A0(\manchester_baby_instance.ram_data_o_18 ),
    .A1(_0197_),
    .S(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0200_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _0689_ (.A(\manchester_baby_instance.ram_data_i_17 ),
    .B(_0191_),
    .Y(_0201_));
 sky130_fd_sc_hd__and2_1 _0690_ (.A(_0108_),
    .B(_0176_),
    .X(_0202_));
 sky130_fd_sc_hd__xnor2_1 _0691_ (.A(_0181_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__clkbuf_4 _0692_ (.A(_0106_),
    .X(_0204_));
 sky130_fd_sc_hd__a32o_1 _0693_ (.A1(_0196_),
    .A2(_0192_),
    .A3(_0201_),
    .B1(_0203_),
    .B2(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(\manchester_baby_instance.ram_data_o_17 ),
    .A1(_0205_),
    .S(_0199_),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _0695_ (.A(_0206_),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_1 _0696_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(_0190_),
    .Y(_0207_));
 sky130_fd_sc_hd__xnor2_1 _0697_ (.A(_0174_),
    .B(_0173_),
    .Y(_0208_));
 sky130_fd_sc_hd__a32o_1 _0698_ (.A1(_0196_),
    .A2(_0191_),
    .A3(_0207_),
    .B1(_0208_),
    .B2(_0204_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _0699_ (.A0(\manchester_baby_instance.ram_data_o_16 ),
    .A1(_0209_),
    .S(_0199_),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0210_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _0701_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B(_0188_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__and2b_1 _0703_ (.A_N(\manchester_baby_instance.ram_data_o_14 ),
    .B(\manchester_baby_instance.ram_data_i_14 ),
    .X(_0213_));
 sky130_fd_sc_hd__nor2_1 _0704_ (.A(_0140_),
    .B(_0160_),
    .Y(_0214_));
 sky130_fd_sc_hd__o21a_1 _0705_ (.A1(_0169_),
    .A2(_0214_),
    .B1(_0144_),
    .X(_0215_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__a31o_1 _0707_ (.A1(_0163_),
    .A2(_0147_),
    .A3(_0216_),
    .B1(_0146_),
    .X(_0217_));
 sky130_fd_sc_hd__o21a_1 _0708_ (.A1(_0213_),
    .A2(_0217_),
    .B1(_0162_),
    .X(_0218_));
 sky130_fd_sc_hd__xnor2_1 _0709_ (.A(_0141_),
    .B(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__a32o_1 _0710_ (.A1(_0196_),
    .A2(_0190_),
    .A3(_0212_),
    .B1(_0219_),
    .B2(_0204_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(\manchester_baby_instance.ram_data_o_15 ),
    .A1(_0220_),
    .S(_0199_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0221_),
    .X(_0097_));
 sky130_fd_sc_hd__nand2_1 _0713_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B(_0188_),
    .Y(_0222_));
 sky130_fd_sc_hd__xnor2_1 _0714_ (.A(_0142_),
    .B(_0217_),
    .Y(_0223_));
 sky130_fd_sc_hd__a32o_1 _0715_ (.A1(_0196_),
    .A2(_0211_),
    .A3(_0222_),
    .B1(_0223_),
    .B2(_0204_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _0716_ (.A0(\manchester_baby_instance.ram_data_o_14 ),
    .A1(_0224_),
    .S(_0199_),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_1 _0717_ (.A(_0225_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _0718_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B(_0187_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _0719_ (.A(_0163_),
    .B(_0216_),
    .Y(_0227_));
 sky130_fd_sc_hd__xnor2_1 _0720_ (.A(_0148_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__clkbuf_4 _0721_ (.A(_0106_),
    .X(_0229_));
 sky130_fd_sc_hd__a32o_1 _0722_ (.A1(_0196_),
    .A2(_0188_),
    .A3(_0226_),
    .B1(_0228_),
    .B2(_0229_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(\manchester_baby_instance.ram_data_o_13 ),
    .A1(_0230_),
    .S(_0199_),
    .X(_0231_));
 sky130_fd_sc_hd__clkbuf_1 _0724_ (.A(_0231_),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _0725_ (.A(\manchester_baby_instance.ram_data_i_10 ),
    .B(_0186_),
    .X(_0232_));
 sky130_fd_sc_hd__or2_1 _0726_ (.A(\manchester_baby_instance.ram_data_i_11 ),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _0727_ (.A(\manchester_baby_instance.ram_data_i_12 ),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__nor2_1 _0728_ (.A(_0169_),
    .B(_0214_),
    .Y(_0235_));
 sky130_fd_sc_hd__xnor2_1 _0729_ (.A(_0144_),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__a32o_1 _0730_ (.A1(_0196_),
    .A2(_0187_),
    .A3(_0234_),
    .B1(_0236_),
    .B2(_0229_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _0731_ (.A0(\manchester_baby_instance.ram_data_o_12 ),
    .A1(_0237_),
    .S(_0199_),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _0732_ (.A(_0238_),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _0733_ (.A(_0195_),
    .X(_0239_));
 sky130_fd_sc_hd__nand2_1 _0734_ (.A(\manchester_baby_instance.ram_data_i_11 ),
    .B(_0232_),
    .Y(_0240_));
 sky130_fd_sc_hd__and2b_1 _0735_ (.A_N(\manchester_baby_instance.ram_data_o_10 ),
    .B(\manchester_baby_instance.ram_data_i_10 ),
    .X(_0241_));
 sky130_fd_sc_hd__nor2_1 _0736_ (.A(_0140_),
    .B(_0155_),
    .Y(_0242_));
 sky130_fd_sc_hd__a31oi_2 _0737_ (.A1(_0156_),
    .A2(_0157_),
    .A3(_0242_),
    .B1(_0166_),
    .Y(_0243_));
 sky130_fd_sc_hd__o21ba_1 _0738_ (.A1(_0241_),
    .A2(_0243_),
    .B1_N(_0167_),
    .X(_0244_));
 sky130_fd_sc_hd__xnor2_1 _0739_ (.A(_0150_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a32o_1 _0740_ (.A1(_0239_),
    .A2(_0233_),
    .A3(_0240_),
    .B1(_0245_),
    .B2(_0229_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _0741_ (.A0(\manchester_baby_instance.ram_data_o_11 ),
    .A1(_0246_),
    .S(_0199_),
    .X(_0247_));
 sky130_fd_sc_hd__clkbuf_1 _0742_ (.A(_0247_),
    .X(_0093_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(\manchester_baby_instance.ram_data_i_10 ),
    .B(_0186_),
    .Y(_0248_));
 sky130_fd_sc_hd__xnor2_1 _0744_ (.A(_0151_),
    .B(_0243_),
    .Y(_0249_));
 sky130_fd_sc_hd__a32o_1 _0745_ (.A1(_0239_),
    .A2(_0232_),
    .A3(_0248_),
    .B1(_0249_),
    .B2(_0229_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_4 _0746_ (.A(_0198_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _0747_ (.A0(\manchester_baby_instance.ram_data_o_10 ),
    .A1(_0250_),
    .S(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__clkbuf_1 _0748_ (.A(_0252_),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0749_ (.A(\manchester_baby_instance.ram_data_i_7 ),
    .B(_0185_),
    .X(_0253_));
 sky130_fd_sc_hd__or2_1 _0750_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B(_0253_),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _0751_ (.A(\manchester_baby_instance.ram_data_i_9 ),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__o21ai_1 _0752_ (.A1(_0140_),
    .A2(_0155_),
    .B1(_0153_),
    .Y(_0256_));
 sky130_fd_sc_hd__xnor2_1 _0753_ (.A(_0158_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__a32o_1 _0754_ (.A1(_0239_),
    .A2(_0186_),
    .A3(_0255_),
    .B1(_0257_),
    .B2(_0229_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _0755_ (.A0(\manchester_baby_instance.ram_data_o_9 ),
    .A1(_0258_),
    .S(_0251_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_1 _0756_ (.A(_0259_),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_1 _0757_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B(_0253_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand3b_4 _0758_ (.A_N(_0101_),
    .B(_0103_),
    .C(_0104_),
    .Y(_0261_));
 sky130_fd_sc_hd__nor2_1 _0759_ (.A(_0261_),
    .B(_0242_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand2_1 _0760_ (.A(_0140_),
    .B(_0155_),
    .Y(_0263_));
 sky130_fd_sc_hd__a32o_1 _0761_ (.A1(_0239_),
    .A2(_0254_),
    .A3(_0260_),
    .B1(_0262_),
    .B2(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(\manchester_baby_instance.ram_data_o_8 ),
    .A1(_0264_),
    .S(_0251_),
    .X(_0265_));
 sky130_fd_sc_hd__clkbuf_1 _0763_ (.A(_0265_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _0764_ (.A(\manchester_baby_instance.ram_data_i_7 ),
    .B(_0185_),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_2 _0765_ (.A(_0112_),
    .Y(_0267_));
 sky130_fd_sc_hd__a21oi_1 _0766_ (.A1(_0116_),
    .A2(_0133_),
    .B1(_0135_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_1 _0767_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_0136_),
    .Y(_0269_));
 sky130_fd_sc_hd__xnor2_1 _0768_ (.A(_0111_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(_0261_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__a31o_1 _0770_ (.A1(_0196_),
    .A2(_0253_),
    .A3(_0266_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(\manchester_baby_instance.ram_data_o_7 ),
    .A1(_0272_),
    .S(_0251_),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(_0273_),
    .X(_0089_));
 sky130_fd_sc_hd__xnor2_1 _0773_ (.A(_0112_),
    .B(_0268_),
    .Y(_0274_));
 sky130_fd_sc_hd__or2_1 _0774_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0184_),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _0775_ (.A(\manchester_baby_instance.ram_data_i_5 ),
    .B(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__nand2_1 _0776_ (.A(\manchester_baby_instance.ram_data_i_6 ),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__and3_1 _0777_ (.A(_0195_),
    .B(_0185_),
    .C(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__a21o_1 _0778_ (.A1(_0204_),
    .A2(_0274_),
    .B1(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _0779_ (.A0(\manchester_baby_instance.ram_data_o_6 ),
    .A1(_0279_),
    .S(_0251_),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_1 _0780_ (.A(_0280_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(\manchester_baby_instance.ram_data_i_5 ),
    .B(_0275_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _0782_ (.A(_0121_),
    .B(_0131_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0783_ (.A(_0132_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _0784_ (.A(_0134_),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__xor2_1 _0785_ (.A(_0116_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__a32o_1 _0786_ (.A1(_0239_),
    .A2(_0276_),
    .A3(_0281_),
    .B1(_0285_),
    .B2(_0229_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _0787_ (.A0(\manchester_baby_instance.ram_data_o_5 ),
    .A1(_0286_),
    .S(_0251_),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_1 _0788_ (.A(_0287_),
    .X(_0087_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(_0132_),
    .B(_0282_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0184_),
    .Y(_0289_));
 sky130_fd_sc_hd__and3_1 _0791_ (.A(_0195_),
    .B(_0275_),
    .C(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__a31o_1 _0792_ (.A1(_0204_),
    .A2(_0283_),
    .A3(_0288_),
    .B1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _0793_ (.A0(\manchester_baby_instance.ram_data_o_4 ),
    .A1(_0291_),
    .S(_0251_),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_1 _0794_ (.A(_0292_),
    .X(_0086_));
 sky130_fd_sc_hd__or2_1 _0795_ (.A(\manchester_baby_instance.ram_data_i_1 ),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _0796_ (.A(_0118_),
    .B(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__nand2_1 _0797_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_1 _0798_ (.A1(_0124_),
    .A2(_0128_),
    .B1(_0122_),
    .Y(_0296_));
 sky130_fd_sc_hd__xnor2_1 _0799_ (.A(_0296_),
    .B(_0130_),
    .Y(_0297_));
 sky130_fd_sc_hd__a32o_1 _0800_ (.A1(_0239_),
    .A2(_0184_),
    .A3(_0295_),
    .B1(_0297_),
    .B2(_0229_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _0801_ (.A0(\manchester_baby_instance.ram_data_o_3 ),
    .A1(_0298_),
    .S(_0251_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(_0299_),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_1 _0803_ (.A(_0118_),
    .B(_0293_),
    .Y(_0300_));
 sky130_fd_sc_hd__xor2_1 _0804_ (.A(_0124_),
    .B(_0128_),
    .X(_0301_));
 sky130_fd_sc_hd__a32o_1 _0805_ (.A1(_0239_),
    .A2(_0294_),
    .A3(_0300_),
    .B1(_0301_),
    .B2(_0229_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(\manchester_baby_instance.ram_data_o_2 ),
    .A1(_0302_),
    .S(_0251_),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _0807_ (.A(_0303_),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_1 _0808_ (.A(\manchester_baby_instance.ram_data_i_1 ),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .Y(_0304_));
 sky130_fd_sc_hd__or2b_1 _0809_ (.A(_0127_),
    .B_N(_0125_),
    .X(_0305_));
 sky130_fd_sc_hd__xnor2_1 _0810_ (.A(_0305_),
    .B(_0126_),
    .Y(_0306_));
 sky130_fd_sc_hd__a32o_1 _0811_ (.A1(_0239_),
    .A2(_0293_),
    .A3(_0304_),
    .B1(_0306_),
    .B2(_0229_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(\manchester_baby_instance.ram_data_o_1 ),
    .A1(_0307_),
    .S(_0251_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _0813_ (.A(_0308_),
    .X(_0083_));
 sky130_fd_sc_hd__or2b_1 _0814_ (.A(_0196_),
    .B_N(\manchester_baby_instance.ram_data_o_0 ),
    .X(_0309_));
 sky130_fd_sc_hd__o21ai_1 _0815_ (.A1(\manchester_baby_instance.ram_data_i_0 ),
    .A2(_0261_),
    .B1(_0199_),
    .Y(_0310_));
 sky130_fd_sc_hd__a32o_1 _0816_ (.A1(\manchester_baby_instance.ram_data_i_0 ),
    .A2(_0199_),
    .A3(_0309_),
    .B1(_0310_),
    .B2(net25),
    .X(_0082_));
 sky130_fd_sc_hd__and3b_1 _0817_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(_0104_),
    .B(_0101_),
    .Y(_0312_));
 sky130_fd_sc_hd__and2_1 _0819_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_1 _0820_ (.A(_0312_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__and2b_1 _0821_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0102_),
    .X(_0315_));
 sky130_fd_sc_hd__o21a_1 _0822_ (.A1(_0311_),
    .A2(_0315_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0316_));
 sky130_fd_sc_hd__a21bo_1 _0823_ (.A1(_0311_),
    .A2(_0314_),
    .B1_N(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__nor2_1 _0824_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0118_),
    .Y(_0318_));
 sky130_fd_sc_hd__buf_2 _0825_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .X(_0319_));
 sky130_fd_sc_hd__xnor2_1 _0826_ (.A(_0319_),
    .B(\manchester_baby_instance.ram_data_i_1 ),
    .Y(_0320_));
 sky130_fd_sc_hd__nand2_1 _0827_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .Y(_0321_));
 sky130_fd_sc_hd__or2_1 _0828_ (.A(_0320_),
    .B(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__a21boi_1 _0829_ (.A1(_0319_),
    .A2(\manchester_baby_instance.ram_data_i_1 ),
    .B1_N(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_1 _0830_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0118_),
    .Y(_0324_));
 sky130_fd_sc_hd__o21ai_1 _0831_ (.A1(_0318_),
    .A2(_0323_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__o21a_1 _0832_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(\manchester_baby_instance.ram_data_i_3 ),
    .B1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__a21o_1 _0833_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(\manchester_baby_instance.ram_data_i_3 ),
    .B1(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_1 _0834_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__and2_1 _0835_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _0836_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0328_),
    .Y(_0330_));
 sky130_fd_sc_hd__clkbuf_4 _0837_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _0838_ (.A(_0331_),
    .B(_0311_),
    .C(_0312_),
    .X(_0332_));
 sky130_fd_sc_hd__o21a_1 _0839_ (.A1(_0329_),
    .A2(_0330_),
    .B1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__and3b_1 _0840_ (.A_N(_0331_),
    .B(_0311_),
    .C(_0313_),
    .X(_0334_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .Y(_0335_));
 sky130_fd_sc_hd__o21a_1 _0842_ (.A1(_0315_),
    .A2(_0334_),
    .B1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__buf_2 _0843_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .X(_0337_));
 sky130_fd_sc_hd__and3_1 _0844_ (.A(_0319_),
    .B(_0337_),
    .C(\manchester_baby_instance.ram_data_o_31 ),
    .X(_0338_));
 sky130_fd_sc_hd__a21boi_1 _0845_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0338_),
    .B1_N(_0334_),
    .Y(_0339_));
 sky130_fd_sc_hd__and3_1 _0846_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0319_),
    .C(_0337_),
    .X(_0340_));
 sky130_fd_sc_hd__and2b_1 _0847_ (.A_N(_0340_),
    .B(_0315_),
    .X(_0341_));
 sky130_fd_sc_hd__o31a_1 _0848_ (.A1(_0336_),
    .A2(_0339_),
    .A3(_0341_),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .X(_0342_));
 sky130_fd_sc_hd__and3b_1 _0849_ (.A_N(_0331_),
    .B(_0311_),
    .C(_0312_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _0850_ (.A1(\manchester_baby_instance.ram_data_o_31 ),
    .A2(_0334_),
    .B1(_0315_),
    .X(_0344_));
 sky130_fd_sc_hd__and4b_1 _0851_ (.A_N(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .C(_0340_),
    .D(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__a21oi_1 _0852_ (.A1(\manchester_baby_instance.ram_data_i_4 ),
    .A2(_0343_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__or3b_1 _0853_ (.A(_0333_),
    .B(_0342_),
    .C_N(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _0854_ (.A1(net26),
    .A2(_0317_),
    .B1(_0347_),
    .B2(_0316_),
    .X(_0081_));
 sky130_fd_sc_hd__xnor2_1 _0855_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .B(\manchester_baby_instance.ram_data_i_3 ),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_1 _0856_ (.A(_0325_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a22o_1 _0857_ (.A1(\manchester_baby_instance.ram_data_i_3 ),
    .A2(_0343_),
    .B1(_0349_),
    .B2(_0332_),
    .X(_0350_));
 sky130_fd_sc_hd__a31o_1 _0858_ (.A1(_0335_),
    .A2(_0340_),
    .A3(_0344_),
    .B1(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__or3_1 _0859_ (.A(_0317_),
    .B(_0339_),
    .C(_0341_),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _0860_ (.A1(_0316_),
    .A2(_0351_),
    .B1(_0352_),
    .B2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .X(_0080_));
 sky130_fd_sc_hd__a21o_1 _0861_ (.A1(_0319_),
    .A2(_0337_),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _0862_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0118_),
    .X(_0354_));
 sky130_fd_sc_hd__nand2_1 _0863_ (.A(_0324_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__xor2_1 _0864_ (.A(_0323_),
    .B(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _0865_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0338_),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _0866_ (.A1(_0332_),
    .A2(_0356_),
    .B1(_0357_),
    .B2(_0339_),
    .X(_0358_));
 sky130_fd_sc_hd__a221o_1 _0867_ (.A1(_0118_),
    .A2(_0343_),
    .B1(_0353_),
    .B2(_0341_),
    .C1(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0317_),
    .B1(_0359_),
    .B2(_0316_),
    .X(_0079_));
 sky130_fd_sc_hd__a21oi_1 _0869_ (.A1(_0337_),
    .A2(\manchester_baby_instance.ram_data_o_31 ),
    .B1(_0319_),
    .Y(_0360_));
 sky130_fd_sc_hd__nor2_1 _0870_ (.A(_0338_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _0871_ (.A(_0320_),
    .B(_0321_),
    .Y(_0362_));
 sky130_fd_sc_hd__xor2_1 _0872_ (.A(_0319_),
    .B(_0337_),
    .X(_0363_));
 sky130_fd_sc_hd__a32o_1 _0873_ (.A1(_0332_),
    .A2(_0322_),
    .A3(_0362_),
    .B1(_0363_),
    .B2(_0315_),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _0874_ (.A1(\manchester_baby_instance.ram_data_i_1 ),
    .A2(_0343_),
    .B1(_0361_),
    .B2(_0334_),
    .C1(_0364_),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _0875_ (.A1(_0319_),
    .A2(_0317_),
    .B1(_0365_),
    .B2(_0316_),
    .X(_0078_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(_0337_),
    .Y(_0366_));
 sky130_fd_sc_hd__and3b_1 _0877_ (.A_N(\manchester_baby_instance.ram_data_o_31 ),
    .B(_0334_),
    .C(_0337_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _0878_ (.A(_0337_),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0368_));
 sky130_fd_sc_hd__a32o_1 _0879_ (.A1(_0332_),
    .A2(_0321_),
    .A3(_0368_),
    .B1(_0343_),
    .B2(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0369_));
 sky130_fd_sc_hd__a211o_1 _0880_ (.A1(_0366_),
    .A2(_0344_),
    .B1(_0367_),
    .C1(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _0881_ (.A1(_0337_),
    .A2(_0317_),
    .B1(_0370_),
    .B2(_0316_),
    .X(_0077_));
 sky130_fd_sc_hd__a41o_1 _0882_ (.A1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .A2(_0331_),
    .A3(_0103_),
    .A4(_0313_),
    .B1(net22),
    .X(_0072_));
 sky130_fd_sc_hd__inv_2 _0883_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ));
 sky130_fd_sc_hd__and4b_1 _0884_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .X(_0371_));
 sky130_fd_sc_hd__buf_2 _0885_ (.A(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(_0104_),
    .A1(\manchester_baby_instance.ram_data_i_15 ),
    .S(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0887_ (.A(_0373_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(_0101_),
    .A1(\manchester_baby_instance.ram_data_i_14 ),
    .S(_0372_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0374_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0890_ (.A0(_0331_),
    .A1(\manchester_baby_instance.ram_data_i_13 ),
    .S(_0372_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0891_ (.A(_0375_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(net30),
    .A1(\manchester_baby_instance.ram_data_i_4 ),
    .S(_0372_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0376_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(net29),
    .A1(\manchester_baby_instance.ram_data_i_3 ),
    .S(_0372_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0377_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(net27),
    .A1(_0118_),
    .S(_0372_),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0378_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(net28),
    .A1(\manchester_baby_instance.ram_data_i_1 ),
    .S(_0372_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0379_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(net31),
    .A1(\manchester_baby_instance.ram_data_i_0 ),
    .S(_0372_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0380_),
    .X(_0063_));
 sky130_fd_sc_hd__and2b_1 _0902_ (.A_N(\manchester_baby_instance.ram_data_i_30 ),
    .B(\manchester_baby_instance.ram_data_o_30 ),
    .X(_0381_));
 sky130_fd_sc_hd__and2b_1 _0903_ (.A_N(\manchester_baby_instance.ram_data_i_28 ),
    .B(\manchester_baby_instance.ram_data_o_28 ),
    .X(_0382_));
 sky130_fd_sc_hd__or2b_1 _0904_ (.A(\manchester_baby_instance.ram_data_i_24 ),
    .B_N(\manchester_baby_instance.ram_data_o_24 ),
    .X(_0383_));
 sky130_fd_sc_hd__or2b_1 _0905_ (.A(\manchester_baby_instance.ram_data_o_24 ),
    .B_N(\manchester_baby_instance.ram_data_i_24 ),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(_0383_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__and2b_1 _0907_ (.A_N(\manchester_baby_instance.ram_data_o_21 ),
    .B(\manchester_baby_instance.ram_data_i_21 ),
    .X(_0386_));
 sky130_fd_sc_hd__or2b_1 _0908_ (.A(\manchester_baby_instance.ram_data_i_21 ),
    .B_N(\manchester_baby_instance.ram_data_o_21 ),
    .X(_0387_));
 sky130_fd_sc_hd__and2b_1 _0909_ (.A_N(_0386_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0910_ (.A(\manchester_baby_instance.ram_data_o_20 ),
    .B(\manchester_baby_instance.ram_data_i_20 ),
    .Y(_0389_));
 sky130_fd_sc_hd__nand2_1 _0911_ (.A(_0388_),
    .B(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__and2b_1 _0912_ (.A_N(\manchester_baby_instance.ram_data_o_22 ),
    .B(\manchester_baby_instance.ram_data_i_22 ),
    .X(_0391_));
 sky130_fd_sc_hd__or2b_1 _0913_ (.A(\manchester_baby_instance.ram_data_i_22 ),
    .B_N(\manchester_baby_instance.ram_data_o_22 ),
    .X(_0392_));
 sky130_fd_sc_hd__or2b_1 _0914_ (.A(_0391_),
    .B_N(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__and2b_1 _0915_ (.A_N(\manchester_baby_instance.ram_data_o_23 ),
    .B(\manchester_baby_instance.ram_data_i_23 ),
    .X(_0394_));
 sky130_fd_sc_hd__or2b_1 _0916_ (.A(\manchester_baby_instance.ram_data_i_23 ),
    .B_N(\manchester_baby_instance.ram_data_o_23 ),
    .X(_0395_));
 sky130_fd_sc_hd__or2b_1 _0917_ (.A(_0394_),
    .B_N(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__or3_1 _0918_ (.A(_0390_),
    .B(_0393_),
    .C(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__xnor2_1 _0919_ (.A(\manchester_baby_instance.ram_data_o_19 ),
    .B(\manchester_baby_instance.ram_data_i_19 ),
    .Y(_0398_));
 sky130_fd_sc_hd__and2_1 _0920_ (.A(_0178_),
    .B(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__nand3_1 _0921_ (.A(_0181_),
    .B(_0174_),
    .C(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__or2b_1 _0922_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B_N(\manchester_baby_instance.ram_data_o_20 ),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _0923_ (.A(\manchester_baby_instance.ram_data_i_19 ),
    .Y(_0402_));
 sky130_fd_sc_hd__and2b_1 _0924_ (.A_N(\manchester_baby_instance.ram_data_i_18 ),
    .B(\manchester_baby_instance.ram_data_o_18 ),
    .X(_0403_));
 sky130_fd_sc_hd__o21a_1 _0925_ (.A1(\manchester_baby_instance.ram_data_o_19 ),
    .A2(_0402_),
    .B1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__a221o_1 _0926_ (.A1(\manchester_baby_instance.ram_data_o_19 ),
    .A2(_0402_),
    .B1(_0182_),
    .B2(_0399_),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _0927_ (.A(_0405_),
    .B(_0389_),
    .Y(_0406_));
 sky130_fd_sc_hd__a311o_1 _0928_ (.A1(_0387_),
    .A2(_0401_),
    .A3(_0406_),
    .B1(_0386_),
    .C1(_0391_),
    .X(_0407_));
 sky130_fd_sc_hd__a31o_1 _0929_ (.A1(_0407_),
    .A2(_0395_),
    .A3(_0392_),
    .B1(_0394_),
    .X(_0408_));
 sky130_fd_sc_hd__o31a_1 _0930_ (.A1(_0173_),
    .A2(_0397_),
    .A3(_0400_),
    .B1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__and2b_1 _0931_ (.A_N(\manchester_baby_instance.ram_data_o_25 ),
    .B(\manchester_baby_instance.ram_data_i_25 ),
    .X(_0410_));
 sky130_fd_sc_hd__or2b_1 _0932_ (.A(\manchester_baby_instance.ram_data_i_25 ),
    .B_N(\manchester_baby_instance.ram_data_o_25 ),
    .X(_0411_));
 sky130_fd_sc_hd__or2b_1 _0933_ (.A(_0410_),
    .B_N(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__and2b_1 _0934_ (.A_N(\manchester_baby_instance.ram_data_i_27 ),
    .B(\manchester_baby_instance.ram_data_o_27 ),
    .X(_0413_));
 sky130_fd_sc_hd__and2b_1 _0935_ (.A_N(\manchester_baby_instance.ram_data_o_27 ),
    .B(\manchester_baby_instance.ram_data_i_27 ),
    .X(_0414_));
 sky130_fd_sc_hd__or2_1 _0936_ (.A(_0413_),
    .B(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__or2b_1 _0937_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B_N(\manchester_baby_instance.ram_data_o_26 ),
    .X(_0416_));
 sky130_fd_sc_hd__or2b_1 _0938_ (.A(\manchester_baby_instance.ram_data_o_26 ),
    .B_N(\manchester_baby_instance.ram_data_i_26 ),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _0940_ (.A(_0415_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__or4_1 _0941_ (.A(_0385_),
    .B(_0409_),
    .C(_0412_),
    .D(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _0942_ (.A1(_0383_),
    .A2(_0411_),
    .B1(_0410_),
    .X(_0421_));
 sky130_fd_sc_hd__o21ba_1 _0943_ (.A1(_0414_),
    .A2(_0416_),
    .B1_N(_0413_),
    .X(_0422_));
 sky130_fd_sc_hd__o21a_1 _0944_ (.A1(_0419_),
    .A2(_0421_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__and2b_1 _0945_ (.A_N(\manchester_baby_instance.ram_data_o_28 ),
    .B(\manchester_baby_instance.ram_data_i_28 ),
    .X(_0424_));
 sky130_fd_sc_hd__or2_1 _0946_ (.A(_0382_),
    .B(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__a21oi_2 _0947_ (.A1(_0420_),
    .A2(_0423_),
    .B1(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__and2b_1 _0948_ (.A_N(\manchester_baby_instance.ram_data_i_29 ),
    .B(\manchester_baby_instance.ram_data_o_29 ),
    .X(_0427_));
 sky130_fd_sc_hd__or2b_1 _0949_ (.A(\manchester_baby_instance.ram_data_o_29 ),
    .B_N(\manchester_baby_instance.ram_data_i_29 ),
    .X(_0428_));
 sky130_fd_sc_hd__and2b_1 _0950_ (.A_N(\manchester_baby_instance.ram_data_o_30 ),
    .B(\manchester_baby_instance.ram_data_i_30 ),
    .X(_0429_));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(_0381_),
    .B(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__inv_2 _0952_ (.A(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__o311a_1 _0953_ (.A1(_0382_),
    .A2(_0426_),
    .A3(_0427_),
    .B1(_0428_),
    .C1(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__nor2_1 _0954_ (.A(\manchester_baby_instance.ram_data_o_31 ),
    .B(\manchester_baby_instance.ram_data_i_31 ),
    .Y(_0433_));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(\manchester_baby_instance.ram_data_o_31 ),
    .B(\manchester_baby_instance.ram_data_i_31 ),
    .X(_0434_));
 sky130_fd_sc_hd__or4_1 _0956_ (.A(_0381_),
    .B(_0432_),
    .C(_0433_),
    .D(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__o22ai_1 _0957_ (.A1(_0381_),
    .A2(_0432_),
    .B1(_0433_),
    .B2(_0434_),
    .Y(_0436_));
 sky130_fd_sc_hd__or4_1 _0958_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(\manchester_baby_instance.ram_data_i_17 ),
    .C(\manchester_baby_instance.ram_data_i_18 ),
    .D(\manchester_baby_instance.ram_data_i_19 ),
    .X(_0437_));
 sky130_fd_sc_hd__or4_2 _0959_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B(_0187_),
    .C(_0189_),
    .D(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__or4_1 _0960_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B(\manchester_baby_instance.ram_data_i_21 ),
    .C(\manchester_baby_instance.ram_data_i_22 ),
    .D(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__or4_1 _0961_ (.A(\manchester_baby_instance.ram_data_i_23 ),
    .B(\manchester_baby_instance.ram_data_i_24 ),
    .C(\manchester_baby_instance.ram_data_i_25 ),
    .D(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__or3_1 _0962_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B(\manchester_baby_instance.ram_data_i_27 ),
    .C(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__or3_1 _0963_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .B(\manchester_baby_instance.ram_data_i_29 ),
    .C(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__or2_1 _0964_ (.A(\manchester_baby_instance.ram_data_i_30 ),
    .B(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__xor2_1 _0965_ (.A(\manchester_baby_instance.ram_data_i_31 ),
    .B(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__a32o_1 _0966_ (.A1(_0106_),
    .A2(_0435_),
    .A3(_0436_),
    .B1(_0196_),
    .B2(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_4 _0967_ (.A(_0198_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(\manchester_baby_instance.ram_data_o_31 ),
    .A1(_0445_),
    .S(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0969_ (.A(_0447_),
    .X(_0062_));
 sky130_fd_sc_hd__nand2_1 _0970_ (.A(\manchester_baby_instance.ram_data_i_30 ),
    .B(_0442_),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2_1 _0971_ (.A(_0261_),
    .B(_0432_),
    .Y(_0449_));
 sky130_fd_sc_hd__o31a_1 _0972_ (.A1(_0382_),
    .A2(_0426_),
    .A3(_0427_),
    .B1(_0428_),
    .X(_0450_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(_0431_),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__a32o_1 _0974_ (.A1(_0239_),
    .A2(_0443_),
    .A3(_0448_),
    .B1(_0449_),
    .B2(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _0975_ (.A0(\manchester_baby_instance.ram_data_o_30 ),
    .A1(_0452_),
    .S(_0446_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0976_ (.A(_0453_),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _0977_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .B(_0441_),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _0978_ (.A(\manchester_baby_instance.ram_data_i_29 ),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__and2b_1 _0979_ (.A_N(\manchester_baby_instance.ram_data_o_29 ),
    .B(\manchester_baby_instance.ram_data_i_29 ),
    .X(_0456_));
 sky130_fd_sc_hd__o22a_1 _0980_ (.A1(_0382_),
    .A2(_0426_),
    .B1(_0427_),
    .B2(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__or4_1 _0981_ (.A(_0456_),
    .B(_0382_),
    .C(_0426_),
    .D(_0427_),
    .X(_0458_));
 sky130_fd_sc_hd__or2b_1 _0982_ (.A(_0457_),
    .B_N(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__a32o_1 _0983_ (.A1(_0239_),
    .A2(_0442_),
    .A3(_0455_),
    .B1(_0459_),
    .B2(_0229_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(\manchester_baby_instance.ram_data_o_29 ),
    .A1(_0460_),
    .S(_0446_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0985_ (.A(_0461_),
    .X(_0060_));
 sky130_fd_sc_hd__nand2_1 _0986_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .B(_0441_),
    .Y(_0462_));
 sky130_fd_sc_hd__and3_1 _0987_ (.A(_0425_),
    .B(_0420_),
    .C(_0423_),
    .X(_0463_));
 sky130_fd_sc_hd__nor2_1 _0988_ (.A(_0426_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__a32o_1 _0989_ (.A1(_0195_),
    .A2(_0454_),
    .A3(_0462_),
    .B1(_0464_),
    .B2(_0106_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _0990_ (.A0(\manchester_baby_instance.ram_data_o_28 ),
    .A1(_0465_),
    .S(_0446_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0991_ (.A(_0466_),
    .X(_0059_));
 sky130_fd_sc_hd__or2_1 _0992_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B(_0440_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _0993_ (.A(\manchester_baby_instance.ram_data_i_27 ),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__or2_1 _0994_ (.A(_0385_),
    .B(_0409_),
    .X(_0469_));
 sky130_fd_sc_hd__a311o_1 _0995_ (.A1(_0383_),
    .A2(_0469_),
    .A3(_0411_),
    .B1(_0418_),
    .C1(_0410_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _0996_ (.A(_0416_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__xnor2_1 _0997_ (.A(_0415_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__a32o_1 _0998_ (.A1(_0195_),
    .A2(_0441_),
    .A3(_0468_),
    .B1(_0472_),
    .B2(_0106_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(\manchester_baby_instance.ram_data_o_27 ),
    .A1(_0473_),
    .S(_0446_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(_0474_),
    .X(_0058_));
 sky130_fd_sc_hd__o211ai_1 _1001_ (.A1(_0469_),
    .A2(_0412_),
    .B1(_0418_),
    .C1(_0421_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B(_0440_),
    .Y(_0476_));
 sky130_fd_sc_hd__and3_1 _1003_ (.A(_0194_),
    .B(_0467_),
    .C(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__a31o_1 _1004_ (.A1(_0204_),
    .A2(_0470_),
    .A3(_0475_),
    .B1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1005_ (.A0(\manchester_baby_instance.ram_data_o_26 ),
    .A1(_0478_),
    .S(_0446_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_1 _1006_ (.A(_0479_),
    .X(_0057_));
 sky130_fd_sc_hd__or2_1 _1007_ (.A(\manchester_baby_instance.ram_data_i_23 ),
    .B(_0439_),
    .X(_0480_));
 sky130_fd_sc_hd__or2_1 _1008_ (.A(\manchester_baby_instance.ram_data_i_24 ),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(\manchester_baby_instance.ram_data_i_25 ),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_1 _1010_ (.A(_0383_),
    .B(_0469_),
    .Y(_0483_));
 sky130_fd_sc_hd__xnor2_1 _1011_ (.A(_0412_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__a32o_1 _1012_ (.A1(_0195_),
    .A2(_0440_),
    .A3(_0482_),
    .B1(_0484_),
    .B2(_0106_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(\manchester_baby_instance.ram_data_o_25 ),
    .A1(_0485_),
    .S(_0446_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _1014_ (.A(_0486_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(_0385_),
    .B(_0409_),
    .Y(_0487_));
 sky130_fd_sc_hd__nand2_1 _1016_ (.A(\manchester_baby_instance.ram_data_i_24 ),
    .B(_0480_),
    .Y(_0488_));
 sky130_fd_sc_hd__and3_1 _1017_ (.A(_0194_),
    .B(_0481_),
    .C(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__a31o_1 _1018_ (.A1(_0204_),
    .A2(_0469_),
    .A3(_0487_),
    .B1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(\manchester_baby_instance.ram_data_o_24 ),
    .A1(_0490_),
    .S(_0446_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(_0491_),
    .X(_0055_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(_0173_),
    .B(_0400_),
    .Y(_0492_));
 sky130_fd_sc_hd__o21a_1 _1022_ (.A1(_0405_),
    .A2(_0492_),
    .B1(_0389_),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a311o_1 _1024_ (.A1(_0387_),
    .A2(_0401_),
    .A3(_0494_),
    .B1(_0393_),
    .C1(_0386_),
    .X(_0495_));
 sky130_fd_sc_hd__a21oi_1 _1025_ (.A1(_0392_),
    .A2(_0495_),
    .B1(_0396_),
    .Y(_0496_));
 sky130_fd_sc_hd__a31o_1 _1026_ (.A1(_0392_),
    .A2(_0396_),
    .A3(_0495_),
    .B1(_0261_),
    .X(_0497_));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(_0195_),
    .B(_0480_),
    .Y(_0498_));
 sky130_fd_sc_hd__a21o_1 _1028_ (.A1(\manchester_baby_instance.ram_data_i_23 ),
    .A2(_0439_),
    .B1(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__o21ai_1 _1029_ (.A1(_0496_),
    .A2(_0497_),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\manchester_baby_instance.ram_data_o_23 ),
    .A1(_0500_),
    .S(_0446_),
    .X(_0501_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0501_),
    .X(_0054_));
 sky130_fd_sc_hd__a31oi_1 _1032_ (.A1(_0387_),
    .A2(_0401_),
    .A3(_0494_),
    .B1(_0386_),
    .Y(_0502_));
 sky130_fd_sc_hd__or2b_1 _1033_ (.A(_0502_),
    .B_N(_0393_),
    .X(_0503_));
 sky130_fd_sc_hd__or2_1 _1034_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B(_0438_),
    .X(_0504_));
 sky130_fd_sc_hd__or2_1 _1035_ (.A(\manchester_baby_instance.ram_data_i_21 ),
    .B(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_1 _1036_ (.A(\manchester_baby_instance.ram_data_i_22 ),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__and3_1 _1037_ (.A(_0194_),
    .B(_0439_),
    .C(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a31o_1 _1038_ (.A1(_0204_),
    .A2(_0495_),
    .A3(_0503_),
    .B1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(\manchester_baby_instance.ram_data_o_22 ),
    .A1(_0508_),
    .S(_0446_),
    .X(_0509_));
 sky130_fd_sc_hd__clkbuf_1 _1040_ (.A(_0509_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _1041_ (.A(\manchester_baby_instance.ram_data_i_21 ),
    .B(_0504_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1042_ (.A(_0401_),
    .B(_0494_),
    .Y(_0511_));
 sky130_fd_sc_hd__xor2_1 _1043_ (.A(_0388_),
    .B(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a32o_1 _1044_ (.A1(_0195_),
    .A2(_0505_),
    .A3(_0510_),
    .B1(_0512_),
    .B2(_0106_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _1045_ (.A0(\manchester_baby_instance.ram_data_o_21 ),
    .A1(_0513_),
    .S(_0198_),
    .X(_0514_));
 sky130_fd_sc_hd__clkbuf_1 _1046_ (.A(_0514_),
    .X(_0052_));
 sky130_fd_sc_hd__or3_1 _1047_ (.A(_0405_),
    .B(_0389_),
    .C(_0492_),
    .X(_0515_));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B(_0438_),
    .Y(_0516_));
 sky130_fd_sc_hd__and3_1 _1049_ (.A(_0194_),
    .B(_0504_),
    .C(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__a31o_1 _1050_ (.A1(_0204_),
    .A2(_0494_),
    .A3(_0515_),
    .B1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _1051_ (.A0(\manchester_baby_instance.ram_data_o_20 ),
    .A1(_0518_),
    .S(_0198_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_1 _1052_ (.A(_0519_),
    .X(_0051_));
 sky130_fd_sc_hd__o31ai_1 _1053_ (.A1(\manchester_baby_instance.ram_data_i_17 ),
    .A2(\manchester_baby_instance.ram_data_i_18 ),
    .A3(_0191_),
    .B1(\manchester_baby_instance.ram_data_i_19 ),
    .Y(_0520_));
 sky130_fd_sc_hd__and2b_1 _1054_ (.A_N(_0403_),
    .B(_0180_),
    .X(_0521_));
 sky130_fd_sc_hd__xnor2_1 _1055_ (.A(_0398_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__a32o_1 _1056_ (.A1(_0195_),
    .A2(_0438_),
    .A3(_0520_),
    .B1(_0522_),
    .B2(_0106_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _1057_ (.A0(\manchester_baby_instance.ram_data_o_19 ),
    .A1(_0523_),
    .S(_0198_),
    .X(_0524_));
 sky130_fd_sc_hd__clkbuf_1 _1058_ (.A(_0524_),
    .X(_0050_));
 sky130_fd_sc_hd__nand2_1 _1059_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_4 _1060_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand4b_4 _1061_ (.A_N(_0104_),
    .B(_0101_),
    .C(_0331_),
    .D(_0526_),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0556_),
    .Y(net8));
 sky130_fd_sc_hd__clkbuf_2 _1063_ (.A(_0104_),
    .X(_0527_));
 sky130_fd_sc_hd__buf_4 _1064_ (.A(_0101_),
    .X(_0528_));
 sky130_fd_sc_hd__buf_4 _1065_ (.A(_0331_),
    .X(_0529_));
 sky130_fd_sc_hd__buf_4 _1066_ (.A(_0526_),
    .X(_0530_));
 sky130_fd_sc_hd__nand4b_2 _1067_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0557_));
 sky130_fd_sc_hd__nand4b_2 _1068_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand4b_2 _1069_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand4b_2 _1070_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand4b_2 _1071_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand4b_2 _1072_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand4b_2 _1073_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand4b_2 _1074_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand4b_2 _1075_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand4b_2 _1076_ (.A_N(_0527_),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .Y(_0566_));
 sky130_fd_sc_hd__clkbuf_2 _1077_ (.A(_0104_),
    .X(_0531_));
 sky130_fd_sc_hd__buf_4 _1078_ (.A(_0101_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_4 _1079_ (.A(_0331_),
    .X(_0533_));
 sky130_fd_sc_hd__buf_4 _1080_ (.A(_0526_),
    .X(_0534_));
 sky130_fd_sc_hd__nand4b_2 _1081_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand4b_2 _1082_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0568_));
 sky130_fd_sc_hd__nand4b_2 _1083_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand4b_2 _1084_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand4b_2 _1085_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand4b_2 _1086_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand4b_2 _1087_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand4b_2 _1088_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand4b_2 _1089_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand4b_2 _1090_ (.A_N(_0531_),
    .B(_0532_),
    .C(_0533_),
    .D(_0534_),
    .Y(_0576_));
 sky130_fd_sc_hd__clkbuf_2 _1091_ (.A(_0104_),
    .X(_0535_));
 sky130_fd_sc_hd__buf_4 _1092_ (.A(_0101_),
    .X(_0536_));
 sky130_fd_sc_hd__buf_4 _1093_ (.A(_0331_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_4 _1094_ (.A(_0526_),
    .X(_0538_));
 sky130_fd_sc_hd__nand4b_2 _1095_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand4b_2 _1096_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand4b_2 _1097_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand4b_2 _1098_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand4b_2 _1099_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand4b_2 _1100_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0582_));
 sky130_fd_sc_hd__nand4b_2 _1101_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand4b_2 _1102_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand4b_2 _1103_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand4b_2 _1104_ (.A_N(_0535_),
    .B(_0536_),
    .C(_0537_),
    .D(_0538_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand4b_2 _1105_ (.A_N(_0104_),
    .B(_0101_),
    .C(_0331_),
    .D(_0526_),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _1106_ (.A(net16),
    .B(net19),
    .X(_0539_));
 sky130_fd_sc_hd__nor2_1 _1107_ (.A(net17),
    .B(_0539_),
    .Y(\manchester_baby_instance.BASE_0.s_tickNext ));
 sky130_fd_sc_hd__and2b_1 _1108_ (.A_N(_0102_),
    .B(_0525_),
    .X(_0540_));
 sky130_fd_sc_hd__clkbuf_1 _1109_ (.A(_0540_),
    .X(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ));
 sky130_fd_sc_hd__and2_1 _1110_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0525_),
    .X(_0541_));
 sky130_fd_sc_hd__or2_1 _1111_ (.A(_0526_),
    .B(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__clkbuf_1 _1112_ (.A(_0542_),
    .X(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ));
 sky130_fd_sc_hd__and2b_1 _1113_ (.A_N(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .B(net15),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1114_ (.A(_0543_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _1115_ (.A_N(net9),
    .B(net2),
    .X(_0544_));
 sky130_fd_sc_hd__buf_1 _1116_ (.A(_0544_),
    .X(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ));
 sky130_fd_sc_hd__nor3_2 _1117_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .Y(_0545_));
 sky130_fd_sc_hd__a22o_1 _1118_ (.A1(_0103_),
    .A2(_0312_),
    .B1(_0314_),
    .B2(_0526_),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _1119_ (.A1(_0337_),
    .A2(_0545_),
    .B1(_0546_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net3));
 sky130_fd_sc_hd__a22o_1 _1120_ (.A1(_0319_),
    .A2(_0545_),
    .B1(_0546_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net4));
 sky130_fd_sc_hd__a22o_1 _1121_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0545_),
    .B1(_0546_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net5));
 sky130_fd_sc_hd__a22o_1 _1122_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0545_),
    .B1(_0546_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net6));
 sky130_fd_sc_hd__a22o_1 _1123_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0545_),
    .B1(_0546_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net7));
 sky130_fd_sc_hd__buf_4 _1124_ (.A(net1),
    .X(_0547_));
 sky130_fd_sc_hd__buf_4 _1125_ (.A(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(_0548_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1127_ (.A(_0548_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(_0548_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1129_ (.A(_0548_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1130_ (.A(_0548_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(_0548_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(_0548_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(_0548_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1134_ (.A(_0548_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(_0548_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_4 _1136_ (.A(net1),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _1137_ (.A(_0549_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1138_ (.A(_0549_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1139_ (.A(_0549_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(_0549_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1141_ (.A(_0549_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1142_ (.A(_0549_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1143_ (.A(_0549_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1144_ (.A(_0549_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(_0549_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(_0549_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_4 _1147_ (.A(net1),
    .X(_0550_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(_0550_),
    .Y(_0021_));
 sky130_fd_sc_hd__or2b_1 _1149_ (.A(net20),
    .B_N(\manchester_baby_instance.BASE_0.s_tickReg ),
    .X(_0551_));
 sky130_fd_sc_hd__xnor2_1 _1150_ (.A(net15),
    .B(net21),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(_0550_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1152_ (.A(_0550_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1153_ (.A(_0550_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1154_ (.A(_0550_),
    .Y(_0025_));
 sky130_fd_sc_hd__and2b_1 _1155_ (.A_N(net24),
    .B(net20),
    .X(_0552_));
 sky130_fd_sc_hd__clkbuf_1 _1156_ (.A(_0552_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(net16),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _1158_ (.A(net16),
    .B(net19),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2_1 _1159_ (.A(_0539_),
    .B(_0553_),
    .Y(_0075_));
 sky130_fd_sc_hd__and2_1 _1160_ (.A(net17),
    .B(_0539_),
    .X(_0554_));
 sky130_fd_sc_hd__clkbuf_1 _1161_ (.A(_0554_),
    .X(_0076_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(_0550_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1163_ (.A(_0550_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(_0550_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(_0550_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(_0550_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_4 _1167_ (.A(net1),
    .X(_0555_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(_0555_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(_0555_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(_0555_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(_0555_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1172_ (.A(_0555_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(_0555_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(_0555_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1175_ (.A(_0555_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1176_ (.A(_0555_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1177_ (.A(_0555_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1178_ (.A(_0547_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(_0547_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(_0547_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1181_ (.A(_0547_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(_0547_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(_0547_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(_0547_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(_0547_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1186_ (.A(_0547_),
    .Y(_0049_));
 sky130_fd_sc_hd__dfrtp_2 _1187_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0050_),
    .RESET_B(_0001_),
    .Q(\manchester_baby_instance.ram_data_o_19 ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0051_),
    .RESET_B(_0002_),
    .Q(\manchester_baby_instance.ram_data_o_20 ));
 sky130_fd_sc_hd__dfrtp_1 _1189_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0052_),
    .RESET_B(_0003_),
    .Q(\manchester_baby_instance.ram_data_o_21 ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0053_),
    .RESET_B(_0004_),
    .Q(\manchester_baby_instance.ram_data_o_22 ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0054_),
    .RESET_B(_0005_),
    .Q(\manchester_baby_instance.ram_data_o_23 ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0055_),
    .RESET_B(_0006_),
    .Q(\manchester_baby_instance.ram_data_o_24 ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0056_),
    .RESET_B(_0007_),
    .Q(\manchester_baby_instance.ram_data_o_25 ));
 sky130_fd_sc_hd__dfrtp_1 _1194_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0057_),
    .RESET_B(_0008_),
    .Q(\manchester_baby_instance.ram_data_o_26 ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0058_),
    .RESET_B(_0009_),
    .Q(\manchester_baby_instance.ram_data_o_27 ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0059_),
    .RESET_B(_0010_),
    .Q(\manchester_baby_instance.ram_data_o_28 ));
 sky130_fd_sc_hd__dfrtp_1 _1197_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0060_),
    .RESET_B(_0011_),
    .Q(\manchester_baby_instance.ram_data_o_29 ));
 sky130_fd_sc_hd__dfrtp_1 _1198_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0061_),
    .RESET_B(_0012_),
    .Q(\manchester_baby_instance.ram_data_o_30 ));
 sky130_fd_sc_hd__dfrtp_4 _1199_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0062_),
    .RESET_B(_0013_),
    .Q(\manchester_baby_instance.ram_data_o_31 ));
 sky130_fd_sc_hd__dfrtp_1 _1200_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0063_),
    .RESET_B(_0014_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1201_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0064_),
    .RESET_B(_0015_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1202_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0065_),
    .RESET_B(_0016_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1203_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0066_),
    .RESET_B(_0017_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1204_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0067_),
    .RESET_B(_0018_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1205_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0068_),
    .RESET_B(_0019_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1206_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0069_),
    .RESET_B(_0020_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1207_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0070_),
    .RESET_B(_0021_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0071_),
    .Q(\manchester_baby_instance.BASE_1.s_derivedClock ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .RESET_B(_0022_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ),
    .RESET_B(_0023_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1211_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ),
    .RESET_B(_0024_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(clknet_2_3__leaf_clock),
    .D(net23),
    .RESET_B(_0025_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(clknet_2_3__leaf_clock),
    .D(net15),
    .Q(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0073_),
    .Q(\manchester_baby_instance.BASE_1.s_counterValue ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0074_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0075_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0076_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(clknet_2_3__leaf_clock),
    .D(net18),
    .Q(\manchester_baby_instance.BASE_0.s_tickReg ));
 sky130_fd_sc_hd__dlxtn_2 _1219_ (.D(ram_data_io[0]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_0 ));
 sky130_fd_sc_hd__dlxtn_2 _1220_ (.D(ram_data_io[1]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_1 ));
 sky130_fd_sc_hd__dlxtn_1 _1221_ (.D(ram_data_io[2]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_2 ));
 sky130_fd_sc_hd__dlxtn_2 _1222_ (.D(ram_data_io[3]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_3 ));
 sky130_fd_sc_hd__dlxtn_2 _1223_ (.D(ram_data_io[4]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_4 ));
 sky130_fd_sc_hd__dlxtn_1 _1224_ (.D(ram_data_io[5]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_5 ));
 sky130_fd_sc_hd__dlxtn_1 _1225_ (.D(ram_data_io[6]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_6 ));
 sky130_fd_sc_hd__dlxtn_1 _1226_ (.D(ram_data_io[7]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_7 ));
 sky130_fd_sc_hd__dlxtn_1 _1227_ (.D(ram_data_io[8]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_8 ));
 sky130_fd_sc_hd__dlxtn_1 _1228_ (.D(ram_data_io[9]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_9 ));
 sky130_fd_sc_hd__dlxtn_1 _1229_ (.D(ram_data_io[10]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_10 ));
 sky130_fd_sc_hd__dlxtn_1 _1230_ (.D(ram_data_io[11]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_11 ));
 sky130_fd_sc_hd__dlxtn_1 _1231_ (.D(ram_data_io[12]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_12 ));
 sky130_fd_sc_hd__dlxtn_1 _1232_ (.D(ram_data_io[13]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_13 ));
 sky130_fd_sc_hd__dlxtn_1 _1233_ (.D(ram_data_io[14]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_14 ));
 sky130_fd_sc_hd__dlxtn_1 _1234_ (.D(ram_data_io[15]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_15 ));
 sky130_fd_sc_hd__dlxtn_1 _1235_ (.D(ram_data_io[16]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_16 ));
 sky130_fd_sc_hd__dlxtn_1 _1236_ (.D(ram_data_io[17]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_17 ));
 sky130_fd_sc_hd__dlxtn_1 _1237_ (.D(ram_data_io[18]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_18 ));
 sky130_fd_sc_hd__dlxtn_1 _1238_ (.D(ram_data_io[19]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_19 ));
 sky130_fd_sc_hd__dlxtn_1 _1239_ (.D(ram_data_io[20]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_20 ));
 sky130_fd_sc_hd__dlxtn_1 _1240_ (.D(ram_data_io[21]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_21 ));
 sky130_fd_sc_hd__dlxtn_1 _1241_ (.D(ram_data_io[22]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_22 ));
 sky130_fd_sc_hd__dlxtn_1 _1242_ (.D(ram_data_io[23]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_23 ));
 sky130_fd_sc_hd__dlxtn_1 _1243_ (.D(ram_data_io[24]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_24 ));
 sky130_fd_sc_hd__dlxtn_1 _1244_ (.D(ram_data_io[25]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_25 ));
 sky130_fd_sc_hd__dlxtn_1 _1245_ (.D(ram_data_io[26]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_26 ));
 sky130_fd_sc_hd__dlxtn_1 _1246_ (.D(ram_data_io[27]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_27 ));
 sky130_fd_sc_hd__dlxtn_1 _1247_ (.D(ram_data_io[28]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_28 ));
 sky130_fd_sc_hd__dlxtn_1 _1248_ (.D(ram_data_io[29]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_29 ));
 sky130_fd_sc_hd__dlxtn_1 _1249_ (.D(ram_data_io[30]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_30 ));
 sky130_fd_sc_hd__dlxtn_1 _1250_ (.D(ram_data_io[31]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_31 ));
 sky130_fd_sc_hd__dfxtp_1 _1251_ (.CLK(clknet_2_3__leaf_clock),
    .D(net14),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_1 _1252_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0000_),
    .Q(\manchester_baby_instance.CIRCUIT_0.Acc.tick ));
 sky130_fd_sc_hd__dfrtp_1 _1253_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0077_),
    .RESET_B(_0026_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1254_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0078_),
    .RESET_B(_0027_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1255_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0079_),
    .RESET_B(_0028_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1256_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0080_),
    .RESET_B(_0029_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1257_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0081_),
    .RESET_B(_0030_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1258_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0082_),
    .RESET_B(_0031_),
    .Q(\manchester_baby_instance.ram_data_o_0 ));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0083_),
    .RESET_B(_0032_),
    .Q(\manchester_baby_instance.ram_data_o_1 ));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0084_),
    .RESET_B(_0033_),
    .Q(\manchester_baby_instance.ram_data_o_2 ));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0085_),
    .RESET_B(_0034_),
    .Q(\manchester_baby_instance.ram_data_o_3 ));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0086_),
    .RESET_B(_0035_),
    .Q(\manchester_baby_instance.ram_data_o_4 ));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0087_),
    .RESET_B(_0036_),
    .Q(\manchester_baby_instance.ram_data_o_5 ));
 sky130_fd_sc_hd__dfrtp_2 _1264_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0088_),
    .RESET_B(_0037_),
    .Q(\manchester_baby_instance.ram_data_o_6 ));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0089_),
    .RESET_B(_0038_),
    .Q(\manchester_baby_instance.ram_data_o_7 ));
 sky130_fd_sc_hd__dfrtp_1 _1266_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0090_),
    .RESET_B(_0039_),
    .Q(\manchester_baby_instance.ram_data_o_8 ));
 sky130_fd_sc_hd__dfrtp_1 _1267_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0091_),
    .RESET_B(_0040_),
    .Q(\manchester_baby_instance.ram_data_o_9 ));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0092_),
    .RESET_B(_0041_),
    .Q(\manchester_baby_instance.ram_data_o_10 ));
 sky130_fd_sc_hd__dfrtp_2 _1269_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0093_),
    .RESET_B(_0042_),
    .Q(\manchester_baby_instance.ram_data_o_11 ));
 sky130_fd_sc_hd__dfrtp_2 _1270_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0094_),
    .RESET_B(_0043_),
    .Q(\manchester_baby_instance.ram_data_o_12 ));
 sky130_fd_sc_hd__dfrtp_1 _1271_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0095_),
    .RESET_B(_0044_),
    .Q(\manchester_baby_instance.ram_data_o_13 ));
 sky130_fd_sc_hd__dfrtp_1 _1272_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0096_),
    .RESET_B(_0045_),
    .Q(\manchester_baby_instance.ram_data_o_14 ));
 sky130_fd_sc_hd__dfrtp_1 _1273_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0097_),
    .RESET_B(_0046_),
    .Q(\manchester_baby_instance.ram_data_o_15 ));
 sky130_fd_sc_hd__dfrtp_2 _1274_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0098_),
    .RESET_B(_0047_),
    .Q(\manchester_baby_instance.ram_data_o_16 ));
 sky130_fd_sc_hd__dfrtp_1 _1275_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0099_),
    .RESET_B(_0048_),
    .Q(\manchester_baby_instance.ram_data_o_17 ));
 sky130_fd_sc_hd__dfrtp_1 _1276_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0100_),
    .RESET_B(_0049_),
    .Q(\manchester_baby_instance.ram_data_o_18 ));
 sky130_fd_sc_hd__ebufn_8 _1277_ (.A(\manchester_baby_instance.ram_data_o_0 ),
    .TE_B(_0556_),
    .Z(ram_data_io[0]));
 sky130_fd_sc_hd__ebufn_8 _1278_ (.A(\manchester_baby_instance.ram_data_o_1 ),
    .TE_B(_0557_),
    .Z(ram_data_io[1]));
 sky130_fd_sc_hd__ebufn_8 _1279_ (.A(\manchester_baby_instance.ram_data_o_2 ),
    .TE_B(_0558_),
    .Z(ram_data_io[2]));
 sky130_fd_sc_hd__ebufn_8 _1280_ (.A(\manchester_baby_instance.ram_data_o_3 ),
    .TE_B(_0559_),
    .Z(ram_data_io[3]));
 sky130_fd_sc_hd__ebufn_8 _1281_ (.A(\manchester_baby_instance.ram_data_o_4 ),
    .TE_B(_0560_),
    .Z(ram_data_io[4]));
 sky130_fd_sc_hd__ebufn_8 _1282_ (.A(\manchester_baby_instance.ram_data_o_5 ),
    .TE_B(_0561_),
    .Z(ram_data_io[5]));
 sky130_fd_sc_hd__ebufn_8 _1283_ (.A(\manchester_baby_instance.ram_data_o_6 ),
    .TE_B(_0562_),
    .Z(ram_data_io[6]));
 sky130_fd_sc_hd__ebufn_8 _1284_ (.A(\manchester_baby_instance.ram_data_o_7 ),
    .TE_B(_0563_),
    .Z(ram_data_io[7]));
 sky130_fd_sc_hd__ebufn_8 _1285_ (.A(\manchester_baby_instance.ram_data_o_8 ),
    .TE_B(_0564_),
    .Z(ram_data_io[8]));
 sky130_fd_sc_hd__ebufn_8 _1286_ (.A(\manchester_baby_instance.ram_data_o_9 ),
    .TE_B(_0565_),
    .Z(ram_data_io[9]));
 sky130_fd_sc_hd__ebufn_8 _1287_ (.A(\manchester_baby_instance.ram_data_o_10 ),
    .TE_B(_0566_),
    .Z(ram_data_io[10]));
 sky130_fd_sc_hd__ebufn_8 _1288_ (.A(\manchester_baby_instance.ram_data_o_11 ),
    .TE_B(_0567_),
    .Z(ram_data_io[11]));
 sky130_fd_sc_hd__ebufn_8 _1289_ (.A(\manchester_baby_instance.ram_data_o_12 ),
    .TE_B(_0568_),
    .Z(ram_data_io[12]));
 sky130_fd_sc_hd__ebufn_8 _1290_ (.A(\manchester_baby_instance.ram_data_o_13 ),
    .TE_B(_0569_),
    .Z(ram_data_io[13]));
 sky130_fd_sc_hd__ebufn_8 _1291_ (.A(\manchester_baby_instance.ram_data_o_14 ),
    .TE_B(_0570_),
    .Z(ram_data_io[14]));
 sky130_fd_sc_hd__ebufn_8 _1292_ (.A(\manchester_baby_instance.ram_data_o_15 ),
    .TE_B(_0571_),
    .Z(ram_data_io[15]));
 sky130_fd_sc_hd__ebufn_8 _1293_ (.A(\manchester_baby_instance.ram_data_o_16 ),
    .TE_B(_0572_),
    .Z(ram_data_io[16]));
 sky130_fd_sc_hd__ebufn_8 _1294_ (.A(\manchester_baby_instance.ram_data_o_17 ),
    .TE_B(_0573_),
    .Z(ram_data_io[17]));
 sky130_fd_sc_hd__ebufn_8 _1295_ (.A(\manchester_baby_instance.ram_data_o_18 ),
    .TE_B(_0574_),
    .Z(ram_data_io[18]));
 sky130_fd_sc_hd__ebufn_8 _1296_ (.A(\manchester_baby_instance.ram_data_o_19 ),
    .TE_B(_0575_),
    .Z(ram_data_io[19]));
 sky130_fd_sc_hd__ebufn_8 _1297_ (.A(\manchester_baby_instance.ram_data_o_20 ),
    .TE_B(_0576_),
    .Z(ram_data_io[20]));
 sky130_fd_sc_hd__ebufn_8 _1298_ (.A(\manchester_baby_instance.ram_data_o_21 ),
    .TE_B(_0577_),
    .Z(ram_data_io[21]));
 sky130_fd_sc_hd__ebufn_8 _1299_ (.A(\manchester_baby_instance.ram_data_o_22 ),
    .TE_B(_0578_),
    .Z(ram_data_io[22]));
 sky130_fd_sc_hd__ebufn_8 _1300_ (.A(\manchester_baby_instance.ram_data_o_23 ),
    .TE_B(_0579_),
    .Z(ram_data_io[23]));
 sky130_fd_sc_hd__ebufn_8 _1301_ (.A(\manchester_baby_instance.ram_data_o_24 ),
    .TE_B(_0580_),
    .Z(ram_data_io[24]));
 sky130_fd_sc_hd__ebufn_8 _1302_ (.A(\manchester_baby_instance.ram_data_o_25 ),
    .TE_B(_0581_),
    .Z(ram_data_io[25]));
 sky130_fd_sc_hd__ebufn_8 _1303_ (.A(\manchester_baby_instance.ram_data_o_26 ),
    .TE_B(_0582_),
    .Z(ram_data_io[26]));
 sky130_fd_sc_hd__ebufn_8 _1304_ (.A(\manchester_baby_instance.ram_data_o_27 ),
    .TE_B(_0583_),
    .Z(ram_data_io[27]));
 sky130_fd_sc_hd__ebufn_8 _1305_ (.A(\manchester_baby_instance.ram_data_o_28 ),
    .TE_B(_0584_),
    .Z(ram_data_io[28]));
 sky130_fd_sc_hd__ebufn_8 _1306_ (.A(\manchester_baby_instance.ram_data_o_29 ),
    .TE_B(_0585_),
    .Z(ram_data_io[29]));
 sky130_fd_sc_hd__ebufn_8 _1307_ (.A(\manchester_baby_instance.ram_data_o_30 ),
    .TE_B(_0586_),
    .Z(ram_data_io[30]));
 sky130_fd_sc_hd__ebufn_8 _1308_ (.A(\manchester_baby_instance.ram_data_o_31 ),
    .TE_B(_0587_),
    .Z(ram_data_io[31]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clock (.A(clock),
    .X(clknet_0_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clock (.A(clknet_0_clock),
    .X(clknet_2_0__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clock (.A(clknet_0_clock),
    .X(clknet_2_1__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clock (.A(clknet_0_clock),
    .X(clknet_2_2__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clock (.A(clknet_0_clock),
    .X(clknet_2_3__leaf_clock));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(net13),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 fanout13 (.A(net8),
    .X(net13));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .X(net14));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0072_),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\manchester_baby_instance.BASE_0.s_tickReg ),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\manchester_baby_instance.ram_data_o_0 ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .X(net15));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .X(net16));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\manchester_baby_instance.BASE_0.s_tickNext ),
    .X(net18));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\manchester_baby_instance.BASE_1.s_counterValue ),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0551_),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net9),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(reset_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 output2 (.A(net2),
    .X(logisim_clock_tree_0_out));
 sky130_fd_sc_hd__clkbuf_4 output3 (.A(net3),
    .X(ram_addr_o[0]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(ram_addr_o[1]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(ram_addr_o[2]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(ram_addr_o[3]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(ram_addr_o[4]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net13),
    .X(ram_rw_en_o));
 sky130_fd_sc_hd__clkbuf_4 output9 (.A(net9),
    .X(stop_lamp_o));
endmodule

