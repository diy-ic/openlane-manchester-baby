magic
tech sky130A
magscale 1 2
timestamp 1702734622
<< viali >>
rect 12449 29257 12483 29291
rect 14381 29257 14415 29291
rect 15761 29257 15795 29291
rect 19441 29257 19475 29291
rect 19993 29257 20027 29291
rect 20913 29257 20947 29291
rect 22201 29257 22235 29291
rect 15025 29189 15059 29223
rect 12725 29121 12759 29155
rect 13185 29121 13219 29155
rect 14657 29121 14691 29155
rect 15669 29121 15703 29155
rect 19349 29121 19383 29155
rect 19901 29121 19935 29155
rect 20821 29121 20855 29155
rect 22109 29121 22143 29155
rect 13001 28985 13035 29019
rect 15209 28985 15243 29019
rect 21189 25857 21223 25891
rect 21281 25653 21315 25687
rect 18797 25449 18831 25483
rect 14565 25313 14599 25347
rect 14841 25313 14875 25347
rect 20177 25313 20211 25347
rect 26433 25313 26467 25347
rect 14473 25245 14507 25279
rect 15853 25245 15887 25279
rect 15945 25245 15979 25279
rect 18889 25245 18923 25279
rect 19349 25245 19383 25279
rect 24133 25245 24167 25279
rect 24409 25245 24443 25279
rect 16221 25177 16255 25211
rect 17969 25177 18003 25211
rect 20453 25177 20487 25211
rect 22201 25177 22235 25211
rect 23857 25177 23891 25211
rect 24685 25177 24719 25211
rect 15761 25109 15795 25143
rect 18429 25109 18463 25143
rect 19441 25109 19475 25143
rect 22385 25109 22419 25143
rect 17233 24905 17267 24939
rect 20269 24905 20303 24939
rect 22017 24905 22051 24939
rect 22937 24905 22971 24939
rect 24409 24905 24443 24939
rect 25237 24905 25271 24939
rect 14749 24837 14783 24871
rect 17325 24769 17359 24803
rect 18153 24769 18187 24803
rect 18337 24769 18371 24803
rect 20453 24769 20487 24803
rect 20545 24769 20579 24803
rect 20637 24769 20671 24803
rect 20821 24769 20855 24803
rect 22201 24769 22235 24803
rect 22293 24769 22327 24803
rect 22385 24769 22419 24803
rect 22569 24769 22603 24803
rect 22845 24769 22879 24803
rect 23857 24769 23891 24803
rect 24041 24769 24075 24803
rect 24133 24769 24167 24803
rect 24225 24769 24259 24803
rect 25145 24769 25179 24803
rect 12357 24701 12391 24735
rect 12633 24701 12667 24735
rect 14381 24701 14415 24735
rect 14473 24701 14507 24735
rect 16497 24701 16531 24735
rect 18429 24701 18463 24735
rect 18705 24701 18739 24735
rect 23121 24701 23155 24735
rect 23673 24701 23707 24735
rect 17969 24565 18003 24599
rect 20177 24565 20211 24599
rect 13185 24361 13219 24395
rect 14197 24361 14231 24395
rect 16129 24361 16163 24395
rect 17693 24361 17727 24395
rect 19073 24361 19107 24395
rect 20269 24361 20303 24395
rect 20545 24361 20579 24395
rect 21189 24361 21223 24395
rect 21833 24361 21867 24395
rect 22063 24361 22097 24395
rect 22661 24361 22695 24395
rect 13093 24293 13127 24327
rect 18061 24293 18095 24327
rect 23397 24293 23431 24327
rect 15393 24225 15427 24259
rect 17785 24225 17819 24259
rect 20729 24225 20763 24259
rect 20821 24225 20855 24259
rect 20914 24225 20948 24259
rect 21925 24225 21959 24259
rect 12909 24157 12943 24191
rect 13369 24157 13403 24191
rect 14289 24157 14323 24191
rect 14473 24157 14507 24191
rect 14841 24157 14875 24191
rect 14933 24157 14967 24191
rect 16037 24157 16071 24191
rect 17049 24157 17083 24191
rect 17325 24157 17359 24191
rect 17417 24157 17451 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 18705 24157 18739 24191
rect 18889 24157 18923 24191
rect 20453 24157 20487 24191
rect 21006 24157 21040 24191
rect 21741 24157 21775 24191
rect 22201 24157 22235 24191
rect 22845 24157 22879 24191
rect 23121 24157 23155 24191
rect 23397 24157 23431 24191
rect 23673 24157 23707 24191
rect 24593 24157 24627 24191
rect 24869 24157 24903 24191
rect 25145 24157 25179 24191
rect 15025 24089 15059 24123
rect 15209 24089 15243 24123
rect 18797 24089 18831 24123
rect 21373 24089 21407 24123
rect 21557 24089 21591 24123
rect 25421 24089 25455 24123
rect 14749 24021 14783 24055
rect 17509 24021 17543 24055
rect 23029 24021 23063 24055
rect 23581 24021 23615 24055
rect 24501 24021 24535 24055
rect 25053 24021 25087 24055
rect 26893 24021 26927 24055
rect 13001 23817 13035 23851
rect 15209 23817 15243 23851
rect 15393 23817 15427 23851
rect 17049 23817 17083 23851
rect 18153 23817 18187 23851
rect 19441 23817 19475 23851
rect 20913 23817 20947 23851
rect 22033 23817 22067 23851
rect 24961 23817 24995 23851
rect 25329 23817 25363 23851
rect 26065 23817 26099 23851
rect 13461 23749 13495 23783
rect 18797 23749 18831 23783
rect 19717 23749 19751 23783
rect 21833 23749 21867 23783
rect 1501 23681 1535 23715
rect 11529 23681 11563 23715
rect 11796 23681 11830 23715
rect 14841 23681 14875 23715
rect 17785 23681 17819 23715
rect 17969 23681 18003 23715
rect 18521 23681 18555 23715
rect 18613 23681 18647 23715
rect 18981 23681 19015 23715
rect 19165 23681 19199 23715
rect 19901 23681 19935 23715
rect 20821 23681 20855 23715
rect 21005 23681 21039 23715
rect 23489 23681 23523 23715
rect 24593 23681 24627 23715
rect 24777 23681 24811 23715
rect 24869 23681 24903 23715
rect 25973 23681 26007 23715
rect 30389 23681 30423 23715
rect 17693 23613 17727 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 19257 23613 19291 23647
rect 19533 23613 19567 23647
rect 23305 23613 23339 23647
rect 23398 23613 23432 23647
rect 23581 23613 23615 23647
rect 23765 23613 23799 23647
rect 23949 23613 23983 23647
rect 24041 23613 24075 23647
rect 24133 23613 24167 23647
rect 24225 23613 24259 23647
rect 25421 23613 25455 23647
rect 25605 23613 25639 23647
rect 1685 23545 1719 23579
rect 12909 23545 12943 23579
rect 13185 23545 13219 23579
rect 16681 23545 16715 23579
rect 22201 23545 22235 23579
rect 30205 23545 30239 23579
rect 15209 23477 15243 23511
rect 17049 23477 17083 23511
rect 17233 23477 17267 23511
rect 22017 23477 22051 23511
rect 23121 23477 23155 23511
rect 24409 23477 24443 23511
rect 12265 23273 12299 23307
rect 15761 23273 15795 23307
rect 23765 23273 23799 23307
rect 25237 23273 25271 23307
rect 11437 23205 11471 23239
rect 16129 23205 16163 23239
rect 22385 23205 22419 23239
rect 10057 23137 10091 23171
rect 11621 23137 11655 23171
rect 14841 23137 14875 23171
rect 15117 23137 15151 23171
rect 15209 23137 15243 23171
rect 16497 23137 16531 23171
rect 19901 23137 19935 23171
rect 20545 23137 20579 23171
rect 22017 23137 22051 23171
rect 23305 23137 23339 23171
rect 12449 23069 12483 23103
rect 16589 23069 16623 23103
rect 16957 23069 16991 23103
rect 17049 23069 17083 23103
rect 17233 23069 17267 23103
rect 19993 23069 20027 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 22201 23069 22235 23103
rect 23581 23069 23615 23103
rect 23673 23069 23707 23103
rect 23857 23069 23891 23103
rect 24041 23069 24075 23103
rect 24593 23069 24627 23103
rect 24741 23069 24775 23103
rect 25099 23069 25133 23103
rect 10302 23001 10336 23035
rect 12716 23001 12750 23035
rect 15326 23001 15360 23035
rect 15761 23001 15795 23035
rect 17417 23001 17451 23035
rect 24869 23001 24903 23035
rect 24961 23001 24995 23035
rect 13829 22933 13863 22967
rect 15485 22933 15519 22967
rect 15577 22933 15611 22967
rect 16865 22933 16899 22967
rect 20361 22933 20395 22967
rect 12817 22729 12851 22763
rect 18521 22729 18555 22763
rect 18889 22729 18923 22763
rect 21189 22729 21223 22763
rect 21557 22729 21591 22763
rect 25881 22729 25915 22763
rect 12265 22661 12299 22695
rect 18429 22661 18463 22695
rect 20821 22661 20855 22695
rect 20913 22661 20947 22695
rect 22385 22661 22419 22695
rect 22937 22661 22971 22695
rect 30205 22661 30239 22695
rect 1685 22593 1719 22627
rect 4813 22593 4847 22627
rect 4997 22593 5031 22627
rect 6745 22593 6779 22627
rect 6929 22593 6963 22627
rect 7757 22593 7791 22627
rect 13001 22593 13035 22627
rect 15301 22593 15335 22627
rect 18337 22593 18371 22627
rect 19073 22593 19107 22627
rect 19165 22593 19199 22627
rect 20545 22593 20579 22627
rect 20693 22593 20727 22627
rect 21010 22593 21044 22627
rect 21281 22593 21315 22627
rect 21373 22593 21407 22627
rect 21661 22599 21695 22633
rect 22109 22593 22143 22627
rect 22293 22593 22327 22627
rect 22477 22593 22511 22627
rect 22595 22593 22629 22627
rect 23029 22593 23063 22627
rect 25421 22593 25455 22627
rect 26249 22593 26283 22627
rect 30481 22593 30515 22627
rect 5181 22525 5215 22559
rect 6837 22525 6871 22559
rect 7573 22525 7607 22559
rect 8309 22525 8343 22559
rect 9965 22525 9999 22559
rect 11621 22525 11655 22559
rect 12725 22525 12759 22559
rect 13829 22525 13863 22559
rect 15025 22525 15059 22559
rect 18797 22525 18831 22559
rect 18889 22525 18923 22559
rect 21465 22525 21499 22559
rect 22753 22525 22787 22559
rect 25513 22525 25547 22559
rect 26157 22525 26191 22559
rect 1501 22457 1535 22491
rect 12541 22457 12575 22491
rect 25789 22457 25823 22491
rect 4905 22389 4939 22423
rect 5733 22389 5767 22423
rect 7021 22389 7055 22423
rect 9413 22389 9447 22423
rect 12173 22389 12207 22423
rect 13277 22389 13311 22423
rect 14749 22389 14783 22423
rect 15025 22389 15059 22423
rect 5181 22185 5215 22219
rect 5641 22185 5675 22219
rect 9229 22185 9263 22219
rect 11621 22185 11655 22219
rect 12436 22185 12470 22219
rect 15761 22185 15795 22219
rect 17417 22185 17451 22219
rect 18153 22185 18187 22219
rect 18613 22185 18647 22219
rect 18797 22185 18831 22219
rect 20453 22185 20487 22219
rect 20637 22185 20671 22219
rect 23673 22185 23707 22219
rect 16405 22117 16439 22151
rect 18337 22117 18371 22151
rect 7665 22049 7699 22083
rect 9413 22049 9447 22083
rect 9505 22049 9539 22083
rect 12173 22049 12207 22083
rect 14749 22049 14783 22083
rect 14958 22049 14992 22083
rect 15485 22049 15519 22083
rect 16497 22049 16531 22083
rect 16773 22049 16807 22083
rect 17785 22049 17819 22083
rect 21281 22049 21315 22083
rect 23121 22049 23155 22083
rect 1685 21981 1719 22015
rect 3801 21981 3835 22015
rect 5825 21981 5859 22015
rect 7481 21981 7515 22015
rect 8769 21981 8803 22015
rect 8953 21981 8987 22015
rect 10241 21981 10275 22015
rect 14289 21981 14323 22015
rect 14473 21981 14507 22015
rect 15393 21981 15427 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 16221 21981 16255 22015
rect 16865 21981 16899 22015
rect 17233 21981 17267 22015
rect 17417 21981 17451 22015
rect 20085 21981 20119 22015
rect 21465 21981 21499 22015
rect 21557 21981 21591 22015
rect 21649 21981 21683 22015
rect 21741 21981 21775 22015
rect 23581 21981 23615 22015
rect 23857 21981 23891 22015
rect 23949 21981 23983 22015
rect 24133 21981 24167 22015
rect 24225 21981 24259 22015
rect 24409 21981 24443 22015
rect 24777 21981 24811 22015
rect 30205 21981 30239 22015
rect 4068 21913 4102 21947
rect 5273 21913 5307 21947
rect 5457 21913 5491 21947
rect 6092 21913 6126 21947
rect 10486 21913 10520 21947
rect 14197 21913 14231 21947
rect 16129 21913 16163 21947
rect 16982 21913 17016 21947
rect 18153 21913 18187 21947
rect 18429 21913 18463 21947
rect 24593 21913 24627 21947
rect 24685 21913 24719 21947
rect 1501 21845 1535 21879
rect 7205 21845 7239 21879
rect 7297 21845 7331 21879
rect 8585 21845 8619 21879
rect 10149 21845 10183 21879
rect 13921 21845 13955 21879
rect 14841 21845 14875 21879
rect 15117 21845 15151 21879
rect 17141 21845 17175 21879
rect 18629 21845 18663 21879
rect 20453 21845 20487 21879
rect 23397 21845 23431 21879
rect 23489 21845 23523 21879
rect 24961 21845 24995 21879
rect 30389 21845 30423 21879
rect 4629 21641 4663 21675
rect 6377 21641 6411 21675
rect 9597 21641 9631 21675
rect 10241 21641 10275 21675
rect 13645 21641 13679 21675
rect 15193 21641 15227 21675
rect 15669 21641 15703 21675
rect 19073 21641 19107 21675
rect 19993 21641 20027 21675
rect 20361 21641 20395 21675
rect 21005 21641 21039 21675
rect 21189 21641 21223 21675
rect 21833 21641 21867 21675
rect 22201 21641 22235 21675
rect 24133 21641 24167 21675
rect 25053 21641 25087 21675
rect 25881 21641 25915 21675
rect 15393 21573 15427 21607
rect 18705 21573 18739 21607
rect 18797 21573 18831 21607
rect 19625 21573 19659 21607
rect 20085 21573 20119 21607
rect 20637 21573 20671 21607
rect 22385 21573 22419 21607
rect 23765 21573 23799 21607
rect 24777 21573 24811 21607
rect 1685 21505 1719 21539
rect 5365 21505 5399 21539
rect 5549 21505 5583 21539
rect 6561 21505 6595 21539
rect 7012 21505 7046 21539
rect 8217 21505 8251 21539
rect 8484 21505 8518 21539
rect 9873 21505 9907 21539
rect 11529 21505 11563 21539
rect 13921 21505 13955 21539
rect 14841 21505 14875 21539
rect 15485 21505 15519 21539
rect 18521 21505 18555 21539
rect 18889 21505 18923 21539
rect 19533 21505 19567 21539
rect 19717 21505 19751 21539
rect 20177 21505 20211 21539
rect 20453 21505 20487 21539
rect 20729 21505 20763 21539
rect 20821 21505 20855 21539
rect 21097 21505 21131 21539
rect 21373 21505 21407 21539
rect 22036 21505 22070 21539
rect 22293 21505 22327 21539
rect 22569 21505 22603 21539
rect 22661 21505 22695 21539
rect 23949 21505 23983 21539
rect 24501 21505 24535 21539
rect 24685 21505 24719 21539
rect 24869 21505 24903 21539
rect 26065 21505 26099 21539
rect 26157 21505 26191 21539
rect 30481 21505 30515 21539
rect 5273 21437 5307 21471
rect 5457 21437 5491 21471
rect 6745 21437 6779 21471
rect 9781 21437 9815 21471
rect 11805 21437 11839 21471
rect 13553 21437 13587 21471
rect 13829 21437 13863 21471
rect 14013 21437 14047 21471
rect 14105 21437 14139 21471
rect 14289 21437 14323 21471
rect 21557 21437 21591 21471
rect 26525 21437 26559 21471
rect 29653 21437 29687 21471
rect 15025 21369 15059 21403
rect 19809 21369 19843 21403
rect 22477 21369 22511 21403
rect 1501 21301 1535 21335
rect 8125 21301 8159 21335
rect 15209 21301 15243 21335
rect 5365 21097 5399 21131
rect 6101 21097 6135 21131
rect 12357 21097 12391 21131
rect 20361 21097 20395 21131
rect 22661 21097 22695 21131
rect 26157 21097 26191 21131
rect 9321 21029 9355 21063
rect 24961 21029 24995 21063
rect 5457 20961 5491 20995
rect 8953 20961 8987 20995
rect 18705 20961 18739 20995
rect 19809 20961 19843 20995
rect 21741 20961 21775 20995
rect 21925 20961 21959 20995
rect 22293 20961 22327 20995
rect 22385 20961 22419 20995
rect 25053 20961 25087 20995
rect 26341 20961 26375 20995
rect 26801 20961 26835 20995
rect 1685 20893 1719 20927
rect 3985 20893 4019 20927
rect 6193 20893 6227 20927
rect 9689 20893 9723 20927
rect 12265 20893 12299 20927
rect 14933 20893 14967 20927
rect 15485 20893 15519 20927
rect 16957 20893 16991 20927
rect 18981 20893 19015 20927
rect 19993 20893 20027 20927
rect 21649 20893 21683 20927
rect 21833 20893 21867 20927
rect 24409 20893 24443 20927
rect 24777 20893 24811 20927
rect 26433 20893 26467 20927
rect 26709 20893 26743 20927
rect 26893 20893 26927 20927
rect 30205 20893 30239 20927
rect 4252 20825 4286 20859
rect 6285 20825 6319 20859
rect 17233 20825 17267 20859
rect 18889 20825 18923 20859
rect 20177 20825 20211 20859
rect 22845 20825 22879 20859
rect 23029 20825 23063 20859
rect 24593 20825 24627 20859
rect 24685 20825 24719 20859
rect 1501 20757 1535 20791
rect 9413 20757 9447 20791
rect 9597 20757 9631 20791
rect 14749 20757 14783 20791
rect 15669 20757 15703 20791
rect 19257 20757 19291 20791
rect 22569 20757 22603 20791
rect 25697 20757 25731 20791
rect 30389 20757 30423 20791
rect 8125 20553 8159 20587
rect 10057 20553 10091 20587
rect 17417 20553 17451 20587
rect 18245 20553 18279 20587
rect 20545 20553 20579 20587
rect 25237 20553 25271 20587
rect 26065 20553 26099 20587
rect 26341 20553 26375 20587
rect 14749 20485 14783 20519
rect 16497 20485 16531 20519
rect 18337 20485 18371 20519
rect 20269 20485 20303 20519
rect 22569 20485 22603 20519
rect 22661 20485 22695 20519
rect 25329 20485 25363 20519
rect 25881 20485 25915 20519
rect 6377 20417 6411 20451
rect 8309 20417 8343 20451
rect 11345 20417 11379 20451
rect 12817 20417 12851 20451
rect 17601 20417 17635 20451
rect 19433 20417 19467 20451
rect 19993 20417 20027 20451
rect 20177 20417 20211 20451
rect 20361 20417 20395 20451
rect 22385 20417 22419 20451
rect 22753 20417 22787 20451
rect 25697 20417 25731 20451
rect 26157 20417 26191 20451
rect 26341 20417 26375 20451
rect 6653 20349 6687 20383
rect 8585 20349 8619 20383
rect 10609 20349 10643 20383
rect 12725 20349 12759 20383
rect 14473 20349 14507 20383
rect 18429 20349 18463 20383
rect 23029 20349 23063 20383
rect 23305 20349 23339 20383
rect 24777 20349 24811 20383
rect 25421 20349 25455 20383
rect 10333 20281 10367 20315
rect 17877 20281 17911 20315
rect 10149 20213 10183 20247
rect 11253 20213 11287 20247
rect 13185 20213 13219 20247
rect 19533 20213 19567 20247
rect 22937 20213 22971 20247
rect 24869 20213 24903 20247
rect 6745 20009 6779 20043
rect 8585 20009 8619 20043
rect 10241 20009 10275 20043
rect 15209 20009 15243 20043
rect 15853 20009 15887 20043
rect 21005 20009 21039 20043
rect 22845 20009 22879 20043
rect 23673 20009 23707 20043
rect 24133 20009 24167 20043
rect 8953 19941 8987 19975
rect 12081 19941 12115 19975
rect 30389 19941 30423 19975
rect 7757 19873 7791 19907
rect 7941 19873 7975 19907
rect 9505 19873 9539 19907
rect 11989 19873 12023 19907
rect 13093 19873 13127 19907
rect 14565 19873 14599 19907
rect 14749 19873 14783 19907
rect 17509 19873 17543 19907
rect 19257 19873 19291 19907
rect 21097 19873 21131 19907
rect 23489 19873 23523 19907
rect 6653 19805 6687 19839
rect 8125 19805 8159 19839
rect 8217 19805 8251 19839
rect 8769 19805 8803 19839
rect 9321 19805 9355 19839
rect 12357 19805 12391 19839
rect 12909 19805 12943 19839
rect 14841 19805 14875 19839
rect 15945 19805 15979 19839
rect 17417 19805 17451 19839
rect 18889 19805 18923 19839
rect 23857 19805 23891 19839
rect 24041 19805 24075 19839
rect 30205 19805 30239 19839
rect 1501 19737 1535 19771
rect 1685 19737 1719 19771
rect 11713 19737 11747 19771
rect 12081 19737 12115 19771
rect 19533 19737 19567 19771
rect 21373 19737 21407 19771
rect 7205 19669 7239 19703
rect 7941 19669 7975 19703
rect 9413 19669 9447 19703
rect 12265 19669 12299 19703
rect 13737 19669 13771 19703
rect 19073 19669 19107 19703
rect 22937 19669 22971 19703
rect 1593 19465 1627 19499
rect 5089 19465 5123 19499
rect 7389 19465 7423 19499
rect 7481 19465 7515 19499
rect 8125 19465 8159 19499
rect 12449 19465 12483 19499
rect 20913 19465 20947 19499
rect 21557 19465 21591 19499
rect 22293 19465 22327 19499
rect 26341 19465 26375 19499
rect 5273 19397 5307 19431
rect 7849 19397 7883 19431
rect 8953 19397 8987 19431
rect 16221 19397 16255 19431
rect 19625 19397 19659 19431
rect 22385 19397 22419 19431
rect 29837 19397 29871 19431
rect 1409 19329 1443 19363
rect 3341 19329 3375 19363
rect 5365 19329 5399 19363
rect 7021 19329 7055 19363
rect 7665 19329 7699 19363
rect 7941 19329 7975 19363
rect 8033 19329 8067 19363
rect 10701 19329 10735 19363
rect 11529 19329 11563 19363
rect 12357 19329 12391 19363
rect 12541 19329 12575 19363
rect 13277 19329 13311 19363
rect 13369 19329 13403 19363
rect 13645 19329 13679 19363
rect 14197 19329 14231 19363
rect 14565 19329 14599 19363
rect 14657 19329 14691 19363
rect 14933 19329 14967 19363
rect 15485 19329 15519 19363
rect 15577 19329 15611 19363
rect 15669 19329 15703 19363
rect 16681 19329 16715 19363
rect 21465 19329 21499 19363
rect 24593 19329 24627 19363
rect 30389 19329 30423 19363
rect 3617 19261 3651 19295
rect 6929 19261 6963 19295
rect 13093 19261 13127 19295
rect 13553 19261 13587 19295
rect 15117 19261 15151 19295
rect 16957 19261 16991 19295
rect 22569 19261 22603 19295
rect 24869 19261 24903 19295
rect 15853 19193 15887 19227
rect 12173 19125 12207 19159
rect 14289 19125 14323 19159
rect 14841 19125 14875 19159
rect 16221 19125 16255 19159
rect 16405 19125 16439 19159
rect 18429 19125 18463 19159
rect 21925 19125 21959 19159
rect 3801 18921 3835 18955
rect 6745 18921 6779 18955
rect 11345 18921 11379 18955
rect 13185 18921 13219 18955
rect 13277 18921 13311 18955
rect 14657 18921 14691 18955
rect 16957 18921 16991 18955
rect 19441 18921 19475 18955
rect 21557 18921 21591 18955
rect 25329 18921 25363 18955
rect 1593 18853 1627 18887
rect 4261 18853 4295 18887
rect 5641 18853 5675 18887
rect 5825 18853 5859 18887
rect 10149 18853 10183 18887
rect 10517 18853 10551 18887
rect 14473 18853 14507 18887
rect 17417 18853 17451 18887
rect 21465 18853 21499 18887
rect 25237 18853 25271 18887
rect 4813 18785 4847 18819
rect 6285 18785 6319 18819
rect 9689 18785 9723 18819
rect 11805 18785 11839 18819
rect 13553 18785 13587 18819
rect 13737 18785 13771 18819
rect 17969 18785 18003 18819
rect 19993 18785 20027 18819
rect 21005 18785 21039 18819
rect 22109 18785 22143 18819
rect 24041 18785 24075 18819
rect 24685 18785 24719 18819
rect 26249 18785 26283 18819
rect 1409 18717 1443 18751
rect 3985 18717 4019 18751
rect 4629 18717 4663 18751
rect 5365 18717 5399 18751
rect 6193 18717 6227 18751
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 6837 18717 6871 18751
rect 6929 18717 6963 18751
rect 7021 18717 7055 18751
rect 9781 18717 9815 18751
rect 10701 18717 10735 18751
rect 11069 18717 11103 18751
rect 11161 18717 11195 18751
rect 11529 18717 11563 18751
rect 11621 18717 11655 18751
rect 11897 18717 11931 18751
rect 12909 18717 12943 18751
rect 13185 18717 13219 18751
rect 13461 18717 13495 18751
rect 13645 18717 13679 18751
rect 14657 18717 14691 18751
rect 15025 18717 15059 18751
rect 16313 18717 16347 18751
rect 17141 18717 17175 18751
rect 21189 18717 21223 18751
rect 21465 18717 21499 18751
rect 21741 18717 21775 18751
rect 24133 18717 24167 18751
rect 24777 18717 24811 18751
rect 25513 18717 25547 18751
rect 26893 18717 26927 18751
rect 30205 18717 30239 18751
rect 9873 18649 9907 18683
rect 10793 18649 10827 18683
rect 10885 18649 10919 18683
rect 13001 18649 13035 18683
rect 17785 18649 17819 18683
rect 19809 18649 19843 18683
rect 20453 18649 20487 18683
rect 22385 18649 22419 18683
rect 24869 18649 24903 18683
rect 25605 18649 25639 18683
rect 4721 18581 4755 18615
rect 10333 18581 10367 18615
rect 16129 18581 16163 18615
rect 17877 18581 17911 18615
rect 19901 18581 19935 18615
rect 21281 18581 21315 18615
rect 23857 18581 23891 18615
rect 26433 18581 26467 18615
rect 30389 18581 30423 18615
rect 1593 18377 1627 18411
rect 7757 18377 7791 18411
rect 7925 18377 7959 18411
rect 8585 18377 8619 18411
rect 9321 18377 9355 18411
rect 11529 18377 11563 18411
rect 12633 18377 12667 18411
rect 13645 18377 13679 18411
rect 20269 18377 20303 18411
rect 21005 18377 21039 18411
rect 22385 18377 22419 18411
rect 22845 18377 22879 18411
rect 25789 18377 25823 18411
rect 5365 18309 5399 18343
rect 8125 18309 8159 18343
rect 21373 18309 21407 18343
rect 25421 18309 25455 18343
rect 1501 18241 1535 18275
rect 7389 18241 7423 18275
rect 8217 18241 8251 18275
rect 10195 18241 10229 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 10885 18241 10919 18275
rect 11161 18241 11195 18275
rect 11345 18241 11379 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 13093 18241 13127 18275
rect 13185 18241 13219 18275
rect 14381 18241 14415 18275
rect 16957 18241 16991 18275
rect 17325 18241 17359 18275
rect 17509 18241 17543 18275
rect 18797 18241 18831 18275
rect 19901 18241 19935 18275
rect 20361 18241 20395 18275
rect 20913 18241 20947 18275
rect 21189 18241 21223 18275
rect 22017 18241 22051 18275
rect 22201 18241 22235 18275
rect 22569 18241 22603 18275
rect 22661 18241 22695 18275
rect 22845 18241 22879 18275
rect 23397 18241 23431 18275
rect 25145 18241 25179 18275
rect 25697 18241 25731 18275
rect 30205 18241 30239 18275
rect 5825 18173 5859 18207
rect 7665 18173 7699 18207
rect 8309 18173 8343 18207
rect 9505 18173 9539 18207
rect 9597 18173 9631 18207
rect 9689 18173 9723 18207
rect 9781 18173 9815 18207
rect 10057 18173 10091 18207
rect 10701 18173 10735 18207
rect 10793 18173 10827 18207
rect 11069 18173 11103 18207
rect 11253 18173 11287 18207
rect 11713 18173 11747 18207
rect 11805 18173 11839 18207
rect 11897 18173 11931 18207
rect 11989 18173 12023 18207
rect 12449 18173 12483 18207
rect 16681 18173 16715 18207
rect 19993 18173 20027 18207
rect 20821 18173 20855 18207
rect 22293 18173 22327 18207
rect 23489 18173 23523 18207
rect 5641 18105 5675 18139
rect 7573 18105 7607 18139
rect 10333 18105 10367 18139
rect 16865 18105 16899 18139
rect 20637 18105 20671 18139
rect 23029 18105 23063 18139
rect 7481 18037 7515 18071
rect 7941 18037 7975 18071
rect 8217 18037 8251 18071
rect 10057 18037 10091 18071
rect 12817 18037 12851 18071
rect 13277 18037 13311 18071
rect 14473 18037 14507 18071
rect 16773 18037 16807 18071
rect 17509 18037 17543 18071
rect 18705 18037 18739 18071
rect 21833 18037 21867 18071
rect 30389 18037 30423 18071
rect 4997 17833 5031 17867
rect 6285 17833 6319 17867
rect 9413 17833 9447 17867
rect 18889 17833 18923 17867
rect 19349 17833 19383 17867
rect 19717 17833 19751 17867
rect 20269 17833 20303 17867
rect 5733 17697 5767 17731
rect 14289 17697 14323 17731
rect 17141 17697 17175 17731
rect 20361 17697 20395 17731
rect 24869 17697 24903 17731
rect 26617 17697 26651 17731
rect 5181 17629 5215 17663
rect 5273 17629 5307 17663
rect 5365 17629 5399 17663
rect 5641 17629 5675 17663
rect 5917 17629 5951 17663
rect 6469 17629 6503 17663
rect 6561 17629 6595 17663
rect 6653 17629 6687 17663
rect 6745 17629 6779 17663
rect 7113 17629 7147 17663
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 9597 17629 9631 17663
rect 9689 17629 9723 17663
rect 9873 17629 9907 17663
rect 9965 17629 9999 17663
rect 13737 17629 13771 17663
rect 16589 17629 16623 17663
rect 16681 17629 16715 17663
rect 16773 17629 16807 17663
rect 16865 17629 16899 17663
rect 19257 17629 19291 17663
rect 20085 17629 20119 17663
rect 27353 17629 27387 17663
rect 27445 17629 27479 17663
rect 5483 17561 5517 17595
rect 6101 17561 6135 17595
rect 14565 17561 14599 17595
rect 16313 17561 16347 17595
rect 17404 17561 17438 17595
rect 25145 17561 25179 17595
rect 27537 17561 27571 17595
rect 7021 17493 7055 17527
rect 7849 17493 7883 17527
rect 13921 17493 13955 17527
rect 17049 17493 17083 17527
rect 19901 17493 19935 17527
rect 26709 17493 26743 17527
rect 4997 17289 5031 17323
rect 5457 17289 5491 17323
rect 6193 17289 6227 17323
rect 6837 17289 6871 17323
rect 8677 17289 8711 17323
rect 11621 17289 11655 17323
rect 12909 17289 12943 17323
rect 14381 17289 14415 17323
rect 14749 17289 14783 17323
rect 15393 17289 15427 17323
rect 16221 17289 16255 17323
rect 17141 17289 17175 17323
rect 20085 17289 20119 17323
rect 22569 17289 22603 17323
rect 24777 17289 24811 17323
rect 7757 17221 7791 17255
rect 7941 17221 7975 17255
rect 9321 17221 9355 17255
rect 9597 17221 9631 17255
rect 10701 17221 10735 17255
rect 12265 17221 12299 17255
rect 14013 17221 14047 17255
rect 4629 17153 4663 17187
rect 5457 17153 5491 17187
rect 5641 17153 5675 17187
rect 6009 17153 6043 17187
rect 6193 17153 6227 17187
rect 6377 17153 6411 17187
rect 6653 17153 6687 17187
rect 7389 17153 7423 17187
rect 7481 17153 7515 17187
rect 7665 17153 7699 17187
rect 8033 17153 8067 17187
rect 8401 17153 8435 17187
rect 8585 17153 8619 17187
rect 8861 17153 8895 17187
rect 9137 17153 9171 17187
rect 9873 17153 9907 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 11529 17153 11563 17187
rect 11805 17153 11839 17187
rect 12412 17153 12446 17187
rect 13093 17153 13127 17187
rect 13185 17153 13219 17187
rect 13277 17153 13311 17187
rect 13553 17153 13587 17187
rect 13737 17153 13771 17187
rect 15301 17153 15335 17187
rect 16129 17153 16163 17187
rect 17325 17153 17359 17187
rect 17509 17153 17543 17187
rect 20729 17153 20763 17187
rect 22201 17153 22235 17187
rect 22661 17153 22695 17187
rect 22845 17153 22879 17187
rect 23581 17153 23615 17187
rect 24961 17153 24995 17187
rect 25053 17153 25087 17187
rect 25329 17153 25363 17187
rect 30205 17153 30239 17187
rect 1409 17085 1443 17119
rect 1685 17085 1719 17119
rect 4721 17085 4755 17119
rect 6469 17085 6503 17119
rect 7297 17085 7331 17119
rect 8953 17085 8987 17119
rect 9045 17085 9079 17119
rect 9413 17085 9447 17119
rect 9505 17085 9539 17119
rect 9689 17085 9723 17119
rect 12633 17085 12667 17119
rect 14841 17085 14875 17119
rect 14933 17085 14967 17119
rect 17601 17085 17635 17119
rect 18337 17085 18371 17119
rect 18613 17085 18647 17119
rect 22017 17085 22051 17119
rect 22109 17085 22143 17119
rect 7757 17017 7791 17051
rect 8493 17017 8527 17051
rect 11805 17017 11839 17051
rect 25237 17017 25271 17051
rect 30389 17017 30423 17051
rect 7297 16949 7331 16983
rect 12541 16949 12575 16983
rect 13415 16949 13449 16983
rect 20177 16949 20211 16983
rect 22753 16949 22787 16983
rect 23673 16949 23707 16983
rect 24041 16949 24075 16983
rect 7849 16745 7883 16779
rect 8217 16745 8251 16779
rect 9597 16745 9631 16779
rect 12909 16745 12943 16779
rect 13093 16745 13127 16779
rect 15577 16745 15611 16779
rect 19349 16745 19383 16779
rect 21511 16745 21545 16779
rect 21649 16745 21683 16779
rect 25605 16745 25639 16779
rect 12449 16677 12483 16711
rect 19533 16677 19567 16711
rect 20361 16677 20395 16711
rect 21005 16677 21039 16711
rect 23397 16677 23431 16711
rect 24133 16677 24167 16711
rect 25697 16677 25731 16711
rect 26157 16677 26191 16711
rect 26617 16677 26651 16711
rect 7941 16609 7975 16643
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 10977 16609 11011 16643
rect 17969 16609 18003 16643
rect 19993 16609 20027 16643
rect 20637 16609 20671 16643
rect 20729 16609 20763 16643
rect 21741 16609 21775 16643
rect 22109 16609 22143 16643
rect 22937 16609 22971 16643
rect 23765 16609 23799 16643
rect 23857 16609 23891 16643
rect 25421 16609 25455 16643
rect 25513 16609 25547 16643
rect 25973 16609 26007 16643
rect 26433 16609 26467 16643
rect 26525 16609 26559 16643
rect 26985 16609 27019 16643
rect 1685 16541 1719 16575
rect 5365 16541 5399 16575
rect 7849 16541 7883 16575
rect 9505 16541 9539 16575
rect 9689 16541 9723 16575
rect 10782 16541 10816 16575
rect 11161 16541 11195 16575
rect 11345 16541 11379 16575
rect 11989 16541 12023 16575
rect 12357 16541 12391 16575
rect 12541 16541 12575 16575
rect 16957 16541 16991 16575
rect 17877 16541 17911 16575
rect 18429 16541 18463 16575
rect 18797 16541 18831 16575
rect 19257 16541 19291 16575
rect 19717 16541 19751 16575
rect 19809 16541 19843 16575
rect 20085 16541 20119 16575
rect 20545 16541 20579 16575
rect 20821 16541 20855 16575
rect 22201 16541 22235 16575
rect 22385 16541 22419 16575
rect 22687 16541 22721 16575
rect 22845 16541 22879 16575
rect 23673 16541 23707 16575
rect 23949 16541 23983 16575
rect 24869 16541 24903 16575
rect 24961 16541 24995 16575
rect 25145 16541 25179 16575
rect 25237 16541 25271 16575
rect 25789 16541 25823 16575
rect 30481 16541 30515 16575
rect 11253 16473 11287 16507
rect 12817 16473 12851 16507
rect 13077 16473 13111 16507
rect 13277 16473 13311 16507
rect 13829 16473 13863 16507
rect 14289 16473 14323 16507
rect 21189 16473 21223 16507
rect 21373 16473 21407 16507
rect 22477 16473 22511 16507
rect 22569 16473 22603 16507
rect 1501 16405 1535 16439
rect 5273 16405 5307 16439
rect 10517 16405 10551 16439
rect 13553 16405 13587 16439
rect 17049 16405 17083 16439
rect 24685 16405 24719 16439
rect 30297 16405 30331 16439
rect 7481 16201 7515 16235
rect 18705 16201 18739 16235
rect 20545 16201 20579 16235
rect 22753 16201 22787 16235
rect 23581 16201 23615 16235
rect 24803 16201 24837 16235
rect 13921 16133 13955 16167
rect 20913 16133 20947 16167
rect 22385 16133 22419 16167
rect 22569 16133 22603 16167
rect 24593 16133 24627 16167
rect 1685 16065 1719 16099
rect 5917 16065 5951 16099
rect 6101 16065 6135 16099
rect 7021 16065 7055 16099
rect 9505 16065 9539 16099
rect 9597 16065 9631 16099
rect 9873 16065 9907 16099
rect 10333 16065 10367 16099
rect 11989 16065 12023 16099
rect 13553 16065 13587 16099
rect 14197 16065 14231 16099
rect 14657 16065 14691 16099
rect 14933 16065 14967 16099
rect 15025 16065 15059 16099
rect 16037 16065 16071 16099
rect 16129 16065 16163 16099
rect 16681 16065 16715 16099
rect 18981 16065 19015 16099
rect 20361 16065 20395 16099
rect 20545 16065 20579 16099
rect 20729 16065 20763 16099
rect 23397 16065 23431 16099
rect 23581 16065 23615 16099
rect 23857 16065 23891 16099
rect 26341 16065 26375 16099
rect 30205 16065 30239 16099
rect 3341 15997 3375 16031
rect 4813 15997 4847 16031
rect 5089 15997 5123 16031
rect 5733 15997 5767 16031
rect 6377 15997 6411 16031
rect 10885 15997 10919 16031
rect 11529 15997 11563 16031
rect 13277 15997 13311 16031
rect 15301 15997 15335 16031
rect 16221 15997 16255 16031
rect 16957 15997 16991 16031
rect 6653 15929 6687 15963
rect 7389 15929 7423 15963
rect 9781 15929 9815 15963
rect 14841 15929 14875 15963
rect 18429 15929 18463 15963
rect 24961 15929 24995 15963
rect 1501 15861 1535 15895
rect 5181 15861 5215 15895
rect 6009 15861 6043 15895
rect 6837 15861 6871 15895
rect 9321 15861 9355 15895
rect 11713 15861 11747 15895
rect 14473 15861 14507 15895
rect 15669 15861 15703 15895
rect 21097 15861 21131 15895
rect 23765 15861 23799 15895
rect 24777 15861 24811 15895
rect 25881 15861 25915 15895
rect 26249 15861 26283 15895
rect 30389 15861 30423 15895
rect 4721 15657 4755 15691
rect 5181 15657 5215 15691
rect 9308 15657 9342 15691
rect 10885 15657 10919 15691
rect 11069 15657 11103 15691
rect 25697 15657 25731 15691
rect 1593 15589 1627 15623
rect 6377 15589 6411 15623
rect 7573 15589 7607 15623
rect 10793 15589 10827 15623
rect 5365 15521 5399 15555
rect 5549 15521 5583 15555
rect 6469 15521 6503 15555
rect 7665 15521 7699 15555
rect 7941 15521 7975 15555
rect 9045 15521 9079 15555
rect 11805 15521 11839 15555
rect 14197 15521 14231 15555
rect 14657 15521 14691 15555
rect 17049 15521 17083 15555
rect 17325 15521 17359 15555
rect 26065 15521 26099 15555
rect 1409 15453 1443 15487
rect 4905 15453 4939 15487
rect 4997 15453 5031 15487
rect 5273 15453 5307 15487
rect 5641 15453 5675 15487
rect 5733 15453 5767 15487
rect 5825 15453 5859 15487
rect 6929 15453 6963 15487
rect 7113 15453 7147 15487
rect 7205 15453 7239 15487
rect 7849 15453 7883 15487
rect 8033 15453 8067 15487
rect 8125 15453 8159 15487
rect 11345 15453 11379 15487
rect 11621 15453 11655 15487
rect 14289 15453 14323 15487
rect 15393 15453 15427 15487
rect 16957 15453 16991 15487
rect 18889 15453 18923 15487
rect 21005 15453 21039 15487
rect 22017 15453 22051 15487
rect 22293 15453 22327 15487
rect 25145 15453 25179 15487
rect 25329 15453 25363 15487
rect 25513 15453 25547 15487
rect 25605 15453 25639 15487
rect 25881 15453 25915 15487
rect 25973 15453 26007 15487
rect 26157 15453 26191 15487
rect 30205 15453 30239 15487
rect 6009 15385 6043 15419
rect 7389 15385 7423 15419
rect 12081 15385 12115 15419
rect 22569 15385 22603 15419
rect 25237 15385 25271 15419
rect 7021 15317 7055 15351
rect 11529 15317 11563 15351
rect 13553 15317 13587 15351
rect 15577 15317 15611 15351
rect 19073 15317 19107 15351
rect 21097 15317 21131 15351
rect 22201 15317 22235 15351
rect 24041 15317 24075 15351
rect 24961 15317 24995 15351
rect 30389 15317 30423 15351
rect 5641 15113 5675 15147
rect 11713 15113 11747 15147
rect 12265 15113 12299 15147
rect 12817 15113 12851 15147
rect 13093 15113 13127 15147
rect 13553 15113 13587 15147
rect 15393 15113 15427 15147
rect 19073 15113 19107 15147
rect 21465 15113 21499 15147
rect 21833 15113 21867 15147
rect 22201 15113 22235 15147
rect 7389 15045 7423 15079
rect 10609 15045 10643 15079
rect 10977 15045 11011 15079
rect 16313 15045 16347 15079
rect 19441 15045 19475 15079
rect 4813 14977 4847 15011
rect 4905 14977 4939 15011
rect 5181 14977 5215 15011
rect 5825 14977 5859 15011
rect 6009 14977 6043 15011
rect 6101 14977 6135 15011
rect 7573 14977 7607 15011
rect 7665 14977 7699 15011
rect 8217 14977 8251 15011
rect 8401 14977 8435 15011
rect 11621 14977 11655 15011
rect 12449 14977 12483 15011
rect 12725 14977 12759 15011
rect 13461 14977 13495 15011
rect 14197 14977 14231 15011
rect 14933 14977 14967 15011
rect 15577 14977 15611 15011
rect 15669 14977 15703 15011
rect 15761 14977 15795 15011
rect 15945 14977 15979 15011
rect 16037 14977 16071 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 18705 14977 18739 15011
rect 19165 14977 19199 15011
rect 21189 14977 21223 15011
rect 24041 14977 24075 15011
rect 13645 14909 13679 14943
rect 15025 14909 15059 14943
rect 16313 14909 16347 14943
rect 18429 14909 18463 14943
rect 18613 14909 18647 14943
rect 22293 14909 22327 14943
rect 22385 14909 22419 14943
rect 5089 14841 5123 14875
rect 7389 14841 7423 14875
rect 15301 14841 15335 14875
rect 20913 14841 20947 14875
rect 4629 14773 4663 14807
rect 8309 14773 8343 14807
rect 9321 14773 9355 14807
rect 11253 14773 11287 14807
rect 14289 14773 14323 14807
rect 16129 14773 16163 14807
rect 16865 14773 16899 14807
rect 24317 14773 24351 14807
rect 24501 14773 24535 14807
rect 4905 14569 4939 14603
rect 6009 14569 6043 14603
rect 6653 14569 6687 14603
rect 7205 14569 7239 14603
rect 8401 14569 8435 14603
rect 9321 14569 9355 14603
rect 9689 14569 9723 14603
rect 14657 14569 14691 14603
rect 16773 14569 16807 14603
rect 17969 14569 18003 14603
rect 20545 14569 20579 14603
rect 22017 14569 22051 14603
rect 24593 14569 24627 14603
rect 26065 14569 26099 14603
rect 5365 14501 5399 14535
rect 7021 14501 7055 14535
rect 9413 14501 9447 14535
rect 18429 14501 18463 14535
rect 30389 14501 30423 14535
rect 5641 14433 5675 14467
rect 7573 14433 7607 14467
rect 8769 14433 8803 14467
rect 9229 14433 9263 14467
rect 16037 14433 16071 14467
rect 16497 14433 16531 14467
rect 16589 14433 16623 14467
rect 18797 14433 18831 14467
rect 22845 14433 22879 14467
rect 25053 14433 25087 14467
rect 25329 14433 25363 14467
rect 1685 14365 1719 14399
rect 4261 14365 4295 14399
rect 5549 14365 5583 14399
rect 5733 14365 5767 14399
rect 5825 14365 5859 14399
rect 6561 14365 6595 14399
rect 7113 14365 7147 14399
rect 7665 14365 7699 14399
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 8585 14365 8619 14399
rect 8953 14365 8987 14399
rect 10517 14365 10551 14399
rect 12265 14365 12299 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 14749 14365 14783 14399
rect 16129 14365 16163 14399
rect 16313 14365 16347 14399
rect 16405 14365 16439 14399
rect 16865 14365 16899 14399
rect 17049 14365 17083 14399
rect 17141 14365 17175 14399
rect 17325 14365 17359 14399
rect 17417 14365 17451 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 19073 14365 19107 14399
rect 19257 14365 19291 14399
rect 21097 14365 21131 14399
rect 21925 14365 21959 14399
rect 22201 14365 22235 14399
rect 22385 14365 22419 14399
rect 22661 14365 22695 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 24869 14365 24903 14399
rect 25421 14365 25455 14399
rect 30205 14365 30239 14399
rect 6193 14297 6227 14331
rect 6377 14297 6411 14331
rect 7757 14297 7791 14331
rect 8309 14297 8343 14331
rect 17601 14297 17635 14331
rect 21373 14297 21407 14331
rect 22293 14297 22327 14331
rect 22523 14297 22557 14331
rect 25697 14297 25731 14331
rect 25881 14297 25915 14331
rect 1501 14229 1535 14263
rect 7941 14229 7975 14263
rect 9045 14229 9079 14263
rect 10609 14229 10643 14263
rect 12357 14229 12391 14263
rect 14197 14229 14231 14263
rect 18337 14229 18371 14263
rect 18981 14229 19015 14263
rect 21741 14229 21775 14263
rect 24409 14229 24443 14263
rect 1593 14025 1627 14059
rect 5641 14025 5675 14059
rect 7941 14025 7975 14059
rect 8109 14025 8143 14059
rect 14381 14025 14415 14059
rect 15025 14025 15059 14059
rect 17601 14025 17635 14059
rect 20361 14025 20395 14059
rect 4721 13957 4755 13991
rect 8309 13957 8343 13991
rect 17417 13957 17451 13991
rect 18797 13957 18831 13991
rect 19717 13957 19751 13991
rect 22845 13957 22879 13991
rect 25053 13957 25087 13991
rect 1409 13889 1443 13923
rect 5549 13889 5583 13923
rect 5733 13889 5767 13923
rect 9505 13889 9539 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14933 13889 14967 13923
rect 15117 13889 15151 13923
rect 17141 13889 17175 13923
rect 17785 13889 17819 13923
rect 17969 13889 18003 13923
rect 18061 13889 18095 13923
rect 18981 13889 19015 13923
rect 20453 13889 20487 13923
rect 20913 13889 20947 13923
rect 22661 13889 22695 13923
rect 24593 13889 24627 13923
rect 24777 13889 24811 13923
rect 25329 13889 25363 13923
rect 30481 13889 30515 13923
rect 4997 13821 5031 13855
rect 9781 13821 9815 13855
rect 11529 13821 11563 13855
rect 11805 13821 11839 13855
rect 14013 13821 14047 13855
rect 17325 13821 17359 13855
rect 19257 13821 19291 13855
rect 25053 13821 25087 13855
rect 19441 13753 19475 13787
rect 3249 13685 3283 13719
rect 8125 13685 8159 13719
rect 11253 13685 11287 13719
rect 13277 13685 13311 13719
rect 16957 13685 16991 13719
rect 17141 13685 17175 13719
rect 19165 13685 19199 13719
rect 21005 13685 21039 13719
rect 22477 13685 22511 13719
rect 24685 13685 24719 13719
rect 25237 13685 25271 13719
rect 30297 13685 30331 13719
rect 4261 13481 4295 13515
rect 6193 13481 6227 13515
rect 8953 13481 8987 13515
rect 10333 13481 10367 13515
rect 11897 13481 11931 13515
rect 15577 13481 15611 13515
rect 15761 13481 15795 13515
rect 17325 13481 17359 13515
rect 9045 13413 9079 13447
rect 10793 13413 10827 13447
rect 15853 13413 15887 13447
rect 21741 13413 21775 13447
rect 23673 13413 23707 13447
rect 5181 13345 5215 13379
rect 5733 13345 5767 13379
rect 13093 13345 13127 13379
rect 17785 13345 17819 13379
rect 18521 13345 18555 13379
rect 19993 13345 20027 13379
rect 22569 13345 22603 13379
rect 23305 13345 23339 13379
rect 23765 13345 23799 13379
rect 25421 13345 25455 13379
rect 1685 13277 1719 13311
rect 4353 13277 4387 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 10517 13277 10551 13311
rect 10609 13277 10643 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11621 13277 11655 13311
rect 12081 13277 12115 13311
rect 12817 13277 12851 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 15301 13277 15335 13311
rect 16037 13277 16071 13311
rect 16221 13277 16255 13311
rect 17325 13277 17359 13311
rect 17417 13277 17451 13311
rect 17693 13277 17727 13311
rect 17877 13277 17911 13311
rect 18613 13277 18647 13311
rect 22109 13277 22143 13311
rect 22201 13277 22235 13311
rect 22845 13277 22879 13311
rect 23029 13277 23063 13311
rect 24409 13277 24443 13311
rect 24685 13277 24719 13311
rect 25513 13277 25547 13311
rect 30205 13277 30239 13311
rect 6009 13209 6043 13243
rect 6225 13209 6259 13243
rect 6561 13209 6595 13243
rect 9413 13209 9447 13243
rect 15025 13209 15059 13243
rect 15393 13209 15427 13243
rect 17601 13209 17635 13243
rect 20269 13209 20303 13243
rect 22293 13209 22327 13243
rect 22431 13209 22465 13243
rect 1501 13141 1535 13175
rect 6377 13141 6411 13175
rect 12449 13141 12483 13175
rect 12909 13141 12943 13175
rect 14657 13141 14691 13175
rect 15301 13141 15335 13175
rect 15593 13141 15627 13175
rect 17141 13141 17175 13175
rect 18981 13141 19015 13175
rect 21925 13141 21959 13175
rect 22661 13141 22695 13175
rect 24501 13141 24535 13175
rect 24869 13141 24903 13175
rect 25145 13141 25179 13175
rect 30389 13141 30423 13175
rect 3249 12937 3283 12971
rect 5365 12937 5399 12971
rect 10609 12937 10643 12971
rect 13277 12937 13311 12971
rect 15117 12937 15151 12971
rect 18797 12937 18831 12971
rect 20545 12937 20579 12971
rect 20913 12937 20947 12971
rect 21281 12937 21315 12971
rect 21373 12937 21407 12971
rect 23857 12937 23891 12971
rect 24961 12937 24995 12971
rect 30297 12937 30331 12971
rect 5181 12869 5215 12903
rect 9045 12869 9079 12903
rect 10425 12869 10459 12903
rect 13921 12869 13955 12903
rect 16865 12869 16899 12903
rect 19283 12869 19317 12903
rect 22201 12869 22235 12903
rect 22753 12869 22787 12903
rect 1685 12801 1719 12835
rect 4997 12801 5031 12835
rect 5273 12801 5307 12835
rect 5549 12801 5583 12835
rect 5733 12801 5767 12835
rect 6377 12801 6411 12835
rect 6837 12801 6871 12835
rect 7021 12801 7055 12835
rect 7113 12801 7147 12835
rect 7389 12801 7423 12835
rect 7481 12801 7515 12835
rect 7757 12801 7791 12835
rect 8861 12801 8895 12835
rect 11529 12801 11563 12835
rect 13461 12801 13495 12835
rect 13737 12801 13771 12835
rect 14105 12801 14139 12835
rect 14197 12801 14231 12835
rect 14749 12801 14783 12835
rect 14933 12801 14967 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 17325 12801 17359 12835
rect 17509 12801 17543 12835
rect 18981 12801 19015 12835
rect 19073 12801 19107 12835
rect 19165 12801 19199 12835
rect 19441 12801 19475 12835
rect 20729 12801 20763 12835
rect 22385 12801 22419 12835
rect 22661 12801 22695 12835
rect 22845 12801 22879 12835
rect 23397 12801 23431 12835
rect 24317 12801 24351 12835
rect 24869 12801 24903 12835
rect 25145 12801 25179 12835
rect 30389 12801 30423 12835
rect 4721 12733 4755 12767
rect 8309 12733 8343 12767
rect 13553 12733 13587 12767
rect 13645 12733 13679 12767
rect 13921 12733 13955 12767
rect 14657 12733 14691 12767
rect 21465 12733 21499 12767
rect 24777 12733 24811 12767
rect 7205 12665 7239 12699
rect 8585 12665 8619 12699
rect 10057 12665 10091 12699
rect 1501 12597 1535 12631
rect 7665 12597 7699 12631
rect 8769 12597 8803 12631
rect 9229 12597 9263 12631
rect 10425 12597 10459 12631
rect 11621 12597 11655 12631
rect 11989 12597 12023 12631
rect 22477 12597 22511 12631
rect 23489 12597 23523 12631
rect 24593 12597 24627 12631
rect 25329 12597 25363 12631
rect 6377 12393 6411 12427
rect 8217 12393 8251 12427
rect 8493 12393 8527 12427
rect 9321 12393 9355 12427
rect 10517 12393 10551 12427
rect 10701 12393 10735 12427
rect 11161 12393 11195 12427
rect 12817 12393 12851 12427
rect 13553 12393 13587 12427
rect 13921 12393 13955 12427
rect 14676 12393 14710 12427
rect 16221 12393 16255 12427
rect 17049 12393 17083 12427
rect 17785 12393 17819 12427
rect 21005 12393 21039 12427
rect 25145 12393 25179 12427
rect 8033 12325 8067 12359
rect 10425 12325 10459 12359
rect 14565 12325 14599 12359
rect 15853 12325 15887 12359
rect 17601 12325 17635 12359
rect 20361 12325 20395 12359
rect 23765 12325 23799 12359
rect 7757 12257 7791 12291
rect 8585 12257 8619 12291
rect 12081 12257 12115 12291
rect 12541 12257 12575 12291
rect 13461 12257 13495 12291
rect 14473 12257 14507 12291
rect 19349 12257 19383 12291
rect 20269 12257 20303 12291
rect 23581 12257 23615 12291
rect 5825 12189 5859 12223
rect 6009 12189 6043 12223
rect 8309 12189 8343 12223
rect 8401 12189 8435 12223
rect 9505 12189 9539 12223
rect 9597 12189 9631 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 9965 12189 9999 12223
rect 10241 12189 10275 12223
rect 11069 12189 11103 12223
rect 11989 12189 12023 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 13001 12189 13035 12223
rect 13093 12189 13127 12223
rect 13829 12189 13863 12223
rect 13921 12189 13955 12223
rect 14841 12189 14875 12223
rect 17233 12189 17267 12223
rect 17509 12189 17543 12223
rect 19257 12189 19291 12223
rect 19441 12189 19475 12223
rect 19901 12189 19935 12223
rect 20545 12189 20579 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 20923 12183 20957 12217
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 25421 12189 25455 12223
rect 25513 12189 25547 12223
rect 6193 12121 6227 12155
rect 10057 12121 10091 12155
rect 10885 12121 10919 12155
rect 13185 12121 13219 12155
rect 13303 12121 13337 12155
rect 16221 12121 16255 12155
rect 17969 12121 18003 12155
rect 20085 12121 20119 12155
rect 24041 12121 24075 12155
rect 24961 12121 24995 12155
rect 25177 12121 25211 12155
rect 25697 12121 25731 12155
rect 6009 12053 6043 12087
rect 6393 12053 6427 12087
rect 6561 12053 6595 12087
rect 10685 12053 10719 12087
rect 11529 12053 11563 12087
rect 12357 12053 12391 12087
rect 14197 12053 14231 12087
rect 16405 12053 16439 12087
rect 17417 12053 17451 12087
rect 17769 12053 17803 12087
rect 21373 12053 21407 12087
rect 25329 12053 25363 12087
rect 25421 12053 25455 12087
rect 5273 11849 5307 11883
rect 6377 11849 6411 11883
rect 7474 11849 7508 11883
rect 7665 11849 7699 11883
rect 9045 11849 9079 11883
rect 9873 11849 9907 11883
rect 13461 11849 13495 11883
rect 17233 11849 17267 11883
rect 17877 11849 17911 11883
rect 19257 11849 19291 11883
rect 23587 11849 23621 11883
rect 23857 11849 23891 11883
rect 7389 11781 7423 11815
rect 20085 11781 20119 11815
rect 20269 11781 20303 11815
rect 24869 11781 24903 11815
rect 1409 11713 1443 11747
rect 2973 11713 3007 11747
rect 5181 11713 5215 11747
rect 5641 11713 5675 11747
rect 6837 11713 6871 11747
rect 7297 11713 7331 11747
rect 7573 11713 7607 11747
rect 8033 11713 8067 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 8861 11713 8895 11747
rect 10241 11713 10275 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 13461 11713 13495 11747
rect 13645 11713 13679 11747
rect 16773 11713 16807 11747
rect 17325 11713 17359 11747
rect 17877 11713 17911 11747
rect 18061 11713 18095 11747
rect 18153 11713 18187 11747
rect 18613 11713 18647 11747
rect 19809 11713 19843 11747
rect 21833 11713 21867 11747
rect 22753 11713 22787 11747
rect 22845 11713 22879 11747
rect 23489 11713 23523 11747
rect 23673 11713 23707 11747
rect 23765 11713 23799 11747
rect 24133 11713 24167 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 24685 11713 24719 11747
rect 24961 11713 24995 11747
rect 25145 11713 25179 11747
rect 25513 11713 25547 11747
rect 25605 11713 25639 11747
rect 25881 11713 25915 11747
rect 26985 11713 27019 11747
rect 27629 11713 27663 11747
rect 30205 11713 30239 11747
rect 3249 11645 3283 11679
rect 5365 11645 5399 11679
rect 6561 11645 6595 11679
rect 6653 11645 6687 11679
rect 6745 11645 6779 11679
rect 7849 11645 7883 11679
rect 7941 11645 7975 11679
rect 8125 11645 8159 11679
rect 8585 11645 8619 11679
rect 10149 11645 10183 11679
rect 11621 11645 11655 11679
rect 15393 11645 15427 11679
rect 17785 11645 17819 11679
rect 18245 11645 18279 11679
rect 18981 11645 19015 11679
rect 19625 11645 19659 11679
rect 19717 11645 19751 11679
rect 19901 11645 19935 11679
rect 22201 11645 22235 11679
rect 22937 11645 22971 11679
rect 23029 11645 23063 11679
rect 24041 11645 24075 11679
rect 24225 11645 24259 11679
rect 25053 11645 25087 11679
rect 4813 11577 4847 11611
rect 18521 11577 18555 11611
rect 20453 11577 20487 11611
rect 22293 11577 22327 11611
rect 23213 11577 23247 11611
rect 30389 11577 30423 11611
rect 1593 11509 1627 11543
rect 4721 11509 4755 11543
rect 5733 11509 5767 11543
rect 6101 11509 6135 11543
rect 10057 11509 10091 11543
rect 15945 11509 15979 11543
rect 17049 11509 17083 11543
rect 17417 11509 17451 11543
rect 18337 11509 18371 11543
rect 18778 11509 18812 11543
rect 18889 11509 18923 11543
rect 19441 11509 19475 11543
rect 21998 11509 22032 11543
rect 22109 11509 22143 11543
rect 25329 11509 25363 11543
rect 25789 11509 25823 11543
rect 3433 11305 3467 11339
rect 4169 11305 4203 11339
rect 4997 11305 5031 11339
rect 6285 11305 6319 11339
rect 7297 11305 7331 11339
rect 8309 11305 8343 11339
rect 8677 11305 8711 11339
rect 13461 11305 13495 11339
rect 14289 11305 14323 11339
rect 16589 11305 16623 11339
rect 18521 11305 18555 11339
rect 21649 11305 21683 11339
rect 22569 11305 22603 11339
rect 23213 11305 23247 11339
rect 23581 11305 23615 11339
rect 27169 11305 27203 11339
rect 24593 11237 24627 11271
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 8217 11169 8251 11203
rect 8401 11169 8435 11203
rect 16037 11169 16071 11203
rect 18613 11169 18647 11203
rect 25697 11169 25731 11203
rect 1685 11101 1719 11135
rect 3617 11101 3651 11135
rect 4261 11101 4295 11135
rect 4905 11101 4939 11135
rect 5549 11101 5583 11135
rect 5733 11101 5767 11135
rect 6193 11101 6227 11135
rect 6377 11101 6411 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 7021 11101 7055 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 8309 11101 8343 11135
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 13185 11101 13219 11135
rect 16313 11101 16347 11135
rect 16405 11101 16439 11135
rect 16681 11101 16715 11135
rect 18337 11101 18371 11135
rect 18429 11101 18463 11135
rect 22753 11101 22787 11135
rect 23121 11101 23155 11135
rect 23305 11101 23339 11135
rect 23489 11101 23523 11135
rect 24501 11101 24535 11135
rect 24685 11101 24719 11135
rect 25421 11101 25455 11135
rect 30481 11101 30515 11135
rect 15761 11033 15795 11067
rect 16129 11033 16163 11067
rect 21281 11033 21315 11067
rect 21465 11033 21499 11067
rect 22937 11033 22971 11067
rect 1501 10965 1535 10999
rect 11621 10965 11655 10999
rect 11989 10965 12023 10999
rect 13645 10965 13679 10999
rect 30297 10965 30331 10999
rect 6469 10761 6503 10795
rect 6837 10761 6871 10795
rect 8585 10761 8619 10795
rect 15209 10761 15243 10795
rect 18153 10761 18187 10795
rect 20069 10761 20103 10795
rect 20637 10761 20671 10795
rect 21189 10761 21223 10795
rect 21481 10761 21515 10795
rect 26249 10761 26283 10795
rect 30297 10761 30331 10795
rect 9413 10693 9447 10727
rect 10977 10693 11011 10727
rect 20269 10693 20303 10727
rect 21281 10693 21315 10727
rect 22477 10693 22511 10727
rect 23581 10693 23615 10727
rect 23765 10693 23799 10727
rect 1685 10625 1719 10659
rect 6653 10625 6687 10659
rect 6929 10625 6963 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 9045 10625 9079 10659
rect 9137 10625 9171 10659
rect 9597 10625 9631 10659
rect 9689 10625 9723 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10241 10625 10275 10659
rect 10333 10625 10367 10659
rect 10609 10625 10643 10659
rect 10885 10625 10919 10659
rect 11069 10625 11103 10659
rect 11253 10625 11287 10659
rect 11345 10625 11379 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 12449 10625 12483 10659
rect 12633 10625 12667 10659
rect 13185 10625 13219 10659
rect 13737 10625 13771 10659
rect 15301 10625 15335 10659
rect 17785 10625 17819 10659
rect 17969 10625 18003 10659
rect 18429 10625 18463 10659
rect 18613 10625 18647 10659
rect 18705 10625 18739 10659
rect 18889 10625 18923 10659
rect 20637 10625 20671 10659
rect 20821 10625 20855 10659
rect 20913 10625 20947 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 22385 10625 22419 10659
rect 22569 10625 22603 10659
rect 22661 10625 22695 10659
rect 22845 10625 22879 10659
rect 22937 10625 22971 10659
rect 23029 10625 23063 10659
rect 24593 10625 24627 10659
rect 26157 10625 26191 10659
rect 30481 10625 30515 10659
rect 8953 10557 8987 10591
rect 9229 10557 9263 10591
rect 11805 10557 11839 10591
rect 21189 10557 21223 10591
rect 23397 10557 23431 10591
rect 10057 10489 10091 10523
rect 10701 10489 10735 10523
rect 13553 10489 13587 10523
rect 14197 10489 14231 10523
rect 21833 10489 21867 10523
rect 23305 10489 23339 10523
rect 1501 10421 1535 10455
rect 8401 10421 8435 10455
rect 8769 10421 8803 10455
rect 10517 10421 10551 10455
rect 13645 10421 13679 10455
rect 13829 10421 13863 10455
rect 18245 10421 18279 10455
rect 18797 10421 18831 10455
rect 19901 10421 19935 10455
rect 20085 10421 20119 10455
rect 21005 10421 21039 10455
rect 21465 10421 21499 10455
rect 21649 10421 21683 10455
rect 22017 10421 22051 10455
rect 24685 10421 24719 10455
rect 25053 10421 25087 10455
rect 7297 10217 7331 10251
rect 9413 10217 9447 10251
rect 9781 10217 9815 10251
rect 21925 10217 21959 10251
rect 23397 10217 23431 10251
rect 23581 10217 23615 10251
rect 23673 10217 23707 10251
rect 30297 10217 30331 10251
rect 17417 10149 17451 10183
rect 23857 10149 23891 10183
rect 25513 10149 25547 10183
rect 5825 10081 5859 10115
rect 5917 10081 5951 10115
rect 6009 10081 6043 10115
rect 7757 10081 7791 10115
rect 8125 10081 8159 10115
rect 8401 10081 8435 10115
rect 14105 10081 14139 10115
rect 17233 10081 17267 10115
rect 18061 10081 18095 10115
rect 19809 10081 19843 10115
rect 20361 10081 20395 10115
rect 20545 10081 20579 10115
rect 24501 10081 24535 10115
rect 24685 10081 24719 10115
rect 24869 10081 24903 10115
rect 25329 10081 25363 10115
rect 1685 10013 1719 10047
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7113 10013 7147 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 8493 10013 8527 10047
rect 8677 10013 8711 10047
rect 9413 10013 9447 10047
rect 9597 10013 9631 10047
rect 9689 10013 9723 10047
rect 9965 10013 9999 10047
rect 11621 10013 11655 10047
rect 11805 10013 11839 10047
rect 11897 10013 11931 10047
rect 11989 10013 12023 10047
rect 12357 10013 12391 10047
rect 12541 10013 12575 10047
rect 16221 10013 16255 10047
rect 16313 10013 16347 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 16865 10013 16899 10047
rect 17141 10013 17175 10047
rect 17509 10013 17543 10047
rect 18153 10013 18187 10047
rect 18245 10013 18279 10047
rect 18337 10013 18371 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 20085 10013 20119 10047
rect 20177 10013 20211 10047
rect 20269 10013 20303 10047
rect 20637 10013 20671 10047
rect 20821 10013 20855 10047
rect 21005 10013 21039 10047
rect 21649 10013 21683 10047
rect 21741 10013 21775 10047
rect 22017 10013 22051 10047
rect 23121 10013 23155 10047
rect 24133 10013 24167 10047
rect 24777 10013 24811 10047
rect 25053 10013 25087 10047
rect 25145 10013 25179 10047
rect 25237 10013 25271 10047
rect 25697 10013 25731 10047
rect 25789 10013 25823 10047
rect 30481 10013 30515 10047
rect 7389 9945 7423 9979
rect 7573 9945 7607 9979
rect 12265 9945 12299 9979
rect 14381 9945 14415 9979
rect 16681 9945 16715 9979
rect 17233 9945 17267 9979
rect 25513 9945 25547 9979
rect 1501 9877 1535 9911
rect 5457 9877 5491 9911
rect 5549 9877 5583 9911
rect 8585 9877 8619 9911
rect 12449 9877 12483 9911
rect 15853 9877 15887 9911
rect 15945 9877 15979 9911
rect 17049 9877 17083 9911
rect 17877 9877 17911 9911
rect 21465 9877 21499 9911
rect 24501 9877 24535 9911
rect 6745 9673 6779 9707
rect 7205 9673 7239 9707
rect 10609 9673 10643 9707
rect 11161 9673 11195 9707
rect 15301 9673 15335 9707
rect 19901 9673 19935 9707
rect 22385 9673 22419 9707
rect 7849 9605 7883 9639
rect 12633 9605 12667 9639
rect 14933 9605 14967 9639
rect 15117 9605 15151 9639
rect 17785 9605 17819 9639
rect 5457 9537 5491 9571
rect 5733 9537 5767 9571
rect 5825 9537 5859 9571
rect 6561 9537 6595 9571
rect 7119 9537 7153 9571
rect 7297 9537 7331 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 10977 9537 11011 9571
rect 11069 9537 11103 9571
rect 11253 9537 11287 9571
rect 12817 9537 12851 9571
rect 13001 9537 13035 9571
rect 14841 9537 14875 9571
rect 15209 9537 15243 9571
rect 15577 9537 15611 9571
rect 15669 9537 15703 9571
rect 17049 9537 17083 9571
rect 17233 9537 17267 9571
rect 17601 9537 17635 9571
rect 19533 9537 19567 9571
rect 20361 9537 20395 9571
rect 21833 9537 21867 9571
rect 3617 9469 3651 9503
rect 5089 9469 5123 9503
rect 5365 9469 5399 9503
rect 6009 9469 6043 9503
rect 6377 9469 6411 9503
rect 10885 9469 10919 9503
rect 17325 9469 17359 9503
rect 17417 9469 17451 9503
rect 19625 9469 19659 9503
rect 20269 9469 20303 9503
rect 23029 9469 23063 9503
rect 23121 9469 23155 9503
rect 23397 9469 23431 9503
rect 24869 9469 24903 9503
rect 25605 9469 25639 9503
rect 7849 9401 7883 9435
rect 15117 9401 15151 9435
rect 19993 9401 20027 9435
rect 5549 9333 5583 9367
rect 10793 9333 10827 9367
rect 19717 9333 19751 9367
rect 20361 9333 20395 9367
rect 22109 9333 22143 9367
rect 22293 9333 22327 9367
rect 24961 9333 24995 9367
rect 1593 9129 1627 9163
rect 4629 9129 4663 9163
rect 6101 9129 6135 9163
rect 10333 9129 10367 9163
rect 16957 9129 16991 9163
rect 18337 9129 18371 9163
rect 19441 9129 19475 9163
rect 21925 9129 21959 9163
rect 22477 9129 22511 9163
rect 23305 9129 23339 9163
rect 23765 9129 23799 9163
rect 30389 9129 30423 9163
rect 5825 9061 5859 9095
rect 8493 9061 8527 9095
rect 10149 9061 10183 9095
rect 13277 9061 13311 9095
rect 18153 9061 18187 9095
rect 18797 9061 18831 9095
rect 19257 9061 19291 9095
rect 20545 9061 20579 9095
rect 8033 8993 8067 9027
rect 8401 8993 8435 9027
rect 10517 8993 10551 9027
rect 13829 8993 13863 9027
rect 15301 8993 15335 9027
rect 15577 8993 15611 9027
rect 17969 8993 18003 9027
rect 20085 8993 20119 9027
rect 20177 8993 20211 9027
rect 21649 8993 21683 9027
rect 1409 8925 1443 8959
rect 4721 8925 4755 8959
rect 5733 8925 5767 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 7573 8925 7607 8959
rect 8622 8925 8656 8959
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 10425 8925 10459 8959
rect 10609 8925 10643 8959
rect 10701 8925 10735 8959
rect 10885 8925 10919 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 13185 8925 13219 8959
rect 13461 8925 13495 8959
rect 13737 8925 13771 8959
rect 13921 8925 13955 8959
rect 15209 8925 15243 8959
rect 17144 8903 17178 8937
rect 17233 8925 17267 8959
rect 17417 8925 17451 8959
rect 17509 8925 17543 8959
rect 18245 8925 18279 8959
rect 18981 8925 19015 8959
rect 19073 8925 19107 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 20729 8925 20763 8959
rect 20821 8925 20855 8959
rect 22109 8925 22143 8959
rect 22385 8925 22419 8959
rect 22569 8925 22603 8959
rect 23489 8925 23523 8959
rect 23581 8925 23615 8959
rect 23857 8925 23891 8959
rect 30205 8925 30239 8959
rect 7757 8857 7791 8891
rect 7941 8857 7975 8891
rect 8769 8857 8803 8891
rect 9413 8857 9447 8891
rect 9505 8857 9539 8891
rect 9643 8857 9677 8891
rect 9873 8857 9907 8891
rect 12817 8857 12851 8891
rect 13027 8857 13061 8891
rect 13645 8857 13679 8891
rect 18521 8857 18555 8891
rect 18705 8857 18739 8891
rect 18797 8857 18831 8891
rect 19625 8857 19659 8891
rect 20545 8857 20579 8891
rect 9137 8789 9171 8823
rect 10793 8789 10827 8823
rect 11529 8789 11563 8823
rect 12541 8789 12575 8823
rect 18245 8789 18279 8823
rect 19425 8789 19459 8823
rect 19901 8789 19935 8823
rect 1593 8585 1627 8619
rect 7021 8585 7055 8619
rect 9045 8585 9079 8619
rect 10425 8585 10459 8619
rect 12725 8585 12759 8619
rect 13277 8585 13311 8619
rect 16037 8585 16071 8619
rect 20821 8585 20855 8619
rect 24317 8585 24351 8619
rect 5825 8517 5859 8551
rect 6041 8517 6075 8551
rect 8125 8517 8159 8551
rect 17693 8517 17727 8551
rect 22109 8517 22143 8551
rect 1409 8449 1443 8483
rect 7297 8449 7331 8483
rect 7389 8449 7423 8483
rect 7647 8449 7681 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 8401 8449 8435 8483
rect 9413 8449 9447 8483
rect 11161 8449 11195 8483
rect 13737 8449 13771 8483
rect 15669 8449 15703 8483
rect 17049 8449 17083 8483
rect 17325 8449 17359 8483
rect 17509 8449 17543 8483
rect 17785 8449 17819 8483
rect 19993 8449 20027 8483
rect 20085 8449 20119 8483
rect 21005 8449 21039 8483
rect 21189 8449 21223 8483
rect 21281 8449 21315 8483
rect 24409 8449 24443 8483
rect 30205 8449 30239 8483
rect 6377 8381 6411 8415
rect 9321 8381 9355 8415
rect 9965 8381 9999 8415
rect 11069 8381 11103 8415
rect 13185 8381 13219 8415
rect 15761 8381 15795 8415
rect 16865 8381 16899 8415
rect 19809 8381 19843 8415
rect 21833 8381 21867 8415
rect 23581 8381 23615 8415
rect 6193 8313 6227 8347
rect 7757 8313 7791 8347
rect 8309 8313 8343 8347
rect 10333 8313 10367 8347
rect 10793 8313 10827 8347
rect 12817 8313 12851 8347
rect 13369 8313 13403 8347
rect 30389 8313 30423 8347
rect 6009 8245 6043 8279
rect 7113 8245 7147 8279
rect 7573 8245 7607 8279
rect 9229 8245 9263 8279
rect 19901 8245 19935 8279
rect 6653 8041 6687 8075
rect 7389 8041 7423 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 17785 8041 17819 8075
rect 18521 8041 18555 8075
rect 20177 8041 20211 8075
rect 21373 8041 21407 8075
rect 21833 8041 21867 8075
rect 22201 8041 22235 8075
rect 22385 8041 22419 8075
rect 23029 8041 23063 8075
rect 7757 7973 7791 8007
rect 21741 7973 21775 8007
rect 22477 7973 22511 8007
rect 4721 7905 4755 7939
rect 6193 7905 6227 7939
rect 12633 7905 12667 7939
rect 12817 7905 12851 7939
rect 18061 7905 18095 7939
rect 1685 7837 1719 7871
rect 6469 7837 6503 7871
rect 6561 7837 6595 7871
rect 6745 7837 6779 7871
rect 7297 7837 7331 7871
rect 7849 7837 7883 7871
rect 17509 7837 17543 7871
rect 17601 7837 17635 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 20269 7837 20303 7871
rect 20545 7837 20579 7871
rect 21097 7837 21131 7871
rect 21281 7837 21315 7871
rect 22293 7837 22327 7871
rect 23121 7837 23155 7871
rect 22845 7769 22879 7803
rect 1501 7701 1535 7735
rect 12173 7701 12207 7735
rect 12541 7701 12575 7735
rect 17325 7701 17359 7735
rect 19717 7701 19751 7735
rect 1593 7497 1627 7531
rect 5733 7497 5767 7531
rect 13277 7497 13311 7531
rect 10517 7429 10551 7463
rect 13461 7429 13495 7463
rect 16957 7429 16991 7463
rect 19349 7429 19383 7463
rect 1409 7361 1443 7395
rect 5641 7361 5675 7395
rect 8309 7361 8343 7395
rect 8585 7361 8619 7395
rect 10609 7361 10643 7395
rect 11529 7361 11563 7395
rect 13369 7361 13403 7395
rect 16681 7361 16715 7395
rect 19073 7361 19107 7395
rect 8861 7293 8895 7327
rect 11805 7293 11839 7327
rect 8493 7225 8527 7259
rect 10333 7157 10367 7191
rect 18429 7157 18463 7191
rect 20821 7157 20855 7191
rect 8953 6953 8987 6987
rect 11897 6953 11931 6987
rect 20085 6953 20119 6987
rect 9413 6817 9447 6851
rect 9597 6817 9631 6851
rect 9321 6749 9355 6783
rect 12081 6749 12115 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 19993 6749 20027 6783
rect 9321 2601 9355 2635
rect 9965 2601 9999 2635
rect 11897 2601 11931 2635
rect 13829 2601 13863 2635
rect 17049 2601 17083 2635
rect 17693 2601 17727 2635
rect 18981 2601 19015 2635
rect 21557 2601 21591 2635
rect 15209 2533 15243 2567
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
rect 11713 2397 11747 2431
rect 12633 2397 12667 2431
rect 13277 2397 13311 2431
rect 13645 2397 13679 2431
rect 15853 2397 15887 2431
rect 16497 2397 16531 2431
rect 18429 2397 18463 2431
rect 18797 2397 18831 2431
rect 21005 2397 21039 2431
rect 21373 2397 21407 2431
rect 15025 2329 15059 2363
rect 16957 2329 16991 2363
rect 17601 2329 17635 2363
rect 10609 2261 10643 2295
rect 12449 2261 12483 2295
rect 13093 2261 13127 2295
rect 15669 2261 15703 2295
rect 16313 2261 16347 2295
rect 18245 2261 18279 2295
rect 20821 2261 20855 2295
<< metal1 >>
rect 1104 29402 30820 29424
rect 1104 29350 5324 29402
rect 5376 29350 5388 29402
rect 5440 29350 5452 29402
rect 5504 29350 5516 29402
rect 5568 29350 5580 29402
rect 5632 29350 12752 29402
rect 12804 29350 12816 29402
rect 12868 29350 12880 29402
rect 12932 29350 12944 29402
rect 12996 29350 13008 29402
rect 13060 29350 20180 29402
rect 20232 29350 20244 29402
rect 20296 29350 20308 29402
rect 20360 29350 20372 29402
rect 20424 29350 20436 29402
rect 20488 29350 27608 29402
rect 27660 29350 27672 29402
rect 27724 29350 27736 29402
rect 27788 29350 27800 29402
rect 27852 29350 27864 29402
rect 27916 29350 30820 29402
rect 1104 29328 30820 29350
rect 12342 29248 12348 29300
rect 12400 29288 12406 29300
rect 12437 29291 12495 29297
rect 12437 29288 12449 29291
rect 12400 29260 12449 29288
rect 12400 29248 12406 29260
rect 12437 29257 12449 29260
rect 12483 29257 12495 29291
rect 12437 29251 12495 29257
rect 13078 29248 13084 29300
rect 13136 29248 13142 29300
rect 14274 29248 14280 29300
rect 14332 29288 14338 29300
rect 14369 29291 14427 29297
rect 14369 29288 14381 29291
rect 14332 29260 14381 29288
rect 14332 29248 14338 29260
rect 14369 29257 14381 29260
rect 14415 29257 14427 29291
rect 14369 29251 14427 29257
rect 15746 29248 15752 29300
rect 15804 29248 15810 29300
rect 18690 29248 18696 29300
rect 18748 29288 18754 29300
rect 19429 29291 19487 29297
rect 19429 29288 19441 29291
rect 18748 29260 19441 29288
rect 18748 29248 18754 29260
rect 19429 29257 19441 29260
rect 19475 29257 19487 29291
rect 19429 29251 19487 29257
rect 19610 29248 19616 29300
rect 19668 29288 19674 29300
rect 19981 29291 20039 29297
rect 19981 29288 19993 29291
rect 19668 29260 19993 29288
rect 19668 29248 19674 29260
rect 19981 29257 19993 29260
rect 20027 29257 20039 29291
rect 19981 29251 20039 29257
rect 20622 29248 20628 29300
rect 20680 29288 20686 29300
rect 20901 29291 20959 29297
rect 20901 29288 20913 29291
rect 20680 29260 20913 29288
rect 20680 29248 20686 29260
rect 20901 29257 20913 29260
rect 20947 29257 20959 29291
rect 20901 29251 20959 29257
rect 21910 29248 21916 29300
rect 21968 29288 21974 29300
rect 22189 29291 22247 29297
rect 22189 29288 22201 29291
rect 21968 29260 22201 29288
rect 21968 29248 21974 29260
rect 22189 29257 22201 29260
rect 22235 29257 22247 29291
rect 22189 29251 22247 29257
rect 12713 29155 12771 29161
rect 12713 29121 12725 29155
rect 12759 29121 12771 29155
rect 13096 29152 13124 29248
rect 14826 29180 14832 29232
rect 14884 29220 14890 29232
rect 15013 29223 15071 29229
rect 15013 29220 15025 29223
rect 14884 29192 15025 29220
rect 14884 29180 14890 29192
rect 15013 29189 15025 29192
rect 15059 29189 15071 29223
rect 15013 29183 15071 29189
rect 13173 29155 13231 29161
rect 13173 29152 13185 29155
rect 13096 29124 13185 29152
rect 12713 29115 12771 29121
rect 13173 29121 13185 29124
rect 13219 29121 13231 29155
rect 13173 29115 13231 29121
rect 12728 29084 12756 29115
rect 14642 29112 14648 29164
rect 14700 29112 14706 29164
rect 15654 29112 15660 29164
rect 15712 29112 15718 29164
rect 19334 29112 19340 29164
rect 19392 29112 19398 29164
rect 19886 29112 19892 29164
rect 19944 29112 19950 29164
rect 20806 29112 20812 29164
rect 20864 29112 20870 29164
rect 22094 29112 22100 29164
rect 22152 29112 22158 29164
rect 13262 29084 13268 29096
rect 12728 29056 13268 29084
rect 13262 29044 13268 29056
rect 13320 29044 13326 29096
rect 12526 28976 12532 29028
rect 12584 29016 12590 29028
rect 12989 29019 13047 29025
rect 12989 29016 13001 29019
rect 12584 28988 13001 29016
rect 12584 28976 12590 28988
rect 12989 28985 13001 28988
rect 13035 28985 13047 29019
rect 12989 28979 13047 28985
rect 15194 28976 15200 29028
rect 15252 28976 15258 29028
rect 1104 28858 30820 28880
rect 1104 28806 4664 28858
rect 4716 28806 4728 28858
rect 4780 28806 4792 28858
rect 4844 28806 4856 28858
rect 4908 28806 4920 28858
rect 4972 28806 12092 28858
rect 12144 28806 12156 28858
rect 12208 28806 12220 28858
rect 12272 28806 12284 28858
rect 12336 28806 12348 28858
rect 12400 28806 19520 28858
rect 19572 28806 19584 28858
rect 19636 28806 19648 28858
rect 19700 28806 19712 28858
rect 19764 28806 19776 28858
rect 19828 28806 26948 28858
rect 27000 28806 27012 28858
rect 27064 28806 27076 28858
rect 27128 28806 27140 28858
rect 27192 28806 27204 28858
rect 27256 28806 30820 28858
rect 1104 28784 30820 28806
rect 1104 28314 30820 28336
rect 1104 28262 5324 28314
rect 5376 28262 5388 28314
rect 5440 28262 5452 28314
rect 5504 28262 5516 28314
rect 5568 28262 5580 28314
rect 5632 28262 12752 28314
rect 12804 28262 12816 28314
rect 12868 28262 12880 28314
rect 12932 28262 12944 28314
rect 12996 28262 13008 28314
rect 13060 28262 20180 28314
rect 20232 28262 20244 28314
rect 20296 28262 20308 28314
rect 20360 28262 20372 28314
rect 20424 28262 20436 28314
rect 20488 28262 27608 28314
rect 27660 28262 27672 28314
rect 27724 28262 27736 28314
rect 27788 28262 27800 28314
rect 27852 28262 27864 28314
rect 27916 28262 30820 28314
rect 1104 28240 30820 28262
rect 1104 27770 30820 27792
rect 1104 27718 4664 27770
rect 4716 27718 4728 27770
rect 4780 27718 4792 27770
rect 4844 27718 4856 27770
rect 4908 27718 4920 27770
rect 4972 27718 12092 27770
rect 12144 27718 12156 27770
rect 12208 27718 12220 27770
rect 12272 27718 12284 27770
rect 12336 27718 12348 27770
rect 12400 27718 19520 27770
rect 19572 27718 19584 27770
rect 19636 27718 19648 27770
rect 19700 27718 19712 27770
rect 19764 27718 19776 27770
rect 19828 27718 26948 27770
rect 27000 27718 27012 27770
rect 27064 27718 27076 27770
rect 27128 27718 27140 27770
rect 27192 27718 27204 27770
rect 27256 27718 30820 27770
rect 1104 27696 30820 27718
rect 1104 27226 30820 27248
rect 1104 27174 5324 27226
rect 5376 27174 5388 27226
rect 5440 27174 5452 27226
rect 5504 27174 5516 27226
rect 5568 27174 5580 27226
rect 5632 27174 12752 27226
rect 12804 27174 12816 27226
rect 12868 27174 12880 27226
rect 12932 27174 12944 27226
rect 12996 27174 13008 27226
rect 13060 27174 20180 27226
rect 20232 27174 20244 27226
rect 20296 27174 20308 27226
rect 20360 27174 20372 27226
rect 20424 27174 20436 27226
rect 20488 27174 27608 27226
rect 27660 27174 27672 27226
rect 27724 27174 27736 27226
rect 27788 27174 27800 27226
rect 27852 27174 27864 27226
rect 27916 27174 30820 27226
rect 1104 27152 30820 27174
rect 1104 26682 30820 26704
rect 1104 26630 4664 26682
rect 4716 26630 4728 26682
rect 4780 26630 4792 26682
rect 4844 26630 4856 26682
rect 4908 26630 4920 26682
rect 4972 26630 12092 26682
rect 12144 26630 12156 26682
rect 12208 26630 12220 26682
rect 12272 26630 12284 26682
rect 12336 26630 12348 26682
rect 12400 26630 19520 26682
rect 19572 26630 19584 26682
rect 19636 26630 19648 26682
rect 19700 26630 19712 26682
rect 19764 26630 19776 26682
rect 19828 26630 26948 26682
rect 27000 26630 27012 26682
rect 27064 26630 27076 26682
rect 27128 26630 27140 26682
rect 27192 26630 27204 26682
rect 27256 26630 30820 26682
rect 1104 26608 30820 26630
rect 1104 26138 30820 26160
rect 1104 26086 5324 26138
rect 5376 26086 5388 26138
rect 5440 26086 5452 26138
rect 5504 26086 5516 26138
rect 5568 26086 5580 26138
rect 5632 26086 12752 26138
rect 12804 26086 12816 26138
rect 12868 26086 12880 26138
rect 12932 26086 12944 26138
rect 12996 26086 13008 26138
rect 13060 26086 20180 26138
rect 20232 26086 20244 26138
rect 20296 26086 20308 26138
rect 20360 26086 20372 26138
rect 20424 26086 20436 26138
rect 20488 26086 27608 26138
rect 27660 26086 27672 26138
rect 27724 26086 27736 26138
rect 27788 26086 27800 26138
rect 27852 26086 27864 26138
rect 27916 26086 30820 26138
rect 1104 26064 30820 26086
rect 20070 25848 20076 25900
rect 20128 25888 20134 25900
rect 21177 25891 21235 25897
rect 21177 25888 21189 25891
rect 20128 25860 21189 25888
rect 20128 25848 20134 25860
rect 21177 25857 21189 25860
rect 21223 25888 21235 25891
rect 22738 25888 22744 25900
rect 21223 25860 22744 25888
rect 21223 25857 21235 25860
rect 21177 25851 21235 25857
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 21174 25644 21180 25696
rect 21232 25684 21238 25696
rect 21269 25687 21327 25693
rect 21269 25684 21281 25687
rect 21232 25656 21281 25684
rect 21232 25644 21238 25656
rect 21269 25653 21281 25656
rect 21315 25653 21327 25687
rect 21269 25647 21327 25653
rect 1104 25594 30820 25616
rect 1104 25542 4664 25594
rect 4716 25542 4728 25594
rect 4780 25542 4792 25594
rect 4844 25542 4856 25594
rect 4908 25542 4920 25594
rect 4972 25542 12092 25594
rect 12144 25542 12156 25594
rect 12208 25542 12220 25594
rect 12272 25542 12284 25594
rect 12336 25542 12348 25594
rect 12400 25542 19520 25594
rect 19572 25542 19584 25594
rect 19636 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 26948 25594
rect 27000 25542 27012 25594
rect 27064 25542 27076 25594
rect 27128 25542 27140 25594
rect 27192 25542 27204 25594
rect 27256 25542 30820 25594
rect 1104 25520 30820 25542
rect 18785 25483 18843 25489
rect 18785 25449 18797 25483
rect 18831 25480 18843 25483
rect 18966 25480 18972 25492
rect 18831 25452 18972 25480
rect 18831 25449 18843 25452
rect 18785 25443 18843 25449
rect 18966 25440 18972 25452
rect 19024 25440 19030 25492
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25313 14611 25347
rect 14553 25307 14611 25313
rect 14461 25279 14519 25285
rect 14461 25245 14473 25279
rect 14507 25245 14519 25279
rect 14568 25276 14596 25307
rect 14734 25304 14740 25356
rect 14792 25344 14798 25356
rect 14829 25347 14887 25353
rect 14829 25344 14841 25347
rect 14792 25316 14841 25344
rect 14792 25304 14798 25316
rect 14829 25313 14841 25316
rect 14875 25313 14887 25347
rect 14829 25307 14887 25313
rect 18414 25304 18420 25356
rect 18472 25344 18478 25356
rect 20165 25347 20223 25353
rect 20165 25344 20177 25347
rect 18472 25316 20177 25344
rect 18472 25304 18478 25316
rect 20165 25313 20177 25316
rect 20211 25344 20223 25347
rect 20211 25316 24164 25344
rect 20211 25313 20223 25316
rect 20165 25307 20223 25313
rect 14918 25276 14924 25288
rect 14568 25248 14924 25276
rect 14461 25239 14519 25245
rect 14476 25208 14504 25239
rect 14918 25236 14924 25248
rect 14976 25236 14982 25288
rect 15841 25279 15899 25285
rect 15841 25245 15853 25279
rect 15887 25245 15899 25279
rect 15841 25239 15899 25245
rect 14826 25208 14832 25220
rect 14476 25180 14832 25208
rect 14826 25168 14832 25180
rect 14884 25168 14890 25220
rect 15856 25208 15884 25239
rect 15930 25236 15936 25288
rect 15988 25236 15994 25288
rect 18877 25279 18935 25285
rect 18877 25276 18889 25279
rect 18800 25248 18889 25276
rect 15856 25180 16068 25208
rect 16040 25152 16068 25180
rect 16206 25168 16212 25220
rect 16264 25168 16270 25220
rect 17218 25168 17224 25220
rect 17276 25168 17282 25220
rect 17862 25168 17868 25220
rect 17920 25208 17926 25220
rect 17957 25211 18015 25217
rect 17957 25208 17969 25211
rect 17920 25180 17969 25208
rect 17920 25168 17926 25180
rect 17957 25177 17969 25180
rect 18003 25177 18015 25211
rect 17957 25171 18015 25177
rect 18800 25152 18828 25248
rect 18877 25245 18889 25248
rect 18923 25245 18935 25279
rect 18877 25239 18935 25245
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25276 19395 25279
rect 20070 25276 20076 25288
rect 19383 25248 20076 25276
rect 19383 25245 19395 25248
rect 19337 25239 19395 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 24136 25285 24164 25316
rect 24210 25304 24216 25356
rect 24268 25344 24274 25356
rect 26421 25347 26479 25353
rect 26421 25344 26433 25347
rect 24268 25316 26433 25344
rect 24268 25304 24274 25316
rect 26421 25313 26433 25316
rect 26467 25313 26479 25347
rect 26421 25307 26479 25313
rect 24121 25279 24179 25285
rect 24121 25245 24133 25279
rect 24167 25276 24179 25279
rect 24397 25279 24455 25285
rect 24397 25276 24409 25279
rect 24167 25248 24409 25276
rect 24167 25245 24179 25248
rect 24121 25239 24179 25245
rect 24397 25245 24409 25248
rect 24443 25245 24455 25279
rect 24397 25239 24455 25245
rect 20441 25211 20499 25217
rect 20441 25177 20453 25211
rect 20487 25208 20499 25211
rect 20530 25208 20536 25220
rect 20487 25180 20536 25208
rect 20487 25177 20499 25180
rect 20441 25171 20499 25177
rect 20530 25168 20536 25180
rect 20588 25168 20594 25220
rect 21174 25168 21180 25220
rect 21232 25168 21238 25220
rect 22189 25211 22247 25217
rect 22189 25177 22201 25211
rect 22235 25177 22247 25211
rect 22189 25171 22247 25177
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 16022 25100 16028 25152
rect 16080 25100 16086 25152
rect 18138 25100 18144 25152
rect 18196 25140 18202 25152
rect 18417 25143 18475 25149
rect 18417 25140 18429 25143
rect 18196 25112 18429 25140
rect 18196 25100 18202 25112
rect 18417 25109 18429 25112
rect 18463 25109 18475 25143
rect 18417 25103 18475 25109
rect 18782 25100 18788 25152
rect 18840 25100 18846 25152
rect 19426 25100 19432 25152
rect 19484 25100 19490 25152
rect 21358 25100 21364 25152
rect 21416 25140 21422 25152
rect 22204 25140 22232 25171
rect 22830 25168 22836 25220
rect 22888 25168 22894 25220
rect 23845 25211 23903 25217
rect 23845 25177 23857 25211
rect 23891 25177 23903 25211
rect 23845 25171 23903 25177
rect 21416 25112 22232 25140
rect 21416 25100 21422 25112
rect 22278 25100 22284 25152
rect 22336 25140 22342 25152
rect 22373 25143 22431 25149
rect 22373 25140 22385 25143
rect 22336 25112 22385 25140
rect 22336 25100 22342 25112
rect 22373 25109 22385 25112
rect 22419 25109 22431 25143
rect 22373 25103 22431 25109
rect 22554 25100 22560 25152
rect 22612 25140 22618 25152
rect 23860 25140 23888 25171
rect 22612 25112 23888 25140
rect 24412 25140 24440 25239
rect 24670 25168 24676 25220
rect 24728 25168 24734 25220
rect 25222 25168 25228 25220
rect 25280 25168 25286 25220
rect 24854 25140 24860 25152
rect 24412 25112 24860 25140
rect 22612 25100 22618 25112
rect 24854 25100 24860 25112
rect 24912 25100 24918 25152
rect 1104 25050 30820 25072
rect 1104 24998 5324 25050
rect 5376 24998 5388 25050
rect 5440 24998 5452 25050
rect 5504 24998 5516 25050
rect 5568 24998 5580 25050
rect 5632 24998 12752 25050
rect 12804 24998 12816 25050
rect 12868 24998 12880 25050
rect 12932 24998 12944 25050
rect 12996 24998 13008 25050
rect 13060 24998 20180 25050
rect 20232 24998 20244 25050
rect 20296 24998 20308 25050
rect 20360 24998 20372 25050
rect 20424 24998 20436 25050
rect 20488 24998 27608 25050
rect 27660 24998 27672 25050
rect 27724 24998 27736 25050
rect 27788 24998 27800 25050
rect 27852 24998 27864 25050
rect 27916 24998 30820 25050
rect 1104 24976 30820 24998
rect 17218 24896 17224 24948
rect 17276 24896 17282 24948
rect 20257 24939 20315 24945
rect 20257 24905 20269 24939
rect 20303 24936 20315 24939
rect 20530 24936 20536 24948
rect 20303 24908 20536 24936
rect 20303 24905 20315 24908
rect 20257 24899 20315 24905
rect 20530 24896 20536 24908
rect 20588 24896 20594 24948
rect 22005 24939 22063 24945
rect 22005 24905 22017 24939
rect 22051 24936 22063 24939
rect 22554 24936 22560 24948
rect 22051 24908 22560 24936
rect 22051 24905 22063 24908
rect 22005 24899 22063 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 22830 24896 22836 24948
rect 22888 24936 22894 24948
rect 22925 24939 22983 24945
rect 22925 24936 22937 24939
rect 22888 24908 22937 24936
rect 22888 24896 22894 24908
rect 22925 24905 22937 24908
rect 22971 24905 22983 24939
rect 22925 24899 22983 24905
rect 24397 24939 24455 24945
rect 24397 24905 24409 24939
rect 24443 24936 24455 24939
rect 24670 24936 24676 24948
rect 24443 24908 24676 24936
rect 24443 24905 24455 24908
rect 24397 24899 24455 24905
rect 24670 24896 24676 24908
rect 24728 24896 24734 24948
rect 25222 24896 25228 24948
rect 25280 24896 25286 24948
rect 14734 24828 14740 24880
rect 14792 24828 14798 24880
rect 15746 24828 15752 24880
rect 15804 24828 15810 24880
rect 19426 24828 19432 24880
rect 19484 24828 19490 24880
rect 20548 24840 21404 24868
rect 14182 24800 14188 24812
rect 13754 24772 14188 24800
rect 14182 24760 14188 24772
rect 14240 24760 14246 24812
rect 16022 24760 16028 24812
rect 16080 24800 16086 24812
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 16080 24772 17325 24800
rect 16080 24760 16086 24772
rect 17313 24769 17325 24772
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 18138 24760 18144 24812
rect 18196 24760 18202 24812
rect 18322 24760 18328 24812
rect 18380 24760 18386 24812
rect 20548 24809 20576 24840
rect 21376 24812 21404 24840
rect 22296 24840 22968 24868
rect 20441 24803 20499 24809
rect 20441 24769 20453 24803
rect 20487 24769 20499 24803
rect 20441 24763 20499 24769
rect 20533 24803 20591 24809
rect 20533 24769 20545 24803
rect 20579 24769 20591 24803
rect 20533 24763 20591 24769
rect 12345 24735 12403 24741
rect 12345 24701 12357 24735
rect 12391 24701 12403 24735
rect 12345 24695 12403 24701
rect 12360 24596 12388 24695
rect 12618 24692 12624 24744
rect 12676 24692 12682 24744
rect 14366 24692 14372 24744
rect 14424 24692 14430 24744
rect 14458 24692 14464 24744
rect 14516 24732 14522 24744
rect 15930 24732 15936 24744
rect 14516 24704 15936 24732
rect 14516 24692 14522 24704
rect 15930 24692 15936 24704
rect 15988 24692 15994 24744
rect 14476 24596 14504 24692
rect 12360 24568 14504 24596
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 16040 24596 16068 24760
rect 16114 24692 16120 24744
rect 16172 24732 16178 24744
rect 16485 24735 16543 24741
rect 16485 24732 16497 24735
rect 16172 24704 16497 24732
rect 16172 24692 16178 24704
rect 16485 24701 16497 24704
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 14608 24568 16068 24596
rect 14608 24556 14614 24568
rect 17954 24556 17960 24608
rect 18012 24556 18018 24608
rect 18156 24596 18184 24760
rect 18414 24692 18420 24744
rect 18472 24692 18478 24744
rect 18690 24692 18696 24744
rect 18748 24692 18754 24744
rect 20456 24732 20484 24763
rect 20622 24760 20628 24812
rect 20680 24760 20686 24812
rect 20809 24803 20867 24809
rect 20809 24769 20821 24803
rect 20855 24769 20867 24803
rect 20809 24763 20867 24769
rect 20456 24704 20576 24732
rect 20548 24664 20576 24704
rect 20714 24692 20720 24744
rect 20772 24732 20778 24744
rect 20824 24732 20852 24763
rect 21358 24760 21364 24812
rect 21416 24760 21422 24812
rect 21818 24760 21824 24812
rect 21876 24800 21882 24812
rect 22296 24809 22324 24840
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 21876 24772 22201 24800
rect 21876 24760 21882 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 22281 24803 22339 24809
rect 22281 24769 22293 24803
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 22296 24732 22324 24763
rect 22370 24760 22376 24812
rect 22428 24760 22434 24812
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 20772 24704 22324 24732
rect 22572 24732 22600 24763
rect 22830 24760 22836 24812
rect 22888 24760 22894 24812
rect 22940 24800 22968 24840
rect 23952 24840 24348 24868
rect 23845 24803 23903 24809
rect 23845 24800 23857 24803
rect 22940 24772 23857 24800
rect 23845 24769 23857 24772
rect 23891 24800 23903 24803
rect 23952 24800 23980 24840
rect 23891 24772 23980 24800
rect 24029 24803 24087 24809
rect 23891 24769 23903 24772
rect 23845 24763 23903 24769
rect 24029 24769 24041 24803
rect 24075 24769 24087 24803
rect 24029 24763 24087 24769
rect 23109 24735 23167 24741
rect 23109 24732 23121 24735
rect 22572 24704 23121 24732
rect 20772 24692 20778 24704
rect 23109 24701 23121 24704
rect 23155 24701 23167 24735
rect 23109 24695 23167 24701
rect 23198 24692 23204 24744
rect 23256 24732 23262 24744
rect 23661 24735 23719 24741
rect 23661 24732 23673 24735
rect 23256 24704 23673 24732
rect 23256 24692 23262 24704
rect 23661 24701 23673 24704
rect 23707 24701 23719 24735
rect 23661 24695 23719 24701
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 24044 24732 24072 24763
rect 24118 24760 24124 24812
rect 24176 24760 24182 24812
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 23808 24704 24072 24732
rect 23808 24692 23814 24704
rect 19720 24636 23336 24664
rect 19720 24596 19748 24636
rect 23308 24608 23336 24636
rect 18156 24568 19748 24596
rect 19978 24556 19984 24608
rect 20036 24596 20042 24608
rect 20165 24599 20223 24605
rect 20165 24596 20177 24599
rect 20036 24568 20177 24596
rect 20036 24556 20042 24568
rect 20165 24565 20177 24568
rect 20211 24565 20223 24599
rect 20165 24559 20223 24565
rect 20438 24556 20444 24608
rect 20496 24596 20502 24608
rect 21910 24596 21916 24608
rect 20496 24568 21916 24596
rect 20496 24556 20502 24568
rect 21910 24556 21916 24568
rect 21968 24556 21974 24608
rect 22278 24556 22284 24608
rect 22336 24596 22342 24608
rect 23198 24596 23204 24608
rect 22336 24568 23204 24596
rect 22336 24556 22342 24568
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23290 24556 23296 24608
rect 23348 24596 23354 24608
rect 24228 24596 24256 24763
rect 23348 24568 24256 24596
rect 24320 24596 24348 24840
rect 25130 24760 25136 24812
rect 25188 24800 25194 24812
rect 25958 24800 25964 24812
rect 25188 24772 25964 24800
rect 25188 24760 25194 24772
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 25590 24596 25596 24608
rect 24320 24568 25596 24596
rect 23348 24556 23354 24568
rect 25590 24556 25596 24568
rect 25648 24556 25654 24608
rect 1104 24506 30820 24528
rect 1104 24454 4664 24506
rect 4716 24454 4728 24506
rect 4780 24454 4792 24506
rect 4844 24454 4856 24506
rect 4908 24454 4920 24506
rect 4972 24454 12092 24506
rect 12144 24454 12156 24506
rect 12208 24454 12220 24506
rect 12272 24454 12284 24506
rect 12336 24454 12348 24506
rect 12400 24454 19520 24506
rect 19572 24454 19584 24506
rect 19636 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 26948 24506
rect 27000 24454 27012 24506
rect 27064 24454 27076 24506
rect 27128 24454 27140 24506
rect 27192 24454 27204 24506
rect 27256 24454 30820 24506
rect 1104 24432 30820 24454
rect 12618 24352 12624 24404
rect 12676 24392 12682 24404
rect 13173 24395 13231 24401
rect 13173 24392 13185 24395
rect 12676 24364 13185 24392
rect 12676 24352 12682 24364
rect 13173 24361 13185 24364
rect 13219 24361 13231 24395
rect 13173 24355 13231 24361
rect 14182 24352 14188 24404
rect 14240 24352 14246 24404
rect 14458 24352 14464 24404
rect 14516 24352 14522 24404
rect 16117 24395 16175 24401
rect 16117 24361 16129 24395
rect 16163 24392 16175 24395
rect 16206 24392 16212 24404
rect 16163 24364 16212 24392
rect 16163 24361 16175 24364
rect 16117 24355 16175 24361
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 17681 24395 17739 24401
rect 17681 24392 17693 24395
rect 17420 24364 17693 24392
rect 13081 24327 13139 24333
rect 13081 24293 13093 24327
rect 13127 24324 13139 24327
rect 14476 24324 14504 24352
rect 13127 24296 14504 24324
rect 13127 24293 13139 24296
rect 13081 24287 13139 24293
rect 15381 24259 15439 24265
rect 15381 24256 15393 24259
rect 13372 24228 15393 24256
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24188 12955 24191
rect 13078 24188 13084 24200
rect 12943 24160 13084 24188
rect 12943 24157 12955 24160
rect 12897 24151 12955 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13372 24197 13400 24228
rect 15381 24225 15393 24228
rect 15427 24225 15439 24259
rect 17420 24256 17448 24364
rect 17681 24361 17693 24364
rect 17727 24361 17739 24395
rect 17681 24355 17739 24361
rect 17954 24352 17960 24404
rect 18012 24352 18018 24404
rect 18690 24352 18696 24404
rect 18748 24392 18754 24404
rect 19061 24395 19119 24401
rect 19061 24392 19073 24395
rect 18748 24364 19073 24392
rect 18748 24352 18754 24364
rect 19061 24361 19073 24364
rect 19107 24361 19119 24395
rect 19061 24355 19119 24361
rect 20070 24352 20076 24404
rect 20128 24392 20134 24404
rect 20257 24395 20315 24401
rect 20257 24392 20269 24395
rect 20128 24364 20269 24392
rect 20128 24352 20134 24364
rect 20257 24361 20269 24364
rect 20303 24361 20315 24395
rect 20257 24355 20315 24361
rect 20533 24395 20591 24401
rect 20533 24361 20545 24395
rect 20579 24392 20591 24395
rect 20622 24392 20628 24404
rect 20579 24364 20628 24392
rect 20579 24361 20591 24364
rect 20533 24355 20591 24361
rect 20622 24352 20628 24364
rect 20680 24352 20686 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 20732 24364 21189 24392
rect 15381 24219 15439 24225
rect 17328 24228 17448 24256
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24157 13415 24191
rect 13357 24151 13415 24157
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 14292 24120 14320 24151
rect 14366 24148 14372 24200
rect 14424 24188 14430 24200
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14424 24160 14473 24188
rect 14424 24148 14430 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14826 24148 14832 24200
rect 14884 24148 14890 24200
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 14976 24160 16037 24188
rect 14976 24148 14982 24160
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17218 24188 17224 24200
rect 17083 24160 17224 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 14550 24120 14556 24132
rect 14292 24092 14556 24120
rect 14292 24064 14320 24092
rect 14550 24080 14556 24092
rect 14608 24080 14614 24132
rect 15013 24123 15071 24129
rect 15013 24120 15025 24123
rect 14752 24092 15025 24120
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14752 24061 14780 24092
rect 15013 24089 15025 24092
rect 15059 24089 15071 24123
rect 15013 24083 15071 24089
rect 15197 24123 15255 24129
rect 15197 24089 15209 24123
rect 15243 24120 15255 24123
rect 15378 24120 15384 24132
rect 15243 24092 15384 24120
rect 15243 24089 15255 24092
rect 15197 24083 15255 24089
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 14737 24055 14795 24061
rect 14737 24021 14749 24055
rect 14783 24021 14795 24055
rect 16040 24052 16068 24151
rect 17218 24148 17224 24160
rect 17276 24148 17282 24200
rect 17328 24197 17356 24228
rect 17494 24216 17500 24268
rect 17552 24256 17558 24268
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 17552 24228 17785 24256
rect 17552 24216 17558 24228
rect 17773 24225 17785 24228
rect 17819 24225 17831 24259
rect 17773 24219 17831 24225
rect 17862 24216 17868 24268
rect 17920 24216 17926 24268
rect 17972 24256 18000 24352
rect 18049 24327 18107 24333
rect 18049 24293 18061 24327
rect 18095 24324 18107 24327
rect 18598 24324 18604 24336
rect 18095 24296 18604 24324
rect 18095 24293 18107 24296
rect 18049 24287 18107 24293
rect 18598 24284 18604 24296
rect 18656 24324 18662 24336
rect 20438 24324 20444 24336
rect 18656 24296 20444 24324
rect 18656 24284 18662 24296
rect 20438 24284 20444 24296
rect 20496 24284 20502 24336
rect 20622 24256 20628 24268
rect 17972 24228 18736 24256
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17405 24191 17463 24197
rect 17405 24157 17417 24191
rect 17451 24188 17463 24191
rect 17681 24191 17739 24197
rect 17681 24188 17693 24191
rect 17451 24160 17693 24188
rect 17451 24157 17463 24160
rect 17405 24151 17463 24157
rect 17681 24157 17693 24160
rect 17727 24188 17739 24191
rect 17880 24188 17908 24216
rect 17727 24160 17908 24188
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 16114 24080 16120 24132
rect 16172 24120 16178 24132
rect 17328 24120 17356 24151
rect 16172 24092 17356 24120
rect 16172 24080 16178 24092
rect 16942 24052 16948 24064
rect 16040 24024 16948 24052
rect 14737 24015 14795 24021
rect 16942 24012 16948 24024
rect 17000 24052 17006 24064
rect 17420 24052 17448 24151
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 18708 24197 18736 24228
rect 19306 24228 20628 24256
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 18138 24080 18144 24132
rect 18196 24120 18202 24132
rect 18782 24120 18788 24132
rect 18196 24092 18788 24120
rect 18196 24080 18202 24092
rect 18782 24080 18788 24092
rect 18840 24120 18846 24132
rect 19306 24120 19334 24228
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 20732 24265 20760 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 21818 24352 21824 24404
rect 21876 24352 21882 24404
rect 21910 24352 21916 24404
rect 21968 24392 21974 24404
rect 22051 24395 22109 24401
rect 22051 24392 22063 24395
rect 21968 24364 22063 24392
rect 21968 24352 21974 24364
rect 22051 24361 22063 24364
rect 22097 24361 22109 24395
rect 22051 24355 22109 24361
rect 22066 24324 22094 24355
rect 22370 24352 22376 24404
rect 22428 24392 22434 24404
rect 22649 24395 22707 24401
rect 22649 24392 22661 24395
rect 22428 24364 22661 24392
rect 22428 24352 22434 24364
rect 22649 24361 22661 24364
rect 22695 24361 22707 24395
rect 22649 24355 22707 24361
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 22888 24364 23796 24392
rect 22888 24352 22894 24364
rect 23385 24327 23443 24333
rect 22066 24296 23244 24324
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24225 20775 24259
rect 20717 24219 20775 24225
rect 20809 24259 20867 24265
rect 20809 24225 20821 24259
rect 20855 24225 20867 24259
rect 20809 24219 20867 24225
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20441 24191 20499 24197
rect 20441 24188 20453 24191
rect 20036 24160 20453 24188
rect 20036 24148 20042 24160
rect 20441 24157 20453 24160
rect 20487 24157 20499 24191
rect 20824 24190 20852 24219
rect 20898 24216 20904 24268
rect 20956 24256 20962 24268
rect 20956 24228 21001 24256
rect 20956 24216 20962 24228
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 21913 24259 21971 24265
rect 21913 24256 21925 24259
rect 21140 24228 21925 24256
rect 21140 24216 21146 24228
rect 21913 24225 21925 24228
rect 21959 24256 21971 24259
rect 21959 24228 23152 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 20441 24151 20499 24157
rect 20732 24162 20852 24190
rect 20994 24191 21052 24197
rect 20732 24132 20760 24162
rect 20994 24157 21006 24191
rect 21040 24157 21052 24191
rect 20994 24151 21052 24157
rect 18840 24092 19334 24120
rect 18840 24080 18846 24092
rect 20714 24080 20720 24132
rect 20772 24080 20778 24132
rect 21013 24120 21041 24151
rect 21726 24148 21732 24200
rect 21784 24148 21790 24200
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22278 24188 22284 24200
rect 22235 24160 22284 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 23124 24197 23152 24228
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24157 23167 24191
rect 23216 24188 23244 24296
rect 23385 24293 23397 24327
rect 23431 24324 23443 24327
rect 23658 24324 23664 24336
rect 23431 24296 23664 24324
rect 23431 24293 23443 24296
rect 23385 24287 23443 24293
rect 23658 24284 23664 24296
rect 23716 24284 23722 24336
rect 23768 24324 23796 24364
rect 25130 24324 25136 24336
rect 23768 24296 25136 24324
rect 25130 24284 25136 24296
rect 25188 24284 25194 24336
rect 25498 24256 25504 24268
rect 24596 24228 25504 24256
rect 24596 24197 24624 24228
rect 25498 24216 25504 24228
rect 25556 24216 25562 24268
rect 23385 24191 23443 24197
rect 23385 24188 23397 24191
rect 23216 24160 23397 24188
rect 23109 24151 23167 24157
rect 23385 24157 23397 24160
rect 23431 24157 23443 24191
rect 23385 24151 23443 24157
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24157 23719 24191
rect 23661 24151 23719 24157
rect 24581 24191 24639 24197
rect 24581 24157 24593 24191
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24188 24915 24191
rect 24946 24188 24952 24200
rect 24903 24160 24952 24188
rect 24903 24157 24915 24160
rect 24857 24151 24915 24157
rect 21266 24120 21272 24132
rect 21013 24092 21272 24120
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 21358 24080 21364 24132
rect 21416 24080 21422 24132
rect 21450 24080 21456 24132
rect 21508 24120 21514 24132
rect 21545 24123 21603 24129
rect 21545 24120 21557 24123
rect 21508 24092 21557 24120
rect 21508 24080 21514 24092
rect 21545 24089 21557 24092
rect 21591 24089 21603 24123
rect 22848 24120 22876 24151
rect 23290 24120 23296 24132
rect 22848 24092 23296 24120
rect 21545 24083 21603 24089
rect 23290 24080 23296 24092
rect 23348 24080 23354 24132
rect 23676 24120 23704 24151
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25133 24191 25191 24197
rect 25133 24157 25145 24191
rect 25179 24157 25191 24191
rect 25133 24151 25191 24157
rect 25148 24120 25176 24151
rect 23400 24092 23704 24120
rect 24872 24092 25176 24120
rect 25409 24123 25467 24129
rect 23400 24064 23428 24092
rect 24872 24064 24900 24092
rect 25409 24089 25421 24123
rect 25455 24089 25467 24123
rect 25409 24083 25467 24089
rect 17000 24024 17448 24052
rect 17000 24012 17006 24024
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 20990 24052 20996 24064
rect 17552 24024 20996 24052
rect 17552 24012 17558 24024
rect 20990 24012 20996 24024
rect 21048 24052 21054 24064
rect 23014 24052 23020 24064
rect 21048 24024 23020 24052
rect 21048 24012 21054 24024
rect 23014 24012 23020 24024
rect 23072 24012 23078 24064
rect 23382 24012 23388 24064
rect 23440 24012 23446 24064
rect 23474 24012 23480 24064
rect 23532 24052 23538 24064
rect 23569 24055 23627 24061
rect 23569 24052 23581 24055
rect 23532 24024 23581 24052
rect 23532 24012 23538 24024
rect 23569 24021 23581 24024
rect 23615 24052 23627 24055
rect 24118 24052 24124 24064
rect 23615 24024 24124 24052
rect 23615 24021 23627 24024
rect 23569 24015 23627 24021
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24486 24012 24492 24064
rect 24544 24012 24550 24064
rect 24854 24012 24860 24064
rect 24912 24012 24918 24064
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25424 24052 25452 24083
rect 26050 24080 26056 24132
rect 26108 24080 26114 24132
rect 25087 24024 25452 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25498 24012 25504 24064
rect 25556 24052 25562 24064
rect 26881 24055 26939 24061
rect 26881 24052 26893 24055
rect 25556 24024 26893 24052
rect 25556 24012 25562 24024
rect 26881 24021 26893 24024
rect 26927 24021 26939 24055
rect 26881 24015 26939 24021
rect 1104 23962 30820 23984
rect 1104 23910 5324 23962
rect 5376 23910 5388 23962
rect 5440 23910 5452 23962
rect 5504 23910 5516 23962
rect 5568 23910 5580 23962
rect 5632 23910 12752 23962
rect 12804 23910 12816 23962
rect 12868 23910 12880 23962
rect 12932 23910 12944 23962
rect 12996 23910 13008 23962
rect 13060 23910 20180 23962
rect 20232 23910 20244 23962
rect 20296 23910 20308 23962
rect 20360 23910 20372 23962
rect 20424 23910 20436 23962
rect 20488 23910 27608 23962
rect 27660 23910 27672 23962
rect 27724 23910 27736 23962
rect 27788 23910 27800 23962
rect 27852 23910 27864 23962
rect 27916 23910 30820 23962
rect 1104 23888 30820 23910
rect 12989 23851 13047 23857
rect 12989 23817 13001 23851
rect 13035 23848 13047 23851
rect 13078 23848 13084 23860
rect 13035 23820 13084 23848
rect 13035 23817 13047 23820
rect 12989 23811 13047 23817
rect 13078 23808 13084 23820
rect 13136 23808 13142 23860
rect 15010 23808 15016 23860
rect 15068 23848 15074 23860
rect 15197 23851 15255 23857
rect 15197 23848 15209 23851
rect 15068 23820 15209 23848
rect 15068 23808 15074 23820
rect 15197 23817 15209 23820
rect 15243 23817 15255 23851
rect 15197 23811 15255 23817
rect 15378 23808 15384 23860
rect 15436 23808 15442 23860
rect 17037 23851 17095 23857
rect 17037 23817 17049 23851
rect 17083 23848 17095 23851
rect 17218 23848 17224 23860
rect 17083 23820 17224 23848
rect 17083 23817 17095 23820
rect 17037 23811 17095 23817
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 17494 23808 17500 23860
rect 17552 23808 17558 23860
rect 18138 23808 18144 23860
rect 18196 23808 18202 23860
rect 18598 23808 18604 23860
rect 18656 23808 18662 23860
rect 18874 23808 18880 23860
rect 18932 23848 18938 23860
rect 19429 23851 19487 23857
rect 19429 23848 19441 23851
rect 18932 23820 19441 23848
rect 18932 23808 18938 23820
rect 19429 23817 19441 23820
rect 19475 23817 19487 23851
rect 20622 23848 20628 23860
rect 19429 23811 19487 23817
rect 19720 23820 20628 23848
rect 11974 23780 11980 23792
rect 11532 23752 11980 23780
rect 1486 23672 1492 23724
rect 1544 23672 1550 23724
rect 11532 23721 11560 23752
rect 11974 23740 11980 23752
rect 12032 23740 12038 23792
rect 13449 23783 13507 23789
rect 13449 23749 13461 23783
rect 13495 23780 13507 23783
rect 13906 23780 13912 23792
rect 13495 23752 13912 23780
rect 13495 23749 13507 23752
rect 13449 23743 13507 23749
rect 13906 23740 13912 23752
rect 13964 23780 13970 23792
rect 14642 23780 14648 23792
rect 13964 23752 14648 23780
rect 13964 23740 13970 23752
rect 14642 23740 14648 23752
rect 14700 23740 14706 23792
rect 11790 23721 11796 23724
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11784 23675 11796 23721
rect 11790 23672 11796 23675
rect 11848 23672 11854 23724
rect 14366 23672 14372 23724
rect 14424 23712 14430 23724
rect 14826 23712 14832 23724
rect 14424 23684 14832 23712
rect 14424 23672 14430 23684
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 17512 23712 17540 23808
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17512 23684 17785 23712
rect 17773 23681 17785 23684
rect 17819 23681 17831 23715
rect 17773 23675 17831 23681
rect 17954 23672 17960 23724
rect 18012 23672 18018 23724
rect 18506 23672 18512 23724
rect 18564 23672 18570 23724
rect 18616 23721 18644 23808
rect 19720 23789 19748 23820
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 20714 23808 20720 23860
rect 20772 23848 20778 23860
rect 20898 23848 20904 23860
rect 20772 23820 20904 23848
rect 20772 23808 20778 23820
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 22021 23851 22079 23857
rect 22021 23848 22033 23851
rect 21008 23820 22033 23848
rect 18785 23783 18843 23789
rect 18785 23749 18797 23783
rect 18831 23780 18843 23783
rect 19705 23783 19763 23789
rect 18831 23752 19012 23780
rect 18831 23749 18843 23752
rect 18785 23743 18843 23749
rect 18984 23721 19012 23752
rect 19705 23749 19717 23783
rect 19751 23749 19763 23783
rect 19705 23743 19763 23749
rect 19978 23740 19984 23792
rect 20036 23780 20042 23792
rect 21008 23780 21036 23820
rect 22021 23817 22033 23820
rect 22067 23817 22079 23851
rect 22021 23811 22079 23817
rect 24118 23808 24124 23860
rect 24176 23848 24182 23860
rect 24176 23820 24900 23848
rect 24176 23808 24182 23820
rect 20036 23752 21036 23780
rect 21821 23783 21879 23789
rect 20036 23740 20042 23752
rect 21821 23749 21833 23783
rect 21867 23780 21879 23783
rect 22278 23780 22284 23792
rect 21867 23752 22284 23780
rect 21867 23749 21879 23752
rect 21821 23743 21879 23749
rect 22278 23740 22284 23752
rect 22336 23740 22342 23792
rect 23382 23780 23388 23792
rect 23216 23752 23388 23780
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 18969 23715 19027 23721
rect 18969 23681 18981 23715
rect 19015 23681 19027 23715
rect 18969 23675 19027 23681
rect 19153 23715 19211 23721
rect 19153 23681 19165 23715
rect 19199 23712 19211 23715
rect 19426 23712 19432 23724
rect 19199 23684 19432 23712
rect 19199 23681 19211 23684
rect 19153 23675 19211 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 19889 23715 19947 23721
rect 19889 23681 19901 23715
rect 19935 23681 19947 23715
rect 19889 23675 19947 23681
rect 20809 23715 20867 23721
rect 20809 23681 20821 23715
rect 20855 23712 20867 23715
rect 20898 23712 20904 23724
rect 20855 23684 20904 23712
rect 20855 23681 20867 23684
rect 20809 23675 20867 23681
rect 17681 23647 17739 23653
rect 17681 23644 17693 23647
rect 17236 23616 17693 23644
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23576 1731 23579
rect 6914 23576 6920 23588
rect 1719 23548 6920 23576
rect 1719 23545 1731 23548
rect 1673 23539 1731 23545
rect 6914 23536 6920 23548
rect 6972 23536 6978 23588
rect 12897 23579 12955 23585
rect 12897 23545 12909 23579
rect 12943 23576 12955 23579
rect 13173 23579 13231 23585
rect 13173 23576 13185 23579
rect 12943 23548 13185 23576
rect 12943 23545 12955 23548
rect 12897 23539 12955 23545
rect 13173 23545 13185 23548
rect 13219 23576 13231 23579
rect 13262 23576 13268 23588
rect 13219 23548 13268 23576
rect 13219 23545 13231 23548
rect 13173 23539 13231 23545
rect 13262 23536 13268 23548
rect 13320 23536 13326 23588
rect 16114 23576 16120 23588
rect 15212 23548 16120 23576
rect 14918 23468 14924 23520
rect 14976 23508 14982 23520
rect 15212 23517 15240 23548
rect 16114 23536 16120 23548
rect 16172 23576 16178 23588
rect 16669 23579 16727 23585
rect 16669 23576 16681 23579
rect 16172 23548 16681 23576
rect 16172 23536 16178 23548
rect 16669 23545 16681 23548
rect 16715 23545 16727 23579
rect 16669 23539 16727 23545
rect 15197 23511 15255 23517
rect 15197 23508 15209 23511
rect 14976 23480 15209 23508
rect 14976 23468 14982 23480
rect 15197 23477 15209 23480
rect 15243 23477 15255 23511
rect 15197 23471 15255 23477
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17037 23511 17095 23517
rect 17037 23508 17049 23511
rect 17000 23480 17049 23508
rect 17000 23468 17006 23480
rect 17037 23477 17049 23480
rect 17083 23477 17095 23511
rect 17037 23471 17095 23477
rect 17126 23468 17132 23520
rect 17184 23508 17190 23520
rect 17236 23517 17264 23616
rect 17681 23613 17693 23616
rect 17727 23613 17739 23647
rect 17681 23607 17739 23613
rect 18524 23576 18552 23672
rect 18782 23604 18788 23656
rect 18840 23604 18846 23656
rect 18874 23604 18880 23656
rect 18932 23644 18938 23656
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18932 23616 19073 23644
rect 18932 23604 18938 23616
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 19245 23647 19303 23653
rect 19245 23613 19257 23647
rect 19291 23644 19303 23647
rect 19521 23647 19579 23653
rect 19521 23644 19533 23647
rect 19291 23616 19533 23644
rect 19291 23613 19303 23616
rect 19245 23607 19303 23613
rect 19521 23613 19533 23616
rect 19567 23613 19579 23647
rect 19521 23607 19579 23613
rect 19904 23644 19932 23675
rect 20898 23672 20904 23684
rect 20956 23672 20962 23724
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21450 23712 21456 23724
rect 21039 23684 21456 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 20070 23644 20076 23656
rect 19904 23616 20076 23644
rect 19904 23576 19932 23616
rect 20070 23604 20076 23616
rect 20128 23644 20134 23656
rect 21192 23644 21220 23684
rect 21450 23672 21456 23684
rect 21508 23672 21514 23724
rect 23216 23644 23244 23752
rect 23382 23740 23388 23752
rect 23440 23780 23446 23792
rect 23440 23752 24808 23780
rect 23440 23740 23446 23752
rect 23474 23672 23480 23724
rect 23532 23672 23538 23724
rect 23658 23672 23664 23724
rect 23716 23712 23722 23724
rect 24780 23721 24808 23752
rect 24872 23721 24900 23820
rect 24946 23808 24952 23860
rect 25004 23808 25010 23860
rect 25317 23851 25375 23857
rect 25317 23817 25329 23851
rect 25363 23848 25375 23851
rect 25498 23848 25504 23860
rect 25363 23820 25504 23848
rect 25363 23817 25375 23820
rect 25317 23811 25375 23817
rect 24581 23715 24639 23721
rect 24581 23712 24593 23715
rect 23716 23684 24593 23712
rect 23716 23672 23722 23684
rect 24581 23681 24593 23684
rect 24627 23681 24639 23715
rect 24581 23675 24639 23681
rect 24765 23715 24823 23721
rect 24765 23681 24777 23715
rect 24811 23681 24823 23715
rect 24765 23675 24823 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 23293 23647 23351 23653
rect 23293 23644 23305 23647
rect 20128 23616 21220 23644
rect 20128 23604 20134 23616
rect 21192 23588 21220 23616
rect 22204 23616 23305 23644
rect 22204 23588 22232 23616
rect 23293 23613 23305 23616
rect 23339 23613 23351 23647
rect 23293 23607 23351 23613
rect 23386 23647 23444 23653
rect 23386 23613 23398 23647
rect 23432 23613 23444 23647
rect 23386 23607 23444 23613
rect 23569 23647 23627 23653
rect 23569 23613 23581 23647
rect 23615 23644 23627 23647
rect 23753 23647 23811 23653
rect 23753 23644 23765 23647
rect 23615 23616 23765 23644
rect 23615 23613 23627 23616
rect 23569 23607 23627 23613
rect 23753 23613 23765 23616
rect 23799 23613 23811 23647
rect 23753 23607 23811 23613
rect 18524 23548 19932 23576
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17184 23480 17233 23508
rect 17184 23468 17190 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 18524 23508 18552 23548
rect 21174 23536 21180 23588
rect 21232 23536 21238 23588
rect 22186 23536 22192 23588
rect 22244 23536 22250 23588
rect 23014 23536 23020 23588
rect 23072 23576 23078 23588
rect 23400 23576 23428 23607
rect 23934 23604 23940 23656
rect 23992 23604 23998 23656
rect 24026 23604 24032 23656
rect 24084 23604 24090 23656
rect 24118 23604 24124 23656
rect 24176 23604 24182 23656
rect 24213 23647 24271 23653
rect 24213 23613 24225 23647
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 23072 23548 23428 23576
rect 24228 23576 24256 23607
rect 25332 23576 25360 23811
rect 25498 23808 25504 23820
rect 25556 23808 25562 23860
rect 26050 23808 26056 23860
rect 26108 23808 26114 23860
rect 25958 23672 25964 23724
rect 26016 23672 26022 23724
rect 30282 23672 30288 23724
rect 30340 23712 30346 23724
rect 30377 23715 30435 23721
rect 30377 23712 30389 23715
rect 30340 23684 30389 23712
rect 30340 23672 30346 23684
rect 30377 23681 30389 23684
rect 30423 23681 30435 23715
rect 30377 23675 30435 23681
rect 25406 23604 25412 23656
rect 25464 23604 25470 23656
rect 25590 23604 25596 23656
rect 25648 23604 25654 23656
rect 24228 23548 25360 23576
rect 23072 23536 23078 23548
rect 26050 23536 26056 23588
rect 26108 23576 26114 23588
rect 30193 23579 30251 23585
rect 30193 23576 30205 23579
rect 26108 23548 30205 23576
rect 26108 23536 26114 23548
rect 30193 23545 30205 23548
rect 30239 23545 30251 23579
rect 30193 23539 30251 23545
rect 18598 23508 18604 23520
rect 18524 23480 18604 23508
rect 17221 23471 17279 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 20346 23468 20352 23520
rect 20404 23508 20410 23520
rect 20898 23508 20904 23520
rect 20404 23480 20904 23508
rect 20404 23468 20410 23480
rect 20898 23468 20904 23480
rect 20956 23508 20962 23520
rect 21358 23508 21364 23520
rect 20956 23480 21364 23508
rect 20956 23468 20962 23480
rect 21358 23468 21364 23480
rect 21416 23508 21422 23520
rect 21542 23508 21548 23520
rect 21416 23480 21548 23508
rect 21416 23468 21422 23480
rect 21542 23468 21548 23480
rect 21600 23508 21606 23520
rect 22005 23511 22063 23517
rect 22005 23508 22017 23511
rect 21600 23480 22017 23508
rect 21600 23468 21606 23480
rect 22005 23477 22017 23480
rect 22051 23477 22063 23511
rect 22005 23471 22063 23477
rect 23109 23511 23167 23517
rect 23109 23477 23121 23511
rect 23155 23508 23167 23511
rect 23474 23508 23480 23520
rect 23155 23480 23480 23508
rect 23155 23477 23167 23480
rect 23109 23471 23167 23477
rect 23474 23468 23480 23480
rect 23532 23468 23538 23520
rect 24118 23468 24124 23520
rect 24176 23508 24182 23520
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24176 23480 24409 23508
rect 24176 23468 24182 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 1104 23418 30820 23440
rect 1104 23366 4664 23418
rect 4716 23366 4728 23418
rect 4780 23366 4792 23418
rect 4844 23366 4856 23418
rect 4908 23366 4920 23418
rect 4972 23366 12092 23418
rect 12144 23366 12156 23418
rect 12208 23366 12220 23418
rect 12272 23366 12284 23418
rect 12336 23366 12348 23418
rect 12400 23366 19520 23418
rect 19572 23366 19584 23418
rect 19636 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 26948 23418
rect 27000 23366 27012 23418
rect 27064 23366 27076 23418
rect 27128 23366 27140 23418
rect 27192 23366 27204 23418
rect 27256 23366 30820 23418
rect 1104 23344 30820 23366
rect 11790 23264 11796 23316
rect 11848 23304 11854 23316
rect 12250 23304 12256 23316
rect 11848 23276 12256 23304
rect 11848 23264 11854 23276
rect 12250 23264 12256 23276
rect 12308 23264 12314 23316
rect 14918 23264 14924 23316
rect 14976 23264 14982 23316
rect 15749 23307 15807 23313
rect 15749 23273 15761 23307
rect 15795 23304 15807 23307
rect 16206 23304 16212 23316
rect 15795 23276 16212 23304
rect 15795 23273 15807 23276
rect 15749 23267 15807 23273
rect 11425 23239 11483 23245
rect 11425 23205 11437 23239
rect 11471 23205 11483 23239
rect 11425 23199 11483 23205
rect 10042 23128 10048 23180
rect 10100 23128 10106 23180
rect 11440 23168 11468 23199
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11440 23140 11621 23168
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 14826 23128 14832 23180
rect 14884 23128 14890 23180
rect 14936 23168 14964 23264
rect 15105 23171 15163 23177
rect 15105 23168 15117 23171
rect 14936 23140 15117 23168
rect 15105 23137 15117 23140
rect 15151 23137 15163 23171
rect 15105 23131 15163 23137
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15764 23168 15792 23267
rect 16206 23264 16212 23276
rect 16264 23264 16270 23316
rect 16298 23264 16304 23316
rect 16356 23304 16362 23316
rect 17954 23304 17960 23316
rect 16356 23276 17960 23304
rect 16356 23264 16362 23276
rect 17954 23264 17960 23276
rect 18012 23264 18018 23316
rect 22186 23264 22192 23316
rect 22244 23264 22250 23316
rect 23658 23264 23664 23316
rect 23716 23304 23722 23316
rect 23753 23307 23811 23313
rect 23753 23304 23765 23307
rect 23716 23276 23765 23304
rect 23716 23264 23722 23276
rect 23753 23273 23765 23276
rect 23799 23273 23811 23307
rect 23753 23267 23811 23273
rect 23934 23264 23940 23316
rect 23992 23264 23998 23316
rect 25225 23307 25283 23313
rect 25225 23273 25237 23307
rect 25271 23304 25283 23307
rect 25406 23304 25412 23316
rect 25271 23276 25412 23304
rect 25271 23273 25283 23276
rect 25225 23267 25283 23273
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 16114 23196 16120 23248
rect 16172 23196 16178 23248
rect 15243 23140 15792 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 11974 23060 11980 23112
rect 12032 23100 12038 23112
rect 12437 23103 12495 23109
rect 12437 23100 12449 23103
rect 12032 23072 12449 23100
rect 12032 23060 12038 23072
rect 12437 23069 12449 23072
rect 12483 23069 12495 23103
rect 14844 23100 14872 23128
rect 16132 23100 16160 23196
rect 16224 23168 16252 23264
rect 17218 23196 17224 23248
rect 17276 23196 17282 23248
rect 16485 23171 16543 23177
rect 16485 23168 16497 23171
rect 16224 23140 16497 23168
rect 16485 23137 16497 23140
rect 16531 23137 16543 23171
rect 17236 23168 17264 23196
rect 16485 23131 16543 23137
rect 16960 23140 17264 23168
rect 16960 23109 16988 23140
rect 19426 23128 19432 23180
rect 19484 23168 19490 23180
rect 19889 23171 19947 23177
rect 19889 23168 19901 23171
rect 19484 23140 19901 23168
rect 19484 23128 19490 23140
rect 19889 23137 19901 23140
rect 19935 23168 19947 23171
rect 20533 23171 20591 23177
rect 20533 23168 20545 23171
rect 19935 23140 20545 23168
rect 19935 23137 19947 23140
rect 19889 23131 19947 23137
rect 20533 23137 20545 23140
rect 20579 23137 20591 23171
rect 20533 23131 20591 23137
rect 20714 23128 20720 23180
rect 20772 23168 20778 23180
rect 22002 23168 22008 23180
rect 20772 23140 22008 23168
rect 20772 23128 20778 23140
rect 22002 23128 22008 23140
rect 22060 23128 22066 23180
rect 16577 23103 16635 23109
rect 16577 23100 16589 23103
rect 14844 23072 15792 23100
rect 16132 23072 16589 23100
rect 12437 23063 12495 23069
rect 9858 22992 9864 23044
rect 9916 23032 9922 23044
rect 10290 23035 10348 23041
rect 10290 23032 10302 23035
rect 9916 23004 10302 23032
rect 9916 22992 9922 23004
rect 10290 23001 10302 23004
rect 10336 23001 10348 23035
rect 10290 22995 10348 23001
rect 12704 23035 12762 23041
rect 12704 23001 12716 23035
rect 12750 23001 12762 23035
rect 15102 23032 15108 23044
rect 12704 22995 12762 23001
rect 13832 23004 15108 23032
rect 12618 22924 12624 22976
rect 12676 22964 12682 22976
rect 12728 22964 12756 22995
rect 13832 22973 13860 23004
rect 15102 22992 15108 23004
rect 15160 23032 15166 23044
rect 15764 23041 15792 23072
rect 16577 23069 16589 23072
rect 16623 23069 16635 23103
rect 16945 23103 17003 23109
rect 16945 23100 16957 23103
rect 16577 23063 16635 23069
rect 16684 23072 16957 23100
rect 15314 23035 15372 23041
rect 15314 23032 15326 23035
rect 15160 23004 15326 23032
rect 15160 22992 15166 23004
rect 15314 23001 15326 23004
rect 15360 23032 15372 23035
rect 15749 23035 15807 23041
rect 15360 23004 15700 23032
rect 15360 23001 15372 23004
rect 15314 22995 15372 23001
rect 12676 22936 12756 22964
rect 13817 22967 13875 22973
rect 12676 22924 12682 22936
rect 13817 22933 13829 22967
rect 13863 22933 13875 22967
rect 13817 22927 13875 22933
rect 15470 22924 15476 22976
rect 15528 22924 15534 22976
rect 15562 22924 15568 22976
rect 15620 22924 15626 22976
rect 15672 22964 15700 23004
rect 15749 23001 15761 23035
rect 15795 23032 15807 23035
rect 16684 23032 16712 23072
rect 16945 23069 16957 23072
rect 16991 23069 17003 23103
rect 16945 23063 17003 23069
rect 17034 23060 17040 23112
rect 17092 23060 17098 23112
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 20346 23100 20352 23112
rect 20027 23072 20352 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 17236 23032 17264 23063
rect 20346 23060 20352 23072
rect 20404 23060 20410 23112
rect 20438 23060 20444 23112
rect 20496 23060 20502 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 21174 23100 21180 23112
rect 20671 23072 21180 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 22204 23109 22232 23264
rect 22373 23239 22431 23245
rect 22373 23205 22385 23239
rect 22419 23236 22431 23239
rect 23382 23236 23388 23248
rect 22419 23208 23388 23236
rect 22419 23205 22431 23208
rect 22373 23199 22431 23205
rect 23382 23196 23388 23208
rect 23440 23236 23446 23248
rect 23952 23236 23980 23264
rect 23440 23208 23980 23236
rect 23440 23196 23446 23208
rect 23293 23171 23351 23177
rect 23293 23137 23305 23171
rect 23339 23168 23351 23171
rect 23339 23140 24624 23168
rect 23339 23137 23351 23140
rect 23293 23131 23351 23137
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23069 22247 23103
rect 22189 23063 22247 23069
rect 23474 23060 23480 23112
rect 23532 23100 23538 23112
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23532 23072 23581 23100
rect 23532 23060 23538 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 23661 23103 23719 23109
rect 23661 23069 23673 23103
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 15795 23004 16712 23032
rect 16776 23004 17264 23032
rect 17405 23035 17463 23041
rect 15795 23001 15807 23004
rect 15749 22995 15807 23001
rect 16298 22964 16304 22976
rect 15672 22936 16304 22964
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 16482 22924 16488 22976
rect 16540 22964 16546 22976
rect 16776 22964 16804 23004
rect 17405 23001 17417 23035
rect 17451 23032 17463 23035
rect 18966 23032 18972 23044
rect 17451 23004 18972 23032
rect 17451 23001 17463 23004
rect 17405 22995 17463 23001
rect 18966 22992 18972 23004
rect 19024 23032 19030 23044
rect 23676 23032 23704 23063
rect 23842 23060 23848 23112
rect 23900 23060 23906 23112
rect 24029 23103 24087 23109
rect 24029 23069 24041 23103
rect 24075 23100 24087 23103
rect 24486 23100 24492 23112
rect 24075 23072 24492 23100
rect 24075 23069 24087 23072
rect 24029 23063 24087 23069
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 24596 23109 24624 23140
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23069 24639 23103
rect 24581 23063 24639 23069
rect 24729 23103 24787 23109
rect 24729 23069 24741 23103
rect 24775 23100 24787 23103
rect 25087 23103 25145 23109
rect 24775 23069 24808 23100
rect 24729 23063 24808 23069
rect 25087 23069 25099 23103
rect 25133 23100 25145 23103
rect 25866 23100 25872 23112
rect 25133 23072 25872 23100
rect 25133 23069 25145 23072
rect 25087 23063 25145 23069
rect 19024 23004 23704 23032
rect 19024 22992 19030 23004
rect 16540 22936 16804 22964
rect 16853 22967 16911 22973
rect 16540 22924 16546 22936
rect 16853 22933 16865 22967
rect 16899 22964 16911 22967
rect 18690 22964 18696 22976
rect 16899 22936 18696 22964
rect 16899 22933 16911 22936
rect 16853 22927 16911 22933
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 20349 22967 20407 22973
rect 20349 22933 20361 22967
rect 20395 22964 20407 22967
rect 20530 22964 20536 22976
rect 20395 22936 20536 22964
rect 20395 22933 20407 22936
rect 20349 22927 20407 22933
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 21082 22924 21088 22976
rect 21140 22964 21146 22976
rect 22278 22964 22284 22976
rect 21140 22936 22284 22964
rect 21140 22924 21146 22936
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 24780 22964 24808 23063
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 24854 22992 24860 23044
rect 24912 22992 24918 23044
rect 24946 22992 24952 23044
rect 25004 22992 25010 23044
rect 25590 22964 25596 22976
rect 24780 22936 25596 22964
rect 25590 22924 25596 22936
rect 25648 22924 25654 22976
rect 1104 22874 30820 22896
rect 1104 22822 5324 22874
rect 5376 22822 5388 22874
rect 5440 22822 5452 22874
rect 5504 22822 5516 22874
rect 5568 22822 5580 22874
rect 5632 22822 12752 22874
rect 12804 22822 12816 22874
rect 12868 22822 12880 22874
rect 12932 22822 12944 22874
rect 12996 22822 13008 22874
rect 13060 22822 20180 22874
rect 20232 22822 20244 22874
rect 20296 22822 20308 22874
rect 20360 22822 20372 22874
rect 20424 22822 20436 22874
rect 20488 22822 27608 22874
rect 27660 22822 27672 22874
rect 27724 22822 27736 22874
rect 27788 22822 27800 22874
rect 27852 22822 27864 22874
rect 27916 22822 30820 22874
rect 1104 22800 30820 22822
rect 12618 22720 12624 22772
rect 12676 22760 12682 22772
rect 12805 22763 12863 22769
rect 12805 22760 12817 22763
rect 12676 22732 12817 22760
rect 12676 22720 12682 22732
rect 12805 22729 12817 22732
rect 12851 22729 12863 22763
rect 12805 22723 12863 22729
rect 14826 22720 14832 22772
rect 14884 22720 14890 22772
rect 18322 22720 18328 22772
rect 18380 22760 18386 22772
rect 18509 22763 18567 22769
rect 18509 22760 18521 22763
rect 18380 22732 18521 22760
rect 18380 22720 18386 22732
rect 18509 22729 18521 22732
rect 18555 22729 18567 22763
rect 18509 22723 18567 22729
rect 12250 22652 12256 22704
rect 12308 22652 12314 22704
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 4430 22624 4436 22636
rect 1719 22596 4436 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 4430 22584 4436 22596
rect 4488 22584 4494 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 6086 22624 6092 22636
rect 5031 22596 6092 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 934 22448 940 22500
rect 992 22488 998 22500
rect 1489 22491 1547 22497
rect 1489 22488 1501 22491
rect 992 22460 1501 22488
rect 992 22448 998 22460
rect 1489 22457 1501 22460
rect 1535 22457 1547 22491
rect 4816 22488 4844 22587
rect 6086 22584 6092 22596
rect 6144 22584 6150 22636
rect 6730 22584 6736 22636
rect 6788 22584 6794 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7650 22624 7656 22636
rect 6963 22596 7656 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7650 22584 7656 22596
rect 7708 22624 7714 22636
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7708 22596 7757 22624
rect 7708 22584 7714 22596
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22593 13047 22627
rect 14844 22624 14872 22720
rect 18417 22695 18475 22701
rect 18417 22692 18429 22695
rect 18248 22664 18429 22692
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 14844 22596 15301 22624
rect 12989 22587 13047 22593
rect 15289 22593 15301 22596
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 5166 22516 5172 22568
rect 5224 22516 5230 22568
rect 6825 22559 6883 22565
rect 6825 22525 6837 22559
rect 6871 22556 6883 22559
rect 7561 22559 7619 22565
rect 7561 22556 7573 22559
rect 6871 22528 7573 22556
rect 6871 22525 6883 22528
rect 6825 22519 6883 22525
rect 7561 22525 7573 22528
rect 7607 22525 7619 22559
rect 7561 22519 7619 22525
rect 8294 22516 8300 22568
rect 8352 22516 8358 22568
rect 9950 22516 9956 22568
rect 10008 22516 10014 22568
rect 11606 22516 11612 22568
rect 11664 22516 11670 22568
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 13004 22556 13032 22587
rect 12759 22528 13032 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 13814 22516 13820 22568
rect 13872 22516 13878 22568
rect 14918 22516 14924 22568
rect 14976 22556 14982 22568
rect 15013 22559 15071 22565
rect 15013 22556 15025 22559
rect 14976 22528 15025 22556
rect 14976 22516 14982 22528
rect 15013 22525 15025 22528
rect 15059 22525 15071 22559
rect 15013 22519 15071 22525
rect 12529 22491 12587 22497
rect 12529 22488 12541 22491
rect 4816 22460 5396 22488
rect 1489 22451 1547 22457
rect 5368 22432 5396 22460
rect 12176 22460 12541 22488
rect 4893 22423 4951 22429
rect 4893 22389 4905 22423
rect 4939 22420 4951 22423
rect 5074 22420 5080 22432
rect 4939 22392 5080 22420
rect 4939 22389 4951 22392
rect 4893 22383 4951 22389
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5350 22380 5356 22432
rect 5408 22420 5414 22432
rect 5721 22423 5779 22429
rect 5721 22420 5733 22423
rect 5408 22392 5733 22420
rect 5408 22380 5414 22392
rect 5721 22389 5733 22392
rect 5767 22389 5779 22423
rect 5721 22383 5779 22389
rect 7006 22380 7012 22432
rect 7064 22380 7070 22432
rect 9398 22380 9404 22432
rect 9456 22380 9462 22432
rect 9858 22380 9864 22432
rect 9916 22420 9922 22432
rect 12176 22429 12204 22460
rect 12529 22457 12541 22460
rect 12575 22457 12587 22491
rect 18248 22488 18276 22664
rect 18417 22661 18429 22664
rect 18463 22661 18475 22695
rect 18417 22655 18475 22661
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22593 18383 22627
rect 18524 22624 18552 22723
rect 18782 22720 18788 22772
rect 18840 22760 18846 22772
rect 18877 22763 18935 22769
rect 18877 22760 18889 22763
rect 18840 22732 18889 22760
rect 18840 22720 18846 22732
rect 18877 22729 18889 22732
rect 18923 22729 18935 22763
rect 18877 22723 18935 22729
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 21177 22763 21235 22769
rect 20588 22732 20852 22760
rect 20588 22720 20594 22732
rect 18966 22652 18972 22704
rect 19024 22692 19030 22704
rect 20824 22701 20852 22732
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 21266 22760 21272 22772
rect 21223 22732 21272 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 21726 22760 21732 22772
rect 21591 22732 21732 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 22554 22720 22560 22772
rect 22612 22760 22618 22772
rect 22612 22732 25820 22760
rect 22612 22720 22618 22732
rect 20809 22695 20867 22701
rect 19024 22664 20760 22692
rect 19024 22652 19030 22664
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 18524 22596 19073 22624
rect 18325 22587 18383 22593
rect 19061 22593 19073 22596
rect 19107 22593 19119 22627
rect 19061 22587 19119 22593
rect 19153 22627 19211 22633
rect 19153 22593 19165 22627
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 18340 22556 18368 22587
rect 18598 22556 18604 22568
rect 18340 22528 18604 22556
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 18782 22516 18788 22568
rect 18840 22516 18846 22568
rect 18877 22559 18935 22565
rect 18877 22525 18889 22559
rect 18923 22525 18935 22559
rect 19168 22556 19196 22587
rect 20530 22584 20536 22636
rect 20588 22584 20594 22636
rect 20732 22633 20760 22664
rect 20809 22661 20821 22695
rect 20855 22661 20867 22695
rect 20809 22655 20867 22661
rect 20901 22695 20959 22701
rect 20901 22661 20913 22695
rect 20947 22692 20959 22695
rect 21082 22692 21088 22704
rect 20947 22664 21088 22692
rect 20947 22661 20959 22664
rect 20901 22655 20959 22661
rect 21082 22652 21088 22664
rect 21140 22652 21146 22704
rect 22373 22695 22431 22701
rect 22373 22661 22385 22695
rect 22419 22692 22431 22695
rect 22925 22695 22983 22701
rect 22925 22692 22937 22695
rect 22419 22664 22937 22692
rect 22419 22661 22431 22664
rect 22373 22655 22431 22661
rect 22925 22661 22937 22664
rect 22971 22661 22983 22695
rect 22925 22655 22983 22661
rect 23198 22652 23204 22704
rect 23256 22692 23262 22704
rect 24026 22692 24032 22704
rect 23256 22664 24032 22692
rect 23256 22652 23262 22664
rect 24026 22652 24032 22664
rect 24084 22652 24090 22704
rect 25792 22692 25820 22732
rect 25866 22720 25872 22772
rect 25924 22720 25930 22772
rect 30193 22695 30251 22701
rect 30193 22692 30205 22695
rect 25792 22664 30205 22692
rect 30193 22661 30205 22664
rect 30239 22661 30251 22695
rect 30193 22655 30251 22661
rect 20681 22627 20760 22633
rect 20681 22593 20693 22627
rect 20727 22624 20760 22627
rect 20727 22596 20944 22624
rect 20727 22593 20739 22596
rect 20681 22587 20739 22593
rect 20916 22568 20944 22596
rect 20990 22584 20996 22636
rect 21048 22633 21054 22636
rect 21048 22587 21056 22633
rect 21048 22584 21054 22587
rect 21266 22584 21272 22636
rect 21324 22584 21330 22636
rect 21649 22633 21707 22639
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22593 21419 22627
rect 21649 22599 21661 22633
rect 21695 22630 21707 22633
rect 21695 22624 21772 22630
rect 22097 22627 22155 22633
rect 22097 22624 22109 22627
rect 21695 22602 22109 22624
rect 21695 22599 21707 22602
rect 21649 22593 21707 22599
rect 21744 22596 22109 22602
rect 22097 22593 22109 22596
rect 22143 22593 22155 22627
rect 21361 22587 21419 22593
rect 22097 22587 22155 22593
rect 18877 22519 18935 22525
rect 19076 22528 19196 22556
rect 18892 22488 18920 22519
rect 19076 22500 19104 22528
rect 20898 22516 20904 22568
rect 20956 22516 20962 22568
rect 18248 22460 18920 22488
rect 12529 22451 12587 22457
rect 12161 22423 12219 22429
rect 12161 22420 12173 22423
rect 9916 22392 12173 22420
rect 9916 22380 9922 22392
rect 12161 22389 12173 22392
rect 12207 22389 12219 22423
rect 12161 22383 12219 22389
rect 12802 22380 12808 22432
rect 12860 22420 12866 22432
rect 13265 22423 13323 22429
rect 13265 22420 13277 22423
rect 12860 22392 13277 22420
rect 12860 22380 12866 22392
rect 13265 22389 13277 22392
rect 13311 22389 13323 22423
rect 13265 22383 13323 22389
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 14737 22423 14795 22429
rect 14737 22420 14749 22423
rect 14608 22392 14749 22420
rect 14608 22380 14614 22392
rect 14737 22389 14749 22392
rect 14783 22389 14795 22423
rect 14737 22383 14795 22389
rect 15010 22380 15016 22432
rect 15068 22380 15074 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 16114 22420 16120 22432
rect 15620 22392 16120 22420
rect 15620 22380 15626 22392
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 17034 22380 17040 22432
rect 17092 22420 17098 22432
rect 17586 22420 17592 22432
rect 17092 22392 17592 22420
rect 17092 22380 17098 22392
rect 17586 22380 17592 22392
rect 17644 22380 17650 22432
rect 18892 22420 18920 22460
rect 19058 22448 19064 22500
rect 19116 22488 19122 22500
rect 21008 22488 21036 22584
rect 19116 22460 21036 22488
rect 21376 22488 21404 22587
rect 22278 22584 22284 22636
rect 22336 22584 22342 22636
rect 22465 22627 22523 22633
rect 22465 22624 22477 22627
rect 22388 22596 22477 22624
rect 21450 22516 21456 22568
rect 21508 22556 21514 22568
rect 22002 22556 22008 22568
rect 21508 22528 22008 22556
rect 21508 22516 21514 22528
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 22186 22488 22192 22500
rect 21376 22460 22192 22488
rect 19116 22448 19122 22460
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 20070 22420 20076 22432
rect 18892 22392 20076 22420
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 22388 22420 22416 22596
rect 22465 22593 22477 22596
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22554 22584 22560 22636
rect 22612 22633 22618 22636
rect 22612 22627 22641 22633
rect 22629 22624 22641 22627
rect 23017 22627 23075 22633
rect 22629 22596 22968 22624
rect 22629 22593 22641 22596
rect 22612 22587 22641 22593
rect 22612 22584 22618 22587
rect 22738 22516 22744 22568
rect 22796 22516 22802 22568
rect 22940 22556 22968 22596
rect 23017 22593 23029 22627
rect 23063 22624 23075 22627
rect 23382 22624 23388 22636
rect 23063 22596 23388 22624
rect 23063 22593 23075 22596
rect 23017 22587 23075 22593
rect 23382 22584 23388 22596
rect 23440 22584 23446 22636
rect 25409 22627 25467 22633
rect 25409 22593 25421 22627
rect 25455 22624 25467 22627
rect 25590 22624 25596 22636
rect 25455 22596 25596 22624
rect 25455 22593 25467 22596
rect 25409 22587 25467 22593
rect 25590 22584 25596 22596
rect 25648 22624 25654 22636
rect 26050 22624 26056 22636
rect 25648 22596 26056 22624
rect 25648 22584 25654 22596
rect 26050 22584 26056 22596
rect 26108 22584 26114 22636
rect 26234 22584 26240 22636
rect 26292 22584 26298 22636
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22624 30527 22627
rect 30926 22624 30932 22636
rect 30515 22596 30932 22624
rect 30515 22593 30527 22596
rect 30469 22587 30527 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 24854 22556 24860 22568
rect 22940 22528 24860 22556
rect 24854 22516 24860 22528
rect 24912 22516 24918 22568
rect 25498 22516 25504 22568
rect 25556 22516 25562 22568
rect 26145 22559 26203 22565
rect 26145 22525 26157 22559
rect 26191 22525 26203 22559
rect 26145 22519 26203 22525
rect 23198 22448 23204 22500
rect 23256 22448 23262 22500
rect 25777 22491 25835 22497
rect 25777 22457 25789 22491
rect 25823 22488 25835 22491
rect 26160 22488 26188 22519
rect 25823 22460 26188 22488
rect 25823 22457 25835 22460
rect 25777 22451 25835 22457
rect 23216 22420 23244 22448
rect 20956 22392 23244 22420
rect 20956 22380 20962 22392
rect 24026 22380 24032 22432
rect 24084 22420 24090 22432
rect 24946 22420 24952 22432
rect 24084 22392 24952 22420
rect 24084 22380 24090 22392
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 1104 22330 30820 22352
rect 1104 22278 4664 22330
rect 4716 22278 4728 22330
rect 4780 22278 4792 22330
rect 4844 22278 4856 22330
rect 4908 22278 4920 22330
rect 4972 22278 12092 22330
rect 12144 22278 12156 22330
rect 12208 22278 12220 22330
rect 12272 22278 12284 22330
rect 12336 22278 12348 22330
rect 12400 22278 19520 22330
rect 19572 22278 19584 22330
rect 19636 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 26948 22330
rect 27000 22278 27012 22330
rect 27064 22278 27076 22330
rect 27128 22278 27140 22330
rect 27192 22278 27204 22330
rect 27256 22278 30820 22330
rect 1104 22256 30820 22278
rect 5166 22176 5172 22228
rect 5224 22176 5230 22228
rect 5629 22219 5687 22225
rect 5629 22185 5641 22219
rect 5675 22216 5687 22219
rect 5718 22216 5724 22228
rect 5675 22188 5724 22216
rect 5675 22185 5687 22188
rect 5629 22179 5687 22185
rect 5718 22176 5724 22188
rect 5776 22216 5782 22228
rect 6730 22216 6736 22228
rect 5776 22188 6736 22216
rect 5776 22176 5782 22188
rect 6730 22176 6736 22188
rect 6788 22216 6794 22228
rect 9217 22219 9275 22225
rect 6788 22188 6914 22216
rect 6788 22176 6794 22188
rect 1670 21972 1676 22024
rect 1728 21972 1734 22024
rect 3786 21972 3792 22024
rect 3844 22012 3850 22024
rect 5810 22012 5816 22024
rect 3844 21984 5816 22012
rect 3844 21972 3850 21984
rect 5810 21972 5816 21984
rect 5868 21972 5874 22024
rect 6886 22012 6914 22188
rect 9217 22185 9229 22219
rect 9263 22216 9275 22219
rect 9398 22216 9404 22228
rect 9263 22188 9404 22216
rect 9263 22185 9275 22188
rect 9217 22179 9275 22185
rect 9398 22176 9404 22188
rect 9456 22176 9462 22228
rect 11606 22176 11612 22228
rect 11664 22176 11670 22228
rect 12424 22219 12482 22225
rect 12424 22185 12436 22219
rect 12470 22216 12482 22219
rect 12802 22216 12808 22228
rect 12470 22188 12808 22216
rect 12470 22185 12482 22188
rect 12424 22179 12482 22185
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 15749 22219 15807 22225
rect 15749 22185 15761 22219
rect 15795 22216 15807 22219
rect 16482 22216 16488 22228
rect 15795 22188 16488 22216
rect 15795 22185 15807 22188
rect 15749 22179 15807 22185
rect 15286 22148 15292 22160
rect 14844 22120 15292 22148
rect 7650 22040 7656 22092
rect 7708 22040 7714 22092
rect 9401 22083 9459 22089
rect 9401 22049 9413 22083
rect 9447 22080 9459 22083
rect 9493 22083 9551 22089
rect 9493 22080 9505 22083
rect 9447 22052 9505 22080
rect 9447 22049 9459 22052
rect 9401 22043 9459 22049
rect 9493 22049 9505 22052
rect 9539 22049 9551 22083
rect 9493 22043 9551 22049
rect 11974 22040 11980 22092
rect 12032 22080 12038 22092
rect 12161 22083 12219 22089
rect 12161 22080 12173 22083
rect 12032 22052 12173 22080
rect 12032 22040 12038 22052
rect 12161 22049 12173 22052
rect 12207 22049 12219 22083
rect 14737 22083 14795 22089
rect 14737 22080 14749 22083
rect 12161 22043 12219 22049
rect 14016 22052 14749 22080
rect 14016 22024 14044 22052
rect 14737 22049 14749 22052
rect 14783 22080 14795 22083
rect 14844 22080 14872 22120
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 15378 22108 15384 22160
rect 15436 22148 15442 22160
rect 15436 22120 15608 22148
rect 15436 22108 15442 22120
rect 14783 22052 14872 22080
rect 14946 22083 15004 22089
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 14946 22049 14958 22083
rect 14992 22080 15004 22083
rect 15396 22080 15424 22108
rect 14992 22052 15424 22080
rect 15473 22083 15531 22089
rect 14992 22049 15004 22052
rect 14946 22043 15004 22049
rect 15473 22049 15485 22083
rect 15519 22049 15531 22083
rect 15473 22043 15531 22049
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 6886 21984 7481 22012
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 8754 21972 8760 22024
rect 8812 21972 8818 22024
rect 8938 21972 8944 22024
rect 8996 21972 9002 22024
rect 9766 21972 9772 22024
rect 9824 22012 9830 22024
rect 9950 22012 9956 22024
rect 9824 21984 9956 22012
rect 9824 21972 9830 21984
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10229 22015 10287 22021
rect 10229 22012 10241 22015
rect 10100 21984 10241 22012
rect 10100 21972 10106 21984
rect 10229 21981 10241 21984
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 13998 21972 14004 22024
rect 14056 21972 14062 22024
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 22012 14519 22015
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 14507 21984 15393 22012
rect 14507 21981 14519 21984
rect 14461 21975 14519 21981
rect 15381 21981 15393 21984
rect 15427 21981 15439 22015
rect 15381 21975 15439 21981
rect 4056 21947 4114 21953
rect 4056 21913 4068 21947
rect 4102 21944 4114 21947
rect 4614 21944 4620 21956
rect 4102 21916 4620 21944
rect 4102 21913 4114 21916
rect 4056 21907 4114 21913
rect 4614 21904 4620 21916
rect 4672 21904 4678 21956
rect 5261 21947 5319 21953
rect 5261 21913 5273 21947
rect 5307 21944 5319 21947
rect 5350 21944 5356 21956
rect 5307 21916 5356 21944
rect 5307 21913 5319 21916
rect 5261 21907 5319 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 5445 21947 5503 21953
rect 5445 21913 5457 21947
rect 5491 21913 5503 21947
rect 5445 21907 5503 21913
rect 6080 21947 6138 21953
rect 6080 21913 6092 21947
rect 6126 21944 6138 21947
rect 6362 21944 6368 21956
rect 6126 21916 6368 21944
rect 6126 21913 6138 21916
rect 6080 21907 6138 21913
rect 934 21836 940 21888
rect 992 21876 998 21888
rect 1489 21879 1547 21885
rect 1489 21876 1501 21879
rect 992 21848 1501 21876
rect 992 21836 998 21848
rect 1489 21845 1501 21848
rect 1535 21845 1547 21879
rect 1489 21839 1547 21845
rect 5166 21836 5172 21888
rect 5224 21876 5230 21888
rect 5460 21876 5488 21907
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 7208 21916 8340 21944
rect 7208 21885 7236 21916
rect 8312 21888 8340 21916
rect 10318 21904 10324 21956
rect 10376 21944 10382 21956
rect 10474 21947 10532 21953
rect 10474 21944 10486 21947
rect 10376 21916 10486 21944
rect 10376 21904 10382 21916
rect 10474 21913 10486 21916
rect 10520 21913 10532 21947
rect 14185 21947 14243 21953
rect 14185 21944 14197 21947
rect 13662 21916 14197 21944
rect 10474 21907 10532 21913
rect 14185 21913 14197 21916
rect 14231 21913 14243 21947
rect 14185 21907 14243 21913
rect 5224 21848 5488 21876
rect 7193 21879 7251 21885
rect 5224 21836 5230 21848
rect 7193 21845 7205 21879
rect 7239 21845 7251 21879
rect 7193 21839 7251 21845
rect 7282 21836 7288 21888
rect 7340 21836 7346 21888
rect 8294 21836 8300 21888
rect 8352 21836 8358 21888
rect 8478 21836 8484 21888
rect 8536 21876 8542 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8536 21848 8585 21876
rect 8536 21836 8542 21848
rect 8573 21845 8585 21848
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 10008 21848 10149 21876
rect 10008 21836 10014 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 10137 21839 10195 21845
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14366 21876 14372 21888
rect 13964 21848 14372 21876
rect 13964 21836 13970 21848
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15105 21879 15163 21885
rect 15105 21845 15117 21879
rect 15151 21876 15163 21879
rect 15286 21876 15292 21888
rect 15151 21848 15292 21876
rect 15151 21845 15163 21848
rect 15105 21839 15163 21845
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 15396 21876 15424 21975
rect 15488 21944 15516 22043
rect 15580 22012 15608 22120
rect 16040 22021 16068 22188
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 16850 22176 16856 22228
rect 16908 22216 16914 22228
rect 17405 22219 17463 22225
rect 17405 22216 17417 22219
rect 16908 22188 17417 22216
rect 16908 22176 16914 22188
rect 17405 22185 17417 22188
rect 17451 22185 17463 22219
rect 17405 22179 17463 22185
rect 16393 22151 16451 22157
rect 16393 22117 16405 22151
rect 16439 22148 16451 22151
rect 17310 22148 17316 22160
rect 16439 22120 17316 22148
rect 16439 22117 16451 22120
rect 16393 22111 16451 22117
rect 17310 22108 17316 22120
rect 17368 22108 17374 22160
rect 16485 22083 16543 22089
rect 16485 22049 16497 22083
rect 16531 22049 16543 22083
rect 16485 22043 16543 22049
rect 16761 22083 16819 22089
rect 16761 22049 16773 22083
rect 16807 22080 16819 22083
rect 17034 22080 17040 22092
rect 16807 22052 17040 22080
rect 16807 22049 16819 22052
rect 16761 22043 16819 22049
rect 15841 22015 15899 22021
rect 15841 22012 15853 22015
rect 15580 21984 15853 22012
rect 15841 21981 15853 21984
rect 15887 21981 15899 22015
rect 15841 21975 15899 21981
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 16209 22015 16267 22021
rect 16209 21981 16221 22015
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 15488 21916 15792 21944
rect 15764 21888 15792 21916
rect 16114 21904 16120 21956
rect 16172 21904 16178 21956
rect 16224 21944 16252 21975
rect 16298 21972 16304 22024
rect 16356 22014 16362 22024
rect 16356 22012 16436 22014
rect 16500 22012 16528 22043
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 17420 22080 17448 22179
rect 17586 22176 17592 22228
rect 17644 22216 17650 22228
rect 18141 22219 18199 22225
rect 18141 22216 18153 22219
rect 17644 22188 18153 22216
rect 17644 22176 17650 22188
rect 18141 22185 18153 22188
rect 18187 22216 18199 22219
rect 18601 22219 18659 22225
rect 18601 22216 18613 22219
rect 18187 22188 18613 22216
rect 18187 22185 18199 22188
rect 18141 22179 18199 22185
rect 18601 22185 18613 22188
rect 18647 22185 18659 22219
rect 18601 22179 18659 22185
rect 18782 22176 18788 22228
rect 18840 22216 18846 22228
rect 20441 22219 20499 22225
rect 20441 22216 20453 22219
rect 18840 22188 20453 22216
rect 18840 22176 18846 22188
rect 20441 22185 20453 22188
rect 20487 22185 20499 22219
rect 20441 22179 20499 22185
rect 18325 22151 18383 22157
rect 18325 22117 18337 22151
rect 18371 22148 18383 22151
rect 19058 22148 19064 22160
rect 18371 22120 19064 22148
rect 18371 22117 18383 22120
rect 18325 22111 18383 22117
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 20456 22148 20484 22179
rect 20530 22176 20536 22228
rect 20588 22216 20594 22228
rect 20625 22219 20683 22225
rect 20625 22216 20637 22219
rect 20588 22188 20637 22216
rect 20588 22176 20594 22188
rect 20625 22185 20637 22188
rect 20671 22185 20683 22219
rect 20625 22179 20683 22185
rect 21450 22176 21456 22228
rect 21508 22176 21514 22228
rect 22278 22176 22284 22228
rect 22336 22176 22342 22228
rect 23661 22219 23719 22225
rect 23661 22185 23673 22219
rect 23707 22216 23719 22219
rect 23750 22216 23756 22228
rect 23707 22188 23756 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 23750 22176 23756 22188
rect 23808 22176 23814 22228
rect 23842 22176 23848 22228
rect 23900 22176 23906 22228
rect 21468 22148 21496 22176
rect 20456 22120 21496 22148
rect 17773 22083 17831 22089
rect 17420 22052 17632 22080
rect 16356 21986 16528 22012
rect 16356 21972 16362 21986
rect 16408 21984 16528 21986
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16632 21984 16865 22012
rect 16632 21972 16638 21984
rect 16853 21981 16865 21984
rect 16899 22012 16911 22015
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 16899 21984 17233 22012
rect 16899 21981 16911 21984
rect 16853 21975 16911 21981
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 21981 17463 22015
rect 17405 21975 17463 21981
rect 16224 21916 16620 21944
rect 15562 21876 15568 21888
rect 15396 21848 15568 21876
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 15746 21836 15752 21888
rect 15804 21836 15810 21888
rect 16592 21876 16620 21916
rect 16666 21904 16672 21956
rect 16724 21944 16730 21956
rect 16970 21947 17028 21953
rect 16970 21944 16982 21947
rect 16724 21916 16982 21944
rect 16724 21904 16730 21916
rect 16970 21913 16982 21916
rect 17016 21944 17028 21947
rect 17420 21944 17448 21975
rect 17016 21916 17448 21944
rect 17604 21944 17632 22052
rect 17773 22049 17785 22083
rect 17819 22080 17831 22083
rect 18414 22080 18420 22092
rect 17819 22052 18420 22080
rect 17819 22049 17831 22052
rect 17773 22043 17831 22049
rect 18414 22040 18420 22052
rect 18472 22040 18478 22092
rect 18690 22040 18696 22092
rect 18748 22080 18754 22092
rect 19150 22080 19156 22092
rect 18748 22052 19156 22080
rect 18748 22040 18754 22052
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 19794 22040 19800 22092
rect 19852 22080 19858 22092
rect 21269 22083 21327 22089
rect 19852 22052 20208 22080
rect 19852 22040 19858 22052
rect 20180 22024 20208 22052
rect 21269 22049 21281 22083
rect 21315 22080 21327 22083
rect 22296 22080 22324 22176
rect 21315 22052 22324 22080
rect 23109 22083 23167 22089
rect 21315 22049 21327 22052
rect 21269 22043 21327 22049
rect 23109 22049 23121 22083
rect 23155 22080 23167 22083
rect 23198 22080 23204 22092
rect 23155 22052 23204 22080
rect 23155 22049 23167 22052
rect 23109 22043 23167 22049
rect 23198 22040 23204 22052
rect 23256 22040 23262 22092
rect 23860 22080 23888 22176
rect 23768 22052 24440 22080
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18874 22012 18880 22024
rect 18288 21984 18880 22012
rect 18288 21972 18294 21984
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 20070 21972 20076 22024
rect 20128 21972 20134 22024
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 20530 22012 20536 22024
rect 20220 21984 20536 22012
rect 20220 21972 20226 21984
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 21174 21972 21180 22024
rect 21232 22012 21238 22024
rect 21453 22015 21511 22021
rect 21453 22012 21465 22015
rect 21232 21984 21465 22012
rect 21232 21972 21238 21984
rect 21453 21981 21465 21984
rect 21499 21981 21511 22015
rect 21453 21975 21511 21981
rect 21542 21972 21548 22024
rect 21600 21972 21606 22024
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21637 21975 21695 21981
rect 21729 22015 21787 22021
rect 21729 21981 21741 22015
rect 21775 22012 21787 22015
rect 22094 22012 22100 22024
rect 21775 21984 22100 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 18141 21947 18199 21953
rect 18141 21944 18153 21947
rect 17604 21916 18153 21944
rect 17016 21913 17028 21916
rect 16970 21907 17028 21913
rect 18141 21913 18153 21916
rect 18187 21913 18199 21947
rect 18141 21907 18199 21913
rect 16850 21876 16856 21888
rect 16592 21848 16856 21876
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 17129 21879 17187 21885
rect 17129 21845 17141 21879
rect 17175 21876 17187 21879
rect 18046 21876 18052 21888
rect 17175 21848 18052 21876
rect 17175 21845 17187 21848
rect 17129 21839 17187 21845
rect 18046 21836 18052 21848
rect 18104 21836 18110 21888
rect 18156 21876 18184 21907
rect 18414 21904 18420 21956
rect 18472 21904 18478 21956
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 20898 21944 20904 21956
rect 20772 21916 20904 21944
rect 20772 21904 20778 21916
rect 20898 21904 20904 21916
rect 20956 21944 20962 21956
rect 21652 21944 21680 21975
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 23440 21984 23581 22012
rect 23440 21972 23446 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23768 21944 23796 22052
rect 23842 21972 23848 22024
rect 23900 21972 23906 22024
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 22012 23995 22015
rect 24026 22012 24032 22024
rect 23983 21984 24032 22012
rect 23983 21981 23995 21984
rect 23937 21975 23995 21981
rect 24026 21972 24032 21984
rect 24084 21972 24090 22024
rect 24118 21972 24124 22024
rect 24176 21972 24182 22024
rect 24412 22021 24440 22052
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 21981 24271 22015
rect 24213 21975 24271 21981
rect 24397 22015 24455 22021
rect 24397 21981 24409 22015
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 22012 24823 22015
rect 24854 22012 24860 22024
rect 24811 21984 24860 22012
rect 24811 21981 24823 21984
rect 24765 21975 24823 21981
rect 20956 21916 21680 21944
rect 23400 21916 23796 21944
rect 20956 21904 20962 21916
rect 18617 21879 18675 21885
rect 18617 21876 18629 21879
rect 18156 21848 18629 21876
rect 18617 21845 18629 21848
rect 18663 21845 18675 21879
rect 18617 21839 18675 21845
rect 20441 21879 20499 21885
rect 20441 21845 20453 21879
rect 20487 21876 20499 21879
rect 20990 21876 20996 21888
rect 20487 21848 20996 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 20990 21836 20996 21848
rect 21048 21836 21054 21888
rect 23400 21885 23428 21916
rect 23385 21879 23443 21885
rect 23385 21845 23397 21879
rect 23431 21845 23443 21879
rect 23385 21839 23443 21845
rect 23474 21836 23480 21888
rect 23532 21836 23538 21888
rect 24228 21876 24256 21975
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 25038 21972 25044 22024
rect 25096 22012 25102 22024
rect 30193 22015 30251 22021
rect 30193 22012 30205 22015
rect 25096 21984 30205 22012
rect 25096 21972 25102 21984
rect 30193 21981 30205 21984
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 24578 21904 24584 21956
rect 24636 21904 24642 21956
rect 24673 21947 24731 21953
rect 24673 21913 24685 21947
rect 24719 21944 24731 21947
rect 26602 21944 26608 21956
rect 24719 21916 26608 21944
rect 24719 21913 24731 21916
rect 24673 21907 24731 21913
rect 26602 21904 26608 21916
rect 26660 21904 26666 21956
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24228 21848 24961 21876
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 30374 21836 30380 21888
rect 30432 21836 30438 21888
rect 1104 21786 30820 21808
rect 1104 21734 5324 21786
rect 5376 21734 5388 21786
rect 5440 21734 5452 21786
rect 5504 21734 5516 21786
rect 5568 21734 5580 21786
rect 5632 21734 12752 21786
rect 12804 21734 12816 21786
rect 12868 21734 12880 21786
rect 12932 21734 12944 21786
rect 12996 21734 13008 21786
rect 13060 21734 20180 21786
rect 20232 21734 20244 21786
rect 20296 21734 20308 21786
rect 20360 21734 20372 21786
rect 20424 21734 20436 21786
rect 20488 21734 27608 21786
rect 27660 21734 27672 21786
rect 27724 21734 27736 21786
rect 27788 21734 27800 21786
rect 27852 21734 27864 21786
rect 27916 21734 30820 21786
rect 1104 21712 30820 21734
rect 4614 21632 4620 21684
rect 4672 21632 4678 21684
rect 6362 21632 6368 21684
rect 6420 21632 6426 21684
rect 7282 21672 7288 21684
rect 6564 21644 7288 21672
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1688 21400 1716 21499
rect 5074 21496 5080 21548
rect 5132 21536 5138 21548
rect 5353 21539 5411 21545
rect 5353 21536 5365 21539
rect 5132 21508 5365 21536
rect 5132 21496 5138 21508
rect 5353 21505 5365 21508
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 5534 21496 5540 21548
rect 5592 21496 5598 21548
rect 6564 21545 6592 21644
rect 7282 21632 7288 21644
rect 7340 21632 7346 21684
rect 9585 21675 9643 21681
rect 9585 21641 9597 21675
rect 9631 21672 9643 21675
rect 9766 21672 9772 21684
rect 9631 21644 9772 21672
rect 9631 21641 9643 21644
rect 9585 21635 9643 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 10229 21675 10287 21681
rect 10229 21641 10241 21675
rect 10275 21672 10287 21675
rect 10318 21672 10324 21684
rect 10275 21644 10324 21672
rect 10275 21641 10287 21644
rect 10229 21635 10287 21641
rect 10318 21632 10324 21644
rect 10376 21632 10382 21684
rect 13633 21675 13691 21681
rect 13633 21641 13645 21675
rect 13679 21672 13691 21675
rect 13814 21672 13820 21684
rect 13679 21644 13820 21672
rect 13679 21641 13691 21644
rect 13633 21635 13691 21641
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 14826 21632 14832 21684
rect 14884 21632 14890 21684
rect 15194 21681 15200 21684
rect 15181 21675 15200 21681
rect 15181 21641 15193 21675
rect 15252 21672 15258 21684
rect 15252 21644 15608 21672
rect 15181 21635 15200 21641
rect 15194 21632 15200 21635
rect 15252 21632 15258 21644
rect 10042 21604 10048 21616
rect 6748 21576 10048 21604
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21468 5319 21471
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 5307 21440 5457 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 5445 21437 5457 21440
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 6748 21477 6776 21576
rect 7006 21545 7012 21548
rect 7000 21536 7012 21545
rect 6967 21508 7012 21536
rect 7000 21499 7012 21508
rect 7006 21496 7012 21499
rect 7064 21496 7070 21548
rect 8220 21545 8248 21576
rect 10042 21564 10048 21576
rect 10100 21564 10106 21616
rect 12434 21564 12440 21616
rect 12492 21564 12498 21616
rect 14844 21604 14872 21632
rect 13924 21576 14964 21604
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21536 8263 21539
rect 8294 21536 8300 21548
rect 8251 21508 8300 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 8294 21496 8300 21508
rect 8352 21496 8358 21548
rect 8478 21545 8484 21548
rect 8472 21499 8484 21545
rect 8478 21496 8484 21499
rect 8536 21496 8542 21548
rect 9858 21496 9864 21548
rect 9916 21496 9922 21548
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10060 21536 10088 21564
rect 11514 21536 11520 21548
rect 10060 21508 11520 21536
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 13924 21545 13952 21576
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21505 13967 21539
rect 13909 21499 13967 21505
rect 14366 21496 14372 21548
rect 14424 21536 14430 21548
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 14424 21508 14841 21536
rect 14424 21496 14430 21508
rect 14829 21505 14841 21508
rect 14875 21505 14887 21539
rect 14936 21536 14964 21576
rect 15010 21564 15016 21616
rect 15068 21604 15074 21616
rect 15381 21607 15439 21613
rect 15381 21604 15393 21607
rect 15068 21576 15393 21604
rect 15068 21564 15074 21576
rect 15381 21573 15393 21576
rect 15427 21573 15439 21607
rect 15580 21604 15608 21644
rect 15654 21632 15660 21684
rect 15712 21632 15718 21684
rect 19061 21675 19119 21681
rect 19061 21641 19073 21675
rect 19107 21672 19119 21675
rect 19886 21672 19892 21684
rect 19107 21644 19892 21672
rect 19107 21641 19119 21644
rect 19061 21635 19119 21641
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20349 21675 20407 21681
rect 20349 21672 20361 21675
rect 20220 21644 20361 21672
rect 20220 21632 20226 21644
rect 20349 21641 20361 21644
rect 20395 21672 20407 21675
rect 20395 21644 20944 21672
rect 20395 21641 20407 21644
rect 20349 21635 20407 21641
rect 16114 21604 16120 21616
rect 15580 21576 16120 21604
rect 15381 21567 15439 21573
rect 16114 21564 16120 21576
rect 16172 21564 16178 21616
rect 17310 21564 17316 21616
rect 17368 21604 17374 21616
rect 18693 21607 18751 21613
rect 18693 21604 18705 21607
rect 17368 21576 18705 21604
rect 17368 21564 17374 21576
rect 18693 21573 18705 21576
rect 18739 21573 18751 21607
rect 18693 21567 18751 21573
rect 14936 21508 15240 21536
rect 14829 21499 14887 21505
rect 6733 21471 6791 21477
rect 6733 21468 6745 21471
rect 5868 21440 6745 21468
rect 5868 21428 5874 21440
rect 6733 21437 6745 21440
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21468 9827 21471
rect 9968 21468 9996 21496
rect 9815 21440 9996 21468
rect 11793 21471 11851 21477
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 11793 21437 11805 21471
rect 11839 21468 11851 21471
rect 11882 21468 11888 21480
rect 11839 21440 11888 21468
rect 11839 21437 11851 21440
rect 11793 21431 11851 21437
rect 11882 21428 11888 21440
rect 11940 21428 11946 21480
rect 13538 21428 13544 21480
rect 13596 21428 13602 21480
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21437 13875 21471
rect 13817 21431 13875 21437
rect 6638 21400 6644 21412
rect 1688 21372 6644 21400
rect 6638 21360 6644 21372
rect 6696 21360 6702 21412
rect 13832 21400 13860 21431
rect 13998 21428 14004 21480
rect 14056 21428 14062 21480
rect 14093 21471 14151 21477
rect 14093 21437 14105 21471
rect 14139 21468 14151 21471
rect 14277 21471 14335 21477
rect 14277 21468 14289 21471
rect 14139 21440 14289 21468
rect 14139 21437 14151 21440
rect 14093 21431 14151 21437
rect 14277 21437 14289 21440
rect 14323 21437 14335 21471
rect 15212 21468 15240 21508
rect 15286 21496 15292 21548
rect 15344 21536 15350 21548
rect 15473 21539 15531 21545
rect 15473 21536 15485 21539
rect 15344 21508 15485 21536
rect 15344 21496 15350 21508
rect 15473 21505 15485 21508
rect 15519 21505 15531 21539
rect 15473 21499 15531 21505
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 15212 21440 15332 21468
rect 14277 21431 14335 21437
rect 15013 21403 15071 21409
rect 15013 21400 15025 21403
rect 13832 21372 15025 21400
rect 15013 21369 15025 21372
rect 15059 21369 15071 21403
rect 15304 21400 15332 21440
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 15746 21468 15752 21480
rect 15436 21440 15752 21468
rect 15436 21428 15442 21440
rect 15746 21428 15752 21440
rect 15804 21468 15810 21480
rect 16206 21468 16212 21480
rect 15804 21440 16212 21468
rect 15804 21428 15810 21440
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 16482 21428 16488 21480
rect 16540 21428 16546 21480
rect 15654 21400 15660 21412
rect 15304 21372 15660 21400
rect 15013 21363 15071 21369
rect 15654 21360 15660 21372
rect 15712 21400 15718 21412
rect 16298 21400 16304 21412
rect 15712 21372 16304 21400
rect 15712 21360 15718 21372
rect 16298 21360 16304 21372
rect 16356 21360 16362 21412
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1489 21335 1547 21341
rect 1489 21332 1501 21335
rect 992 21304 1501 21332
rect 992 21292 998 21304
rect 1489 21301 1501 21304
rect 1535 21301 1547 21335
rect 1489 21295 1547 21301
rect 1670 21292 1676 21344
rect 1728 21332 1734 21344
rect 6914 21332 6920 21344
rect 1728 21304 6920 21332
rect 1728 21292 1734 21304
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 8113 21335 8171 21341
rect 8113 21301 8125 21335
rect 8159 21332 8171 21335
rect 8938 21332 8944 21344
rect 8159 21304 8944 21332
rect 8159 21301 8171 21304
rect 8113 21295 8171 21301
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 15197 21335 15255 21341
rect 15197 21301 15209 21335
rect 15243 21332 15255 21335
rect 15562 21332 15568 21344
rect 15243 21304 15568 21332
rect 15243 21301 15255 21304
rect 15197 21295 15255 21301
rect 15562 21292 15568 21304
rect 15620 21332 15626 21344
rect 16500 21332 16528 21428
rect 15620 21304 16528 21332
rect 18524 21332 18552 21499
rect 18708 21468 18736 21567
rect 18782 21564 18788 21616
rect 18840 21564 18846 21616
rect 19613 21607 19671 21613
rect 19613 21573 19625 21607
rect 19659 21604 19671 21607
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 19659 21576 20085 21604
rect 19659 21573 19671 21576
rect 19613 21567 19671 21573
rect 20073 21573 20085 21576
rect 20119 21604 20131 21607
rect 20625 21607 20683 21613
rect 20625 21604 20637 21607
rect 20119 21576 20637 21604
rect 20119 21573 20131 21576
rect 20073 21567 20131 21573
rect 20625 21573 20637 21576
rect 20671 21573 20683 21607
rect 20916 21604 20944 21644
rect 20990 21632 20996 21684
rect 21048 21632 21054 21684
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 21140 21644 21189 21672
rect 21140 21632 21146 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 21266 21632 21272 21684
rect 21324 21672 21330 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21324 21644 21833 21672
rect 21324 21632 21330 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 21821 21635 21879 21641
rect 22189 21675 22247 21681
rect 22189 21641 22201 21675
rect 22235 21672 22247 21675
rect 22235 21644 22508 21672
rect 22235 21641 22247 21644
rect 22189 21635 22247 21641
rect 20916 21576 21404 21604
rect 20625 21567 20683 21573
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21536 18935 21539
rect 19150 21536 19156 21548
rect 18923 21508 19156 21536
rect 18923 21505 18935 21508
rect 18877 21499 18935 21505
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21536 19763 21539
rect 19886 21536 19892 21548
rect 19751 21508 19892 21536
rect 19751 21505 19763 21508
rect 19705 21499 19763 21505
rect 19536 21468 19564 21499
rect 19886 21496 19892 21508
rect 19944 21496 19950 21548
rect 20165 21539 20223 21545
rect 20165 21505 20177 21539
rect 20211 21536 20223 21539
rect 20346 21536 20352 21548
rect 20211 21508 20352 21536
rect 20211 21505 20223 21508
rect 20165 21499 20223 21505
rect 20346 21496 20352 21508
rect 20404 21536 20410 21548
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 20404 21508 20453 21536
rect 20404 21496 20410 21508
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 20530 21496 20536 21548
rect 20588 21536 20594 21548
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 20588 21508 20729 21536
rect 20588 21496 20594 21508
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21536 20867 21539
rect 20990 21536 20996 21548
rect 20855 21508 20996 21536
rect 20855 21505 20867 21508
rect 20809 21499 20867 21505
rect 20990 21496 20996 21508
rect 21048 21496 21054 21548
rect 21376 21545 21404 21576
rect 21542 21564 21548 21616
rect 21600 21564 21606 21616
rect 22370 21604 22376 21616
rect 22036 21576 22376 21604
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21361 21539 21419 21545
rect 21131 21508 21220 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 19978 21468 19984 21480
rect 18708 21440 19334 21468
rect 19536 21440 19984 21468
rect 18690 21332 18696 21344
rect 18524 21304 18696 21332
rect 15620 21292 15626 21304
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 19306 21332 19334 21440
rect 19978 21428 19984 21440
rect 20036 21468 20042 21480
rect 21192 21468 21220 21508
rect 21361 21505 21373 21539
rect 21407 21505 21419 21539
rect 21560 21536 21588 21564
rect 22036 21545 22064 21576
rect 22370 21564 22376 21576
rect 22428 21564 22434 21616
rect 22480 21604 22508 21644
rect 23382 21632 23388 21684
rect 23440 21672 23446 21684
rect 24121 21675 24179 21681
rect 23440 21644 23796 21672
rect 23440 21632 23446 21644
rect 22480 21576 22692 21604
rect 22664 21548 22692 21576
rect 23474 21564 23480 21616
rect 23532 21564 23538 21616
rect 23768 21613 23796 21644
rect 24121 21641 24133 21675
rect 24167 21672 24179 21675
rect 24578 21672 24584 21684
rect 24167 21644 24584 21672
rect 24167 21641 24179 21644
rect 24121 21635 24179 21641
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 25038 21632 25044 21684
rect 25096 21632 25102 21684
rect 25869 21675 25927 21681
rect 25869 21641 25881 21675
rect 25915 21672 25927 21675
rect 26234 21672 26240 21684
rect 25915 21644 26240 21672
rect 25915 21641 25927 21644
rect 25869 21635 25927 21641
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 23753 21607 23811 21613
rect 23753 21573 23765 21607
rect 23799 21573 23811 21607
rect 23753 21567 23811 21573
rect 24765 21607 24823 21613
rect 24765 21573 24777 21607
rect 24811 21604 24823 21607
rect 25314 21604 25320 21616
rect 24811 21576 25320 21604
rect 24811 21573 24823 21576
rect 24765 21567 24823 21573
rect 25314 21564 25320 21576
rect 25372 21564 25378 21616
rect 22024 21542 22082 21545
rect 21361 21499 21419 21505
rect 21468 21508 21588 21536
rect 21928 21539 22082 21542
rect 21928 21514 22036 21539
rect 21468 21468 21496 21508
rect 20036 21440 21496 21468
rect 21545 21471 21603 21477
rect 20036 21428 20042 21440
rect 21545 21437 21557 21471
rect 21591 21468 21603 21471
rect 21928 21468 21956 21514
rect 22024 21505 22036 21514
rect 22070 21505 22082 21539
rect 22024 21499 22082 21505
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21505 22339 21539
rect 22281 21499 22339 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22296 21468 22324 21499
rect 22572 21468 22600 21499
rect 22646 21496 22652 21548
rect 22704 21496 22710 21548
rect 23492 21536 23520 21564
rect 23934 21536 23940 21548
rect 23492 21508 23940 21536
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24486 21496 24492 21548
rect 24544 21496 24550 21548
rect 24578 21496 24584 21548
rect 24636 21536 24642 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 24636 21508 24685 21536
rect 24636 21496 24642 21508
rect 24673 21505 24685 21508
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 24854 21496 24860 21548
rect 24912 21496 24918 21548
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 26053 21499 26111 21505
rect 21591 21440 21956 21468
rect 22204 21440 22600 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 19794 21360 19800 21412
rect 19852 21360 19858 21412
rect 19886 21360 19892 21412
rect 19944 21400 19950 21412
rect 21082 21400 21088 21412
rect 19944 21372 21088 21400
rect 19944 21360 19950 21372
rect 21082 21360 21088 21372
rect 21140 21360 21146 21412
rect 22204 21344 22232 21440
rect 26068 21412 26096 21499
rect 26142 21496 26148 21548
rect 26200 21496 26206 21548
rect 30466 21496 30472 21548
rect 30524 21496 30530 21548
rect 26326 21428 26332 21480
rect 26384 21468 26390 21480
rect 26513 21471 26571 21477
rect 26513 21468 26525 21471
rect 26384 21440 26525 21468
rect 26384 21428 26390 21440
rect 26513 21437 26525 21440
rect 26559 21437 26571 21471
rect 26513 21431 26571 21437
rect 26602 21428 26608 21480
rect 26660 21468 26666 21480
rect 29641 21471 29699 21477
rect 29641 21468 29653 21471
rect 26660 21440 29653 21468
rect 26660 21428 26666 21440
rect 29641 21437 29653 21440
rect 29687 21437 29699 21471
rect 29641 21431 29699 21437
rect 22278 21360 22284 21412
rect 22336 21400 22342 21412
rect 22465 21403 22523 21409
rect 22465 21400 22477 21403
rect 22336 21372 22477 21400
rect 22336 21360 22342 21372
rect 22465 21369 22477 21372
rect 22511 21369 22523 21403
rect 22465 21363 22523 21369
rect 26050 21360 26056 21412
rect 26108 21360 26114 21412
rect 20070 21332 20076 21344
rect 19306 21304 20076 21332
rect 20070 21292 20076 21304
rect 20128 21292 20134 21344
rect 22186 21292 22192 21344
rect 22244 21292 22250 21344
rect 24394 21292 24400 21344
rect 24452 21332 24458 21344
rect 26234 21332 26240 21344
rect 24452 21304 26240 21332
rect 24452 21292 24458 21304
rect 26234 21292 26240 21304
rect 26292 21292 26298 21344
rect 1104 21242 30820 21264
rect 1104 21190 4664 21242
rect 4716 21190 4728 21242
rect 4780 21190 4792 21242
rect 4844 21190 4856 21242
rect 4908 21190 4920 21242
rect 4972 21190 12092 21242
rect 12144 21190 12156 21242
rect 12208 21190 12220 21242
rect 12272 21190 12284 21242
rect 12336 21190 12348 21242
rect 12400 21190 19520 21242
rect 19572 21190 19584 21242
rect 19636 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 26948 21242
rect 27000 21190 27012 21242
rect 27064 21190 27076 21242
rect 27128 21190 27140 21242
rect 27192 21190 27204 21242
rect 27256 21190 30820 21242
rect 1104 21168 30820 21190
rect 5166 21088 5172 21140
rect 5224 21128 5230 21140
rect 5353 21131 5411 21137
rect 5353 21128 5365 21131
rect 5224 21100 5365 21128
rect 5224 21088 5230 21100
rect 5353 21097 5365 21100
rect 5399 21097 5411 21131
rect 5353 21091 5411 21097
rect 5368 20992 5396 21091
rect 6086 21088 6092 21140
rect 6144 21088 6150 21140
rect 6638 21088 6644 21140
rect 6696 21088 6702 21140
rect 8938 21088 8944 21140
rect 8996 21088 9002 21140
rect 12345 21131 12403 21137
rect 12345 21097 12357 21131
rect 12391 21128 12403 21131
rect 12434 21128 12440 21140
rect 12391 21100 12440 21128
rect 12391 21097 12403 21100
rect 12345 21091 12403 21097
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 13538 21088 13544 21140
rect 13596 21128 13602 21140
rect 13596 21100 18276 21128
rect 13596 21088 13602 21100
rect 5445 20995 5503 21001
rect 5445 20992 5457 20995
rect 5368 20964 5457 20992
rect 5445 20961 5457 20964
rect 5491 20961 5503 20995
rect 5445 20955 5503 20961
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20893 1731 20927
rect 1673 20887 1731 20893
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 1688 20788 1716 20887
rect 3326 20884 3332 20936
rect 3384 20924 3390 20936
rect 3786 20924 3792 20936
rect 3384 20896 3792 20924
rect 3384 20884 3390 20896
rect 3786 20884 3792 20896
rect 3844 20924 3850 20936
rect 3973 20927 4031 20933
rect 3973 20924 3985 20927
rect 3844 20896 3985 20924
rect 3844 20884 3850 20896
rect 3973 20893 3985 20896
rect 4019 20893 4031 20927
rect 6104 20924 6132 21088
rect 6181 20927 6239 20933
rect 6181 20924 6193 20927
rect 6104 20896 6193 20924
rect 3973 20887 4031 20893
rect 6181 20893 6193 20896
rect 6227 20893 6239 20927
rect 6181 20887 6239 20893
rect 4240 20859 4298 20865
rect 4240 20825 4252 20859
rect 4286 20856 4298 20859
rect 6273 20859 6331 20865
rect 6273 20856 6285 20859
rect 4286 20828 6285 20856
rect 4286 20825 4298 20828
rect 4240 20819 4298 20825
rect 6273 20825 6285 20828
rect 6319 20825 6331 20859
rect 6656 20856 6684 21088
rect 8956 21001 8984 21088
rect 9309 21063 9367 21069
rect 9309 21029 9321 21063
rect 9355 21060 9367 21063
rect 9398 21060 9404 21072
rect 9355 21032 9404 21060
rect 9355 21029 9367 21032
rect 9309 21023 9367 21029
rect 9398 21020 9404 21032
rect 9456 21020 9462 21072
rect 14274 21020 14280 21072
rect 14332 21060 14338 21072
rect 15746 21060 15752 21072
rect 14332 21032 15752 21060
rect 14332 21020 14338 21032
rect 15746 21020 15752 21032
rect 15804 21020 15810 21072
rect 18248 21060 18276 21100
rect 20346 21088 20352 21140
rect 20404 21088 20410 21140
rect 20898 21088 20904 21140
rect 20956 21088 20962 21140
rect 22186 21128 22192 21140
rect 21928 21100 22192 21128
rect 20916 21060 20944 21088
rect 18248 21032 20944 21060
rect 8941 20995 8999 21001
rect 8941 20961 8953 20995
rect 8987 20961 8999 20995
rect 8941 20955 8999 20961
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 11388 20964 18460 20992
rect 11388 20952 11394 20964
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9766 20924 9772 20936
rect 9723 20896 9772 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9766 20884 9772 20896
rect 9824 20884 9830 20936
rect 12268 20933 12296 20964
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20924 12311 20927
rect 14921 20927 14979 20933
rect 12299 20896 12333 20924
rect 12299 20893 12311 20896
rect 12253 20887 12311 20893
rect 14921 20893 14933 20927
rect 14967 20924 14979 20927
rect 15194 20924 15200 20936
rect 14967 20896 15200 20924
rect 14967 20893 14979 20896
rect 14921 20887 14979 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15470 20884 15476 20936
rect 15528 20884 15534 20936
rect 16945 20927 17003 20933
rect 16945 20893 16957 20927
rect 16991 20893 17003 20927
rect 18432 20924 18460 20964
rect 18690 20952 18696 21004
rect 18748 20992 18754 21004
rect 21928 21001 21956 21100
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 22646 21088 22652 21140
rect 22704 21088 22710 21140
rect 23842 21088 23848 21140
rect 23900 21128 23906 21140
rect 26145 21131 26203 21137
rect 26145 21128 26157 21131
rect 23900 21100 26157 21128
rect 23900 21088 23906 21100
rect 26145 21097 26157 21100
rect 26191 21097 26203 21131
rect 26145 21091 26203 21097
rect 22664 21060 22692 21088
rect 24854 21060 24860 21072
rect 22296 21032 22692 21060
rect 22756 21032 24860 21060
rect 22296 21001 22324 21032
rect 22756 21004 22784 21032
rect 19797 20995 19855 21001
rect 19797 20992 19809 20995
rect 18748 20964 19809 20992
rect 18748 20952 18754 20964
rect 19797 20961 19809 20964
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 21913 20995 21971 21001
rect 21913 20992 21925 20995
rect 21775 20964 21925 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 21913 20961 21925 20964
rect 21959 20961 21971 20995
rect 21913 20955 21971 20961
rect 22281 20995 22339 21001
rect 22281 20961 22293 20995
rect 22327 20961 22339 20995
rect 22281 20955 22339 20961
rect 22370 20952 22376 21004
rect 22428 20952 22434 21004
rect 22738 20952 22744 21004
rect 22796 20952 22802 21004
rect 23952 20964 24624 20992
rect 23952 20936 23980 20964
rect 18969 20927 19027 20933
rect 18969 20924 18981 20927
rect 18432 20896 18981 20924
rect 16945 20887 17003 20893
rect 18969 20893 18981 20896
rect 19015 20924 19027 20927
rect 19426 20924 19432 20936
rect 19015 20896 19432 20924
rect 19015 20893 19027 20896
rect 18969 20887 19027 20893
rect 10226 20856 10232 20868
rect 6656 20828 10232 20856
rect 6273 20819 6331 20825
rect 10226 20816 10232 20828
rect 10284 20816 10290 20868
rect 16960 20856 16988 20887
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19886 20884 19892 20936
rect 19944 20884 19950 20936
rect 19978 20884 19984 20936
rect 20036 20884 20042 20936
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 21821 20927 21879 20933
rect 21821 20893 21833 20927
rect 21867 20924 21879 20927
rect 22094 20924 22100 20936
rect 21867 20896 22100 20924
rect 21867 20893 21879 20896
rect 21821 20887 21879 20893
rect 16960 20828 17080 20856
rect 17052 20800 17080 20828
rect 17218 20816 17224 20868
rect 17276 20816 17282 20868
rect 18877 20859 18935 20865
rect 18877 20856 18889 20859
rect 18446 20828 18889 20856
rect 18877 20825 18889 20828
rect 18923 20825 18935 20859
rect 19904 20856 19932 20884
rect 20165 20859 20223 20865
rect 20165 20856 20177 20859
rect 19904 20828 20177 20856
rect 18877 20819 18935 20825
rect 20165 20825 20177 20828
rect 20211 20825 20223 20859
rect 21652 20856 21680 20887
rect 22094 20884 22100 20896
rect 22152 20924 22158 20936
rect 22152 20896 22968 20924
rect 22152 20884 22158 20896
rect 22940 20868 22968 20896
rect 23934 20884 23940 20936
rect 23992 20884 23998 20936
rect 24394 20884 24400 20936
rect 24452 20884 24458 20936
rect 24596 20924 24624 20964
rect 24744 20933 24772 21032
rect 24854 21020 24860 21032
rect 24912 21020 24918 21072
rect 24949 21063 25007 21069
rect 24949 21029 24961 21063
rect 24995 21060 25007 21063
rect 24995 21032 30236 21060
rect 24995 21029 25007 21032
rect 24949 21023 25007 21029
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24872 20964 25053 20992
rect 24744 20927 24823 20933
rect 24596 20896 24716 20924
rect 24744 20896 24777 20927
rect 24688 20868 24716 20896
rect 24765 20893 24777 20896
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 24872 20868 24900 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 26050 20992 26056 21004
rect 25041 20955 25099 20961
rect 25180 20964 26056 20992
rect 22186 20856 22192 20868
rect 21652 20828 22192 20856
rect 20165 20819 20223 20825
rect 22186 20816 22192 20828
rect 22244 20856 22250 20868
rect 22830 20856 22836 20868
rect 22244 20828 22836 20856
rect 22244 20816 22250 20828
rect 22830 20816 22836 20828
rect 22888 20816 22894 20868
rect 22922 20816 22928 20868
rect 22980 20856 22986 20868
rect 23017 20859 23075 20865
rect 23017 20856 23029 20859
rect 22980 20828 23029 20856
rect 22980 20816 22986 20828
rect 23017 20825 23029 20828
rect 23063 20825 23075 20859
rect 23017 20819 23075 20825
rect 23106 20816 23112 20868
rect 23164 20856 23170 20868
rect 24578 20856 24584 20868
rect 23164 20828 24584 20856
rect 23164 20816 23170 20828
rect 24578 20816 24584 20828
rect 24636 20816 24642 20868
rect 24670 20816 24676 20868
rect 24728 20816 24734 20868
rect 24854 20816 24860 20868
rect 24912 20816 24918 20868
rect 8478 20788 8484 20800
rect 1688 20760 8484 20788
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 8754 20748 8760 20800
rect 8812 20788 8818 20800
rect 9401 20791 9459 20797
rect 9401 20788 9413 20791
rect 8812 20760 9413 20788
rect 8812 20748 8818 20760
rect 9401 20757 9413 20760
rect 9447 20757 9459 20791
rect 9401 20751 9459 20757
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 9674 20788 9680 20800
rect 9631 20760 9680 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 14734 20748 14740 20800
rect 14792 20748 14798 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 15657 20791 15715 20797
rect 15657 20788 15669 20791
rect 15528 20760 15669 20788
rect 15528 20748 15534 20760
rect 15657 20757 15669 20760
rect 15703 20757 15715 20791
rect 15657 20751 15715 20757
rect 17034 20748 17040 20800
rect 17092 20748 17098 20800
rect 19242 20748 19248 20800
rect 19300 20748 19306 20800
rect 22557 20791 22615 20797
rect 22557 20757 22569 20791
rect 22603 20788 22615 20791
rect 25180 20788 25208 20964
rect 26050 20952 26056 20964
rect 26108 20992 26114 21004
rect 26329 20995 26387 21001
rect 26329 20992 26341 20995
rect 26108 20964 26341 20992
rect 26108 20952 26114 20964
rect 26329 20961 26341 20964
rect 26375 20961 26387 20995
rect 26789 20995 26847 21001
rect 26789 20992 26801 20995
rect 26329 20955 26387 20961
rect 26436 20964 26801 20992
rect 26436 20933 26464 20964
rect 26789 20961 26801 20964
rect 26835 20961 26847 20995
rect 26789 20955 26847 20961
rect 30208 20933 30236 21032
rect 26421 20927 26479 20933
rect 26421 20893 26433 20927
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20893 26755 20927
rect 26697 20887 26755 20893
rect 26881 20927 26939 20933
rect 26881 20893 26893 20927
rect 26927 20893 26939 20927
rect 26881 20887 26939 20893
rect 30193 20927 30251 20933
rect 30193 20893 30205 20927
rect 30239 20893 30251 20927
rect 30193 20887 30251 20893
rect 26326 20816 26332 20868
rect 26384 20856 26390 20868
rect 26712 20856 26740 20887
rect 26384 20828 26740 20856
rect 26384 20816 26390 20828
rect 22603 20760 25208 20788
rect 22603 20757 22615 20760
rect 22557 20751 22615 20757
rect 25682 20748 25688 20800
rect 25740 20748 25746 20800
rect 26142 20748 26148 20800
rect 26200 20788 26206 20800
rect 26896 20788 26924 20887
rect 26200 20760 26924 20788
rect 26200 20748 26206 20760
rect 30282 20748 30288 20800
rect 30340 20788 30346 20800
rect 30377 20791 30435 20797
rect 30377 20788 30389 20791
rect 30340 20760 30389 20788
rect 30340 20748 30346 20760
rect 30377 20757 30389 20760
rect 30423 20757 30435 20791
rect 30377 20751 30435 20757
rect 1104 20698 30820 20720
rect 1104 20646 5324 20698
rect 5376 20646 5388 20698
rect 5440 20646 5452 20698
rect 5504 20646 5516 20698
rect 5568 20646 5580 20698
rect 5632 20646 12752 20698
rect 12804 20646 12816 20698
rect 12868 20646 12880 20698
rect 12932 20646 12944 20698
rect 12996 20646 13008 20698
rect 13060 20646 20180 20698
rect 20232 20646 20244 20698
rect 20296 20646 20308 20698
rect 20360 20646 20372 20698
rect 20424 20646 20436 20698
rect 20488 20646 27608 20698
rect 27660 20646 27672 20698
rect 27724 20646 27736 20698
rect 27788 20646 27800 20698
rect 27852 20646 27864 20698
rect 27916 20646 30820 20698
rect 1104 20624 30820 20646
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7650 20584 7656 20596
rect 6972 20556 7656 20584
rect 6972 20544 6978 20556
rect 7650 20544 7656 20556
rect 7708 20584 7714 20596
rect 8113 20587 8171 20593
rect 8113 20584 8125 20587
rect 7708 20556 8125 20584
rect 7708 20544 7714 20556
rect 8113 20553 8125 20556
rect 8159 20553 8171 20587
rect 8113 20547 8171 20553
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 9306 20584 9312 20596
rect 8536 20556 9312 20584
rect 8536 20544 8542 20556
rect 9306 20544 9312 20556
rect 9364 20584 9370 20596
rect 10045 20587 10103 20593
rect 10045 20584 10057 20587
rect 9364 20556 10057 20584
rect 9364 20544 9370 20556
rect 10045 20553 10057 20556
rect 10091 20584 10103 20587
rect 10318 20584 10324 20596
rect 10091 20556 10324 20584
rect 10091 20553 10103 20556
rect 10045 20547 10103 20553
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17405 20587 17463 20593
rect 17405 20584 17417 20587
rect 17276 20556 17417 20584
rect 17276 20544 17282 20556
rect 17405 20553 17417 20556
rect 17451 20553 17463 20587
rect 17405 20547 17463 20553
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 19242 20584 19248 20596
rect 18279 20556 19248 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19518 20544 19524 20596
rect 19576 20544 19582 20596
rect 19978 20544 19984 20596
rect 20036 20544 20042 20596
rect 20070 20544 20076 20596
rect 20128 20584 20134 20596
rect 20533 20587 20591 20593
rect 20128 20556 20484 20584
rect 20128 20544 20134 20556
rect 7098 20476 7104 20528
rect 7156 20476 7162 20528
rect 14734 20476 14740 20528
rect 14792 20476 14798 20528
rect 16482 20476 16488 20528
rect 16540 20476 16546 20528
rect 18325 20519 18383 20525
rect 18325 20485 18337 20519
rect 18371 20516 18383 20519
rect 18966 20516 18972 20528
rect 18371 20488 18972 20516
rect 18371 20485 18383 20488
rect 18325 20479 18383 20485
rect 18966 20476 18972 20488
rect 19024 20516 19030 20528
rect 19536 20516 19564 20544
rect 19024 20488 19564 20516
rect 19996 20516 20024 20544
rect 20257 20519 20315 20525
rect 20257 20516 20269 20519
rect 19996 20488 20269 20516
rect 19024 20476 19030 20488
rect 20257 20485 20269 20488
rect 20303 20485 20315 20519
rect 20456 20516 20484 20556
rect 20533 20553 20545 20587
rect 20579 20584 20591 20587
rect 20806 20584 20812 20596
rect 20579 20556 20812 20584
rect 20579 20553 20591 20556
rect 20533 20547 20591 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 23106 20584 23112 20596
rect 22572 20556 23112 20584
rect 22572 20525 22600 20556
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 25225 20587 25283 20593
rect 25225 20553 25237 20587
rect 25271 20584 25283 20587
rect 25682 20584 25688 20596
rect 25271 20556 25688 20584
rect 25271 20553 25283 20556
rect 25225 20547 25283 20553
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 26053 20587 26111 20593
rect 26053 20553 26065 20587
rect 26099 20584 26111 20587
rect 26142 20584 26148 20596
rect 26099 20556 26148 20584
rect 26099 20553 26111 20556
rect 26053 20547 26111 20553
rect 26142 20544 26148 20556
rect 26200 20544 26206 20596
rect 26326 20544 26332 20596
rect 26384 20544 26390 20596
rect 22557 20519 22615 20525
rect 22557 20516 22569 20519
rect 20456 20488 22569 20516
rect 20257 20479 20315 20485
rect 22557 20485 22569 20488
rect 22603 20485 22615 20519
rect 22557 20479 22615 20485
rect 22649 20519 22707 20525
rect 22649 20485 22661 20519
rect 22695 20516 22707 20519
rect 22922 20516 22928 20528
rect 22695 20488 22928 20516
rect 22695 20485 22707 20488
rect 22649 20479 22707 20485
rect 22922 20476 22928 20488
rect 22980 20476 22986 20528
rect 24026 20476 24032 20528
rect 24084 20476 24090 20528
rect 24670 20476 24676 20528
rect 24728 20476 24734 20528
rect 25314 20476 25320 20528
rect 25372 20516 25378 20528
rect 25590 20516 25596 20528
rect 25372 20488 25596 20516
rect 25372 20476 25378 20488
rect 25590 20476 25596 20488
rect 25648 20476 25654 20528
rect 25869 20519 25927 20525
rect 25869 20485 25881 20519
rect 25915 20516 25927 20519
rect 26602 20516 26608 20528
rect 25915 20488 26608 20516
rect 25915 20485 25927 20488
rect 25869 20479 25927 20485
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5868 20420 6377 20448
rect 5868 20408 5874 20420
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 8294 20408 8300 20460
rect 8352 20408 8358 20460
rect 9674 20408 9680 20460
rect 9732 20408 9738 20460
rect 11330 20448 11336 20460
rect 9784 20420 11336 20448
rect 6638 20340 6644 20392
rect 6696 20340 6702 20392
rect 8570 20340 8576 20392
rect 8628 20340 8634 20392
rect 9784 20256 9812 20420
rect 11330 20408 11336 20420
rect 11388 20408 11394 20460
rect 12618 20408 12624 20460
rect 12676 20448 12682 20460
rect 12805 20451 12863 20457
rect 12805 20448 12817 20451
rect 12676 20420 12817 20448
rect 12676 20408 12682 20420
rect 12805 20417 12817 20420
rect 12851 20448 12863 20451
rect 13538 20448 13544 20460
rect 12851 20420 13544 20448
rect 12851 20417 12863 20420
rect 12805 20411 12863 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 19426 20457 19432 20460
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20448 17647 20451
rect 19421 20448 19432 20457
rect 17635 20420 17908 20448
rect 19387 20420 19432 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 10042 20340 10048 20392
rect 10100 20380 10106 20392
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 10100 20352 10609 20380
rect 10100 20340 10106 20352
rect 10597 20349 10609 20352
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12713 20383 12771 20389
rect 12713 20380 12725 20383
rect 12584 20352 12725 20380
rect 12584 20340 12590 20352
rect 12713 20349 12725 20352
rect 12759 20349 12771 20383
rect 12713 20343 12771 20349
rect 14274 20340 14280 20392
rect 14332 20380 14338 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 14332 20352 14473 20380
rect 14332 20340 14338 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 10318 20272 10324 20324
rect 10376 20272 10382 20324
rect 17880 20321 17908 20420
rect 19421 20411 19432 20420
rect 19426 20408 19432 20411
rect 19484 20408 19490 20460
rect 19978 20408 19984 20460
rect 20036 20408 20042 20460
rect 20070 20408 20076 20460
rect 20128 20448 20134 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 20128 20420 20177 20448
rect 20128 20408 20134 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18417 20383 18475 20389
rect 18417 20380 18429 20383
rect 18012 20352 18429 20380
rect 18012 20340 18018 20352
rect 18417 20349 18429 20352
rect 18463 20349 18475 20383
rect 18417 20343 18475 20349
rect 20364 20380 20392 20411
rect 22370 20408 22376 20460
rect 22428 20408 22434 20460
rect 22738 20408 22744 20460
rect 22796 20408 22802 20460
rect 24688 20448 24716 20476
rect 26344 20457 26372 20488
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 25685 20451 25743 20457
rect 25685 20448 25697 20451
rect 24688 20420 25697 20448
rect 25685 20417 25697 20420
rect 25731 20448 25743 20451
rect 26145 20451 26203 20457
rect 26145 20448 26157 20451
rect 25731 20420 26157 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 26145 20417 26157 20420
rect 26191 20417 26203 20451
rect 26145 20411 26203 20417
rect 26329 20451 26387 20457
rect 26329 20417 26341 20451
rect 26375 20417 26387 20451
rect 26329 20411 26387 20417
rect 22756 20380 22784 20408
rect 20364 20352 22784 20380
rect 17865 20315 17923 20321
rect 17865 20281 17877 20315
rect 17911 20281 17923 20315
rect 17865 20275 17923 20281
rect 19150 20272 19156 20324
rect 19208 20312 19214 20324
rect 20364 20312 20392 20352
rect 23014 20340 23020 20392
rect 23072 20340 23078 20392
rect 23290 20340 23296 20392
rect 23348 20340 23354 20392
rect 24486 20340 24492 20392
rect 24544 20380 24550 20392
rect 24765 20383 24823 20389
rect 24765 20380 24777 20383
rect 24544 20352 24777 20380
rect 24544 20340 24550 20352
rect 24765 20349 24777 20352
rect 24811 20380 24823 20383
rect 24854 20380 24860 20392
rect 24811 20352 24860 20380
rect 24811 20349 24823 20352
rect 24765 20343 24823 20349
rect 24854 20340 24860 20352
rect 24912 20340 24918 20392
rect 25409 20383 25467 20389
rect 25409 20349 25421 20383
rect 25455 20349 25467 20383
rect 25409 20343 25467 20349
rect 19208 20284 20392 20312
rect 19208 20272 19214 20284
rect 24946 20272 24952 20324
rect 25004 20312 25010 20324
rect 25424 20312 25452 20343
rect 25004 20284 25452 20312
rect 25004 20272 25010 20284
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 9766 20244 9772 20256
rect 7432 20216 9772 20244
rect 7432 20204 7438 20216
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 10134 20204 10140 20256
rect 10192 20204 10198 20256
rect 11238 20204 11244 20256
rect 11296 20204 11302 20256
rect 13173 20247 13231 20253
rect 13173 20213 13185 20247
rect 13219 20244 13231 20247
rect 13262 20244 13268 20256
rect 13219 20216 13268 20244
rect 13219 20213 13231 20216
rect 13173 20207 13231 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 19521 20247 19579 20253
rect 19521 20213 19533 20247
rect 19567 20244 19579 20247
rect 19978 20244 19984 20256
rect 19567 20216 19984 20244
rect 19567 20213 19579 20216
rect 19521 20207 19579 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20990 20244 20996 20256
rect 20128 20216 20996 20244
rect 20128 20204 20134 20216
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 22925 20247 22983 20253
rect 22925 20213 22937 20247
rect 22971 20244 22983 20247
rect 24670 20244 24676 20256
rect 22971 20216 24676 20244
rect 22971 20213 22983 20216
rect 22925 20207 22983 20213
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 24854 20204 24860 20256
rect 24912 20204 24918 20256
rect 1104 20154 30820 20176
rect 1104 20102 4664 20154
rect 4716 20102 4728 20154
rect 4780 20102 4792 20154
rect 4844 20102 4856 20154
rect 4908 20102 4920 20154
rect 4972 20102 12092 20154
rect 12144 20102 12156 20154
rect 12208 20102 12220 20154
rect 12272 20102 12284 20154
rect 12336 20102 12348 20154
rect 12400 20102 19520 20154
rect 19572 20102 19584 20154
rect 19636 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 26948 20154
rect 27000 20102 27012 20154
rect 27064 20102 27076 20154
rect 27128 20102 27140 20154
rect 27192 20102 27204 20154
rect 27256 20102 30820 20154
rect 1104 20080 30820 20102
rect 6733 20043 6791 20049
rect 6733 20009 6745 20043
rect 6779 20040 6791 20043
rect 7098 20040 7104 20052
rect 6779 20012 7104 20040
rect 6779 20009 6791 20012
rect 6733 20003 6791 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8570 20000 8576 20052
rect 8628 20000 8634 20052
rect 10042 20040 10048 20052
rect 8864 20012 10048 20040
rect 8864 19972 8892 20012
rect 10042 20000 10048 20012
rect 10100 20000 10106 20052
rect 10226 20000 10232 20052
rect 10284 20040 10290 20052
rect 10962 20040 10968 20052
rect 10284 20012 10968 20040
rect 10284 20000 10290 20012
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 11572 20012 12020 20040
rect 11572 20000 11578 20012
rect 2746 19944 8892 19972
rect 8941 19975 8999 19981
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 992 19740 1501 19768
rect 992 19728 998 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 1489 19731 1547 19737
rect 1673 19771 1731 19777
rect 1673 19737 1685 19771
rect 1719 19768 1731 19771
rect 2746 19768 2774 19944
rect 8941 19941 8953 19975
rect 8987 19941 8999 19975
rect 8941 19935 8999 19941
rect 7650 19864 7656 19916
rect 7708 19904 7714 19916
rect 7745 19907 7803 19913
rect 7745 19904 7757 19907
rect 7708 19876 7757 19904
rect 7708 19864 7714 19876
rect 7745 19873 7757 19876
rect 7791 19873 7803 19907
rect 7745 19867 7803 19873
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 1719 19740 2774 19768
rect 5184 19808 6653 19836
rect 1719 19737 1731 19740
rect 1673 19731 1731 19737
rect 5184 19712 5212 19808
rect 6641 19805 6653 19808
rect 6687 19836 6699 19839
rect 7374 19836 7380 19848
rect 6687 19808 7380 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 7760 19768 7788 19867
rect 7926 19864 7932 19916
rect 7984 19864 7990 19916
rect 8110 19796 8116 19848
rect 8168 19796 8174 19848
rect 8205 19839 8263 19845
rect 8205 19805 8217 19839
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 8956 19836 8984 19935
rect 9490 19864 9496 19916
rect 9548 19904 9554 19916
rect 11992 19913 12020 20012
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 15838 20000 15844 20052
rect 15896 20000 15902 20052
rect 20806 20040 20812 20052
rect 18064 20012 20812 20040
rect 12066 19932 12072 19984
rect 12124 19932 12130 19984
rect 15470 19972 15476 19984
rect 14568 19944 15476 19972
rect 11977 19907 12035 19913
rect 9548 19876 10456 19904
rect 9548 19864 9554 19876
rect 8803 19808 8984 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 7834 19768 7840 19780
rect 7760 19740 7840 19768
rect 7834 19728 7840 19740
rect 7892 19768 7898 19780
rect 8220 19768 8248 19799
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 9858 19836 9864 19848
rect 9364 19808 9864 19836
rect 9364 19796 9370 19808
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 7892 19740 8248 19768
rect 7892 19728 7898 19740
rect 5166 19660 5172 19712
rect 5224 19660 5230 19712
rect 7190 19660 7196 19712
rect 7248 19660 7254 19712
rect 7929 19703 7987 19709
rect 7929 19669 7941 19703
rect 7975 19700 7987 19703
rect 8754 19700 8760 19712
rect 7975 19672 8760 19700
rect 7975 19669 7987 19672
rect 7929 19663 7987 19669
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 9398 19660 9404 19712
rect 9456 19660 9462 19712
rect 10428 19700 10456 19876
rect 11977 19873 11989 19907
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 13078 19864 13084 19916
rect 13136 19864 13142 19916
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14568 19913 14596 19944
rect 15470 19932 15476 19944
rect 15528 19972 15534 19984
rect 17954 19972 17960 19984
rect 15528 19944 17960 19972
rect 15528 19932 15534 19944
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 14553 19907 14611 19913
rect 14553 19904 14565 19907
rect 14516 19876 14565 19904
rect 14516 19864 14522 19876
rect 14553 19873 14565 19876
rect 14599 19873 14611 19907
rect 14553 19867 14611 19873
rect 14737 19907 14795 19913
rect 14737 19873 14749 19907
rect 14783 19904 14795 19907
rect 15102 19904 15108 19916
rect 14783 19876 15108 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15102 19864 15108 19876
rect 15160 19864 15166 19916
rect 17494 19864 17500 19916
rect 17552 19864 17558 19916
rect 12345 19839 12403 19845
rect 11992 19808 12296 19836
rect 11238 19728 11244 19780
rect 11296 19728 11302 19780
rect 11698 19728 11704 19780
rect 11756 19728 11762 19780
rect 11992 19768 12020 19808
rect 11900 19740 12020 19768
rect 11900 19700 11928 19740
rect 12066 19728 12072 19780
rect 12124 19728 12130 19780
rect 12268 19768 12296 19808
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 12434 19836 12440 19848
rect 12391 19808 12440 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 12526 19796 12532 19848
rect 12584 19796 12590 19848
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 12897 19799 12955 19805
rect 12544 19768 12572 19796
rect 12912 19768 12940 19799
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15562 19836 15568 19848
rect 14884 19808 15568 19836
rect 14884 19796 14890 19808
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15746 19796 15752 19848
rect 15804 19836 15810 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15804 19808 15945 19836
rect 15804 19796 15810 19808
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 15979 19808 17417 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 17405 19805 17417 19808
rect 17451 19836 17463 19839
rect 18064 19836 18092 20012
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 20990 20000 20996 20052
rect 21048 20000 21054 20052
rect 22370 20000 22376 20052
rect 22428 20040 22434 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 22428 20012 22845 20040
rect 22428 20000 22434 20012
rect 22833 20009 22845 20012
rect 22879 20009 22891 20043
rect 22833 20003 22891 20009
rect 22848 19972 22876 20003
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 23348 20012 23673 20040
rect 23348 20000 23354 20012
rect 23661 20009 23673 20012
rect 23707 20009 23719 20043
rect 23661 20003 23719 20009
rect 24026 20000 24032 20052
rect 24084 20040 24090 20052
rect 24121 20043 24179 20049
rect 24121 20040 24133 20043
rect 24084 20012 24133 20040
rect 24084 20000 24090 20012
rect 24121 20009 24133 20012
rect 24167 20009 24179 20043
rect 24121 20003 24179 20009
rect 24762 20000 24768 20052
rect 24820 20000 24826 20052
rect 24854 20000 24860 20052
rect 24912 20000 24918 20052
rect 24780 19972 24808 20000
rect 22848 19944 23520 19972
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 17451 19808 18092 19836
rect 18156 19876 19257 19904
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 16022 19768 16028 19780
rect 12268 19740 12434 19768
rect 12544 19740 12940 19768
rect 13648 19740 16028 19768
rect 12406 19712 12434 19740
rect 10428 19672 11928 19700
rect 11974 19660 11980 19712
rect 12032 19700 12038 19712
rect 12253 19703 12311 19709
rect 12253 19700 12265 19703
rect 12032 19672 12265 19700
rect 12032 19660 12038 19672
rect 12253 19669 12265 19672
rect 12299 19669 12311 19703
rect 12253 19663 12311 19669
rect 12342 19660 12348 19712
rect 12400 19700 12434 19712
rect 13648 19700 13676 19740
rect 16022 19728 16028 19740
rect 16080 19728 16086 19780
rect 17034 19728 17040 19780
rect 17092 19768 17098 19780
rect 18156 19768 18184 19876
rect 19245 19873 19257 19876
rect 19291 19904 19303 19907
rect 21085 19907 21143 19913
rect 19291 19876 20760 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 18874 19796 18880 19848
rect 18932 19796 18938 19848
rect 20732 19836 20760 19876
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 22094 19904 22100 19916
rect 21131 19876 22100 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 20898 19836 20904 19848
rect 20732 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19836 20962 19848
rect 21100 19836 21128 19867
rect 22094 19864 22100 19876
rect 22152 19904 22158 19916
rect 23492 19913 23520 19944
rect 23584 19944 24808 19972
rect 23477 19907 23535 19913
rect 22152 19876 22600 19904
rect 22152 19864 22158 19876
rect 20956 19808 21128 19836
rect 22572 19836 22600 19876
rect 23477 19873 23489 19907
rect 23523 19873 23535 19907
rect 23477 19867 23535 19873
rect 23014 19836 23020 19848
rect 22572 19808 23020 19836
rect 20956 19796 20962 19808
rect 23014 19796 23020 19808
rect 23072 19836 23078 19848
rect 23584 19836 23612 19944
rect 24872 19904 24900 20000
rect 30374 19932 30380 19984
rect 30432 19932 30438 19984
rect 23860 19876 24900 19904
rect 23860 19845 23888 19876
rect 23072 19808 23612 19836
rect 23845 19839 23903 19845
rect 23072 19796 23078 19808
rect 23845 19805 23857 19839
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 24029 19839 24087 19845
rect 24029 19805 24041 19839
rect 24075 19805 24087 19839
rect 24029 19799 24087 19805
rect 19521 19771 19579 19777
rect 19521 19768 19533 19771
rect 17092 19740 18184 19768
rect 19352 19740 19533 19768
rect 17092 19728 17098 19740
rect 12400 19672 13676 19700
rect 12400 19660 12406 19672
rect 13722 19660 13728 19712
rect 13780 19660 13786 19712
rect 19061 19703 19119 19709
rect 19061 19669 19073 19703
rect 19107 19700 19119 19703
rect 19352 19700 19380 19740
rect 19521 19737 19533 19740
rect 19567 19737 19579 19771
rect 19521 19731 19579 19737
rect 19978 19728 19984 19780
rect 20036 19728 20042 19780
rect 20806 19728 20812 19780
rect 20864 19728 20870 19780
rect 21358 19728 21364 19780
rect 21416 19728 21422 19780
rect 21818 19728 21824 19780
rect 21876 19728 21882 19780
rect 24044 19768 24072 19799
rect 24670 19796 24676 19848
rect 24728 19836 24734 19848
rect 30193 19839 30251 19845
rect 30193 19836 30205 19839
rect 24728 19808 30205 19836
rect 24728 19796 24734 19808
rect 30193 19805 30205 19808
rect 30239 19805 30251 19839
rect 30193 19799 30251 19805
rect 25038 19768 25044 19780
rect 22848 19740 25044 19768
rect 19107 19672 19380 19700
rect 20824 19700 20852 19728
rect 22848 19700 22876 19740
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 20824 19672 22876 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 22922 19660 22928 19712
rect 22980 19660 22986 19712
rect 1104 19610 30820 19632
rect 1104 19558 5324 19610
rect 5376 19558 5388 19610
rect 5440 19558 5452 19610
rect 5504 19558 5516 19610
rect 5568 19558 5580 19610
rect 5632 19558 12752 19610
rect 12804 19558 12816 19610
rect 12868 19558 12880 19610
rect 12932 19558 12944 19610
rect 12996 19558 13008 19610
rect 13060 19558 20180 19610
rect 20232 19558 20244 19610
rect 20296 19558 20308 19610
rect 20360 19558 20372 19610
rect 20424 19558 20436 19610
rect 20488 19558 27608 19610
rect 27660 19558 27672 19610
rect 27724 19558 27736 19610
rect 27788 19558 27800 19610
rect 27852 19558 27864 19610
rect 27916 19558 30820 19610
rect 1104 19536 30820 19558
rect 1581 19499 1639 19505
rect 1581 19465 1593 19499
rect 1627 19496 1639 19499
rect 4338 19496 4344 19508
rect 1627 19468 4344 19496
rect 1627 19465 1639 19468
rect 1581 19459 1639 19465
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 5077 19499 5135 19505
rect 5077 19496 5089 19499
rect 4488 19468 5089 19496
rect 4488 19456 4494 19468
rect 5077 19465 5089 19468
rect 5123 19465 5135 19499
rect 7006 19496 7012 19508
rect 5077 19459 5135 19465
rect 6932 19468 7012 19496
rect 5261 19431 5319 19437
rect 5261 19428 5273 19431
rect 4830 19400 5273 19428
rect 5261 19397 5273 19400
rect 5307 19397 5319 19431
rect 5261 19391 5319 19397
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 3326 19320 3332 19372
rect 3384 19320 3390 19372
rect 4614 19320 4620 19372
rect 4672 19320 4678 19372
rect 5166 19360 5172 19372
rect 4816 19332 5172 19360
rect 3602 19252 3608 19304
rect 3660 19252 3666 19304
rect 4632 19292 4660 19320
rect 4816 19292 4844 19332
rect 5166 19320 5172 19332
rect 5224 19360 5230 19372
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 5224 19332 5365 19360
rect 5224 19320 5230 19332
rect 5353 19329 5365 19332
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 4632 19264 4844 19292
rect 6362 19252 6368 19304
rect 6420 19292 6426 19304
rect 6932 19301 6960 19468
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7374 19456 7380 19508
rect 7432 19456 7438 19508
rect 7469 19499 7527 19505
rect 7469 19465 7481 19499
rect 7515 19496 7527 19499
rect 7926 19496 7932 19508
rect 7515 19468 7932 19496
rect 7515 19465 7527 19468
rect 7469 19459 7527 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8110 19456 8116 19508
rect 8168 19456 8174 19508
rect 8294 19456 8300 19508
rect 8352 19456 8358 19508
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12437 19499 12495 19505
rect 12437 19496 12449 19499
rect 12124 19468 12449 19496
rect 12124 19456 12130 19468
rect 12437 19465 12449 19468
rect 12483 19465 12495 19499
rect 15562 19496 15568 19508
rect 12437 19459 12495 19465
rect 14200 19468 15568 19496
rect 7834 19428 7840 19440
rect 7024 19400 7840 19428
rect 7024 19369 7052 19400
rect 7834 19388 7840 19400
rect 7892 19388 7898 19440
rect 8128 19428 8156 19456
rect 7944 19400 8156 19428
rect 8312 19428 8340 19456
rect 8941 19431 8999 19437
rect 8941 19428 8953 19431
rect 8312 19400 8953 19428
rect 7009 19363 7067 19369
rect 7009 19329 7021 19363
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 7944 19369 7972 19400
rect 8941 19397 8953 19400
rect 8987 19397 8999 19431
rect 14200 19428 14228 19468
rect 15562 19456 15568 19468
rect 15620 19496 15626 19508
rect 15620 19468 19656 19496
rect 15620 19456 15626 19468
rect 16209 19431 16267 19437
rect 8941 19391 8999 19397
rect 10704 19400 14228 19428
rect 14292 19400 16160 19428
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 6917 19295 6975 19301
rect 6917 19292 6929 19295
rect 6420 19264 6929 19292
rect 6420 19252 6426 19264
rect 6917 19261 6929 19264
rect 6963 19292 6975 19295
rect 8036 19292 8064 19323
rect 10594 19320 10600 19372
rect 10652 19360 10658 19372
rect 10704 19369 10732 19400
rect 14292 19372 14320 19400
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10652 19332 10701 19360
rect 10652 19320 10658 19332
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10689 19323 10747 19329
rect 10962 19320 10968 19372
rect 11020 19360 11026 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11020 19332 11529 19360
rect 11020 19320 11026 19332
rect 11517 19329 11529 19332
rect 11563 19360 11575 19363
rect 11606 19360 11612 19372
rect 11563 19332 11612 19360
rect 11563 19329 11575 19332
rect 11517 19323 11575 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 12342 19320 12348 19372
rect 12400 19320 12406 19372
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12618 19360 12624 19372
rect 12575 19332 12624 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 13170 19320 13176 19372
rect 13228 19360 13234 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 13228 19332 13277 19360
rect 13228 19320 13234 19332
rect 13265 19329 13277 19332
rect 13311 19329 13323 19363
rect 13265 19323 13323 19329
rect 13354 19320 13360 19372
rect 13412 19320 13418 19372
rect 13633 19363 13691 19369
rect 13633 19329 13645 19363
rect 13679 19360 13691 19363
rect 13679 19332 13952 19360
rect 13679 19329 13691 19332
rect 13633 19323 13691 19329
rect 6963 19264 8064 19292
rect 12452 19292 12480 19320
rect 13081 19295 13139 19301
rect 13081 19292 13093 19295
rect 12452 19264 13093 19292
rect 6963 19261 6975 19264
rect 6917 19255 6975 19261
rect 13081 19261 13093 19264
rect 13127 19261 13139 19295
rect 13081 19255 13139 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13722 19292 13728 19304
rect 13587 19264 13728 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 12434 19224 12440 19236
rect 6604 19196 12440 19224
rect 6604 19184 6610 19196
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 13924 19224 13952 19332
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 14185 19363 14243 19369
rect 14185 19360 14197 19363
rect 14056 19332 14197 19360
rect 14056 19320 14062 19332
rect 14185 19329 14197 19332
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 14200 19292 14228 19323
rect 14274 19320 14280 19372
rect 14332 19320 14338 19372
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19360 14703 19363
rect 14826 19360 14832 19372
rect 14691 19332 14832 19360
rect 14691 19329 14703 19332
rect 14645 19323 14703 19329
rect 14826 19320 14832 19332
rect 14884 19360 14890 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14884 19332 14933 19360
rect 14884 19320 14890 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15286 19320 15292 19372
rect 15344 19360 15350 19372
rect 15473 19363 15531 19369
rect 15473 19360 15485 19363
rect 15344 19332 15485 19360
rect 15344 19320 15350 19332
rect 15473 19329 15485 19332
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15565 19363 15623 19369
rect 15565 19329 15577 19363
rect 15611 19329 15623 19363
rect 15565 19323 15623 19329
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14200 19264 14688 19292
rect 14660 19236 14688 19264
rect 14936 19264 15117 19292
rect 14936 19236 14964 19264
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 13924 19196 14412 19224
rect 5442 19116 5448 19168
rect 5500 19156 5506 19168
rect 9490 19156 9496 19168
rect 5500 19128 9496 19156
rect 5500 19116 5506 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10778 19156 10784 19168
rect 9732 19128 10784 19156
rect 9732 19116 9738 19128
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 11940 19128 12173 19156
rect 11940 19116 11946 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12161 19119 12219 19125
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 14277 19159 14335 19165
rect 14277 19156 14289 19159
rect 14240 19128 14289 19156
rect 14240 19116 14246 19128
rect 14277 19125 14289 19128
rect 14323 19125 14335 19159
rect 14384 19156 14412 19196
rect 14642 19184 14648 19236
rect 14700 19184 14706 19236
rect 14918 19184 14924 19236
rect 14976 19184 14982 19236
rect 14829 19159 14887 19165
rect 14829 19156 14841 19159
rect 14384 19128 14841 19156
rect 14277 19119 14335 19125
rect 14829 19125 14841 19128
rect 14875 19156 14887 19159
rect 15194 19156 15200 19168
rect 14875 19128 15200 19156
rect 14875 19125 14887 19128
rect 14829 19119 14887 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15304 19156 15332 19320
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15580 19292 15608 19323
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 16132 19360 16160 19400
rect 16209 19397 16221 19431
rect 16255 19428 16267 19431
rect 16482 19428 16488 19440
rect 16255 19400 16488 19428
rect 16255 19397 16267 19400
rect 16209 19391 16267 19397
rect 16482 19388 16488 19400
rect 16540 19388 16546 19440
rect 17034 19428 17040 19440
rect 16684 19400 17040 19428
rect 16684 19369 16712 19400
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 17494 19388 17500 19440
rect 17552 19388 17558 19440
rect 18874 19388 18880 19440
rect 18932 19428 18938 19440
rect 19426 19428 19432 19440
rect 18932 19400 19432 19428
rect 18932 19388 18938 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 19518 19388 19524 19440
rect 19576 19388 19582 19440
rect 19628 19437 19656 19468
rect 20898 19456 20904 19508
rect 20956 19456 20962 19508
rect 21545 19499 21603 19505
rect 21545 19465 21557 19499
rect 21591 19496 21603 19499
rect 21818 19496 21824 19508
rect 21591 19468 21824 19496
rect 21591 19465 21603 19468
rect 21545 19459 21603 19465
rect 21818 19456 21824 19468
rect 21876 19456 21882 19508
rect 22281 19499 22339 19505
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 22922 19496 22928 19508
rect 22327 19468 22928 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 22922 19456 22928 19468
rect 22980 19456 22986 19508
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 23440 19468 26188 19496
rect 23440 19456 23446 19468
rect 19613 19431 19671 19437
rect 19613 19397 19625 19431
rect 19659 19397 19671 19431
rect 19613 19391 19671 19397
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 22244 19400 22385 19428
rect 22244 19388 22250 19400
rect 22373 19397 22385 19400
rect 22419 19428 22431 19431
rect 23400 19428 23428 19456
rect 24762 19428 24768 19440
rect 22419 19400 23428 19428
rect 24596 19400 24768 19428
rect 22419 19397 22431 19400
rect 22373 19391 22431 19397
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16132 19332 16681 19360
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 19536 19360 19564 19388
rect 24596 19369 24624 19400
rect 24762 19388 24768 19400
rect 24820 19388 24826 19440
rect 25866 19388 25872 19440
rect 25924 19388 25930 19440
rect 26160 19428 26188 19468
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 26292 19468 26341 19496
rect 26292 19456 26298 19468
rect 26329 19465 26341 19468
rect 26375 19465 26387 19499
rect 26329 19459 26387 19465
rect 29825 19431 29883 19437
rect 29825 19428 29837 19431
rect 26160 19400 29837 19428
rect 29825 19397 29837 19400
rect 29871 19397 29883 19431
rect 29825 19391 29883 19397
rect 21453 19363 21511 19369
rect 21453 19360 21465 19363
rect 19536 19332 21465 19360
rect 16669 19323 16727 19329
rect 21453 19329 21465 19332
rect 21499 19329 21511 19363
rect 21453 19323 21511 19329
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 30282 19320 30288 19372
rect 30340 19360 30346 19372
rect 30377 19363 30435 19369
rect 30377 19360 30389 19363
rect 30340 19332 30389 19360
rect 30340 19320 30346 19332
rect 30377 19329 30389 19332
rect 30423 19329 30435 19363
rect 30377 19323 30435 19329
rect 15436 19264 15884 19292
rect 15436 19252 15442 19264
rect 15856 19236 15884 19264
rect 16942 19252 16948 19304
rect 17000 19252 17006 19304
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 20956 19264 22569 19292
rect 20956 19252 20962 19264
rect 22557 19261 22569 19264
rect 22603 19292 22615 19295
rect 22603 19264 22692 19292
rect 22603 19261 22615 19264
rect 22557 19255 22615 19261
rect 15838 19184 15844 19236
rect 15896 19184 15902 19236
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 15304 19128 16221 19156
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16390 19116 16396 19168
rect 16448 19116 16454 19168
rect 18414 19116 18420 19168
rect 18472 19116 18478 19168
rect 21910 19116 21916 19168
rect 21968 19116 21974 19168
rect 22664 19156 22692 19264
rect 24854 19252 24860 19304
rect 24912 19252 24918 19304
rect 24946 19156 24952 19168
rect 22664 19128 24952 19156
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 1104 19066 30820 19088
rect 1104 19014 4664 19066
rect 4716 19014 4728 19066
rect 4780 19014 4792 19066
rect 4844 19014 4856 19066
rect 4908 19014 4920 19066
rect 4972 19014 12092 19066
rect 12144 19014 12156 19066
rect 12208 19014 12220 19066
rect 12272 19014 12284 19066
rect 12336 19014 12348 19066
rect 12400 19014 19520 19066
rect 19572 19014 19584 19066
rect 19636 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 26948 19066
rect 27000 19014 27012 19066
rect 27064 19014 27076 19066
rect 27128 19014 27140 19066
rect 27192 19014 27204 19066
rect 27256 19014 30820 19066
rect 1104 18992 30820 19014
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3660 18924 3801 18952
rect 3660 18912 3666 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 6546 18952 6552 18964
rect 3789 18915 3847 18921
rect 4172 18924 6552 18952
rect 1581 18887 1639 18893
rect 1581 18853 1593 18887
rect 1627 18884 1639 18887
rect 4172 18884 4200 18924
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 6696 18924 6745 18952
rect 6696 18912 6702 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 11146 18952 11152 18964
rect 6733 18915 6791 18921
rect 10152 18924 11152 18952
rect 1627 18856 4200 18884
rect 4249 18887 4307 18893
rect 1627 18853 1639 18856
rect 1581 18847 1639 18853
rect 4249 18853 4261 18887
rect 4295 18853 4307 18887
rect 4249 18847 4307 18853
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 3973 18751 4031 18757
rect 3973 18717 3985 18751
rect 4019 18748 4031 18751
rect 4264 18748 4292 18847
rect 4338 18844 4344 18896
rect 4396 18884 4402 18896
rect 5074 18884 5080 18896
rect 4396 18856 5080 18884
rect 4396 18844 4402 18856
rect 5074 18844 5080 18856
rect 5132 18884 5138 18896
rect 5629 18887 5687 18893
rect 5629 18884 5641 18887
rect 5132 18856 5641 18884
rect 5132 18844 5138 18856
rect 5629 18853 5641 18856
rect 5675 18853 5687 18887
rect 5629 18847 5687 18853
rect 5813 18887 5871 18893
rect 5813 18853 5825 18887
rect 5859 18884 5871 18887
rect 9950 18884 9956 18896
rect 5859 18856 6684 18884
rect 5859 18853 5871 18856
rect 5813 18847 5871 18853
rect 4801 18819 4859 18825
rect 4801 18816 4813 18819
rect 4019 18720 4292 18748
rect 4356 18788 4813 18816
rect 4019 18717 4031 18720
rect 3973 18711 4031 18717
rect 4356 18624 4384 18788
rect 4801 18785 4813 18788
rect 4847 18816 4859 18819
rect 5442 18816 5448 18828
rect 4847 18788 5448 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 6273 18819 6331 18825
rect 6273 18816 6285 18819
rect 6104 18788 6285 18816
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 4488 18720 4629 18748
rect 4488 18708 4494 18720
rect 4617 18717 4629 18720
rect 4663 18748 4675 18751
rect 5166 18748 5172 18760
rect 4663 18720 5172 18748
rect 4663 18717 4675 18720
rect 4617 18711 4675 18717
rect 5166 18708 5172 18720
rect 5224 18748 5230 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5224 18720 5365 18748
rect 5224 18708 5230 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 6104 18624 6132 18788
rect 6273 18785 6285 18788
rect 6319 18785 6331 18819
rect 6273 18779 6331 18785
rect 6181 18751 6239 18757
rect 6181 18717 6193 18751
rect 6227 18717 6239 18751
rect 6181 18711 6239 18717
rect 6196 18680 6224 18711
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 6546 18708 6552 18760
rect 6604 18708 6610 18760
rect 6656 18748 6684 18856
rect 6748 18856 9956 18884
rect 6748 18828 6776 18856
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 10042 18844 10048 18896
rect 10100 18884 10106 18896
rect 10152 18893 10180 18924
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 11333 18955 11391 18961
rect 11333 18921 11345 18955
rect 11379 18952 11391 18955
rect 11698 18952 11704 18964
rect 11379 18924 11704 18952
rect 11379 18921 11391 18924
rect 11333 18915 11391 18921
rect 11698 18912 11704 18924
rect 11756 18912 11762 18964
rect 11790 18912 11796 18964
rect 11848 18912 11854 18964
rect 13170 18912 13176 18964
rect 13228 18912 13234 18964
rect 13265 18955 13323 18961
rect 13265 18921 13277 18955
rect 13311 18952 13323 18955
rect 13354 18952 13360 18964
rect 13311 18924 13360 18952
rect 13311 18921 13323 18924
rect 13265 18915 13323 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14608 18924 14657 18952
rect 14608 18912 14614 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 16942 18912 16948 18964
rect 17000 18912 17006 18964
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 21358 18912 21364 18964
rect 21416 18952 21422 18964
rect 21545 18955 21603 18961
rect 21545 18952 21557 18955
rect 21416 18924 21557 18952
rect 21416 18912 21422 18924
rect 21545 18921 21557 18924
rect 21591 18921 21603 18955
rect 21545 18915 21603 18921
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 25317 18955 25375 18961
rect 25317 18952 25329 18955
rect 24912 18924 25329 18952
rect 24912 18912 24918 18924
rect 25317 18921 25329 18924
rect 25363 18921 25375 18955
rect 25317 18915 25375 18921
rect 10137 18887 10195 18893
rect 10137 18884 10149 18887
rect 10100 18856 10149 18884
rect 10100 18844 10106 18856
rect 10137 18853 10149 18856
rect 10183 18853 10195 18887
rect 10137 18847 10195 18853
rect 10505 18887 10563 18893
rect 10505 18853 10517 18887
rect 10551 18884 10563 18887
rect 11808 18884 11836 18912
rect 14366 18884 14372 18896
rect 10551 18856 12940 18884
rect 10551 18853 10563 18856
rect 10505 18847 10563 18853
rect 6730 18776 6736 18828
rect 6788 18776 6794 18828
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 9723 18788 10732 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6656 18720 6837 18748
rect 6825 18717 6837 18720
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 6914 18708 6920 18760
rect 6972 18708 6978 18760
rect 7006 18708 7012 18760
rect 7064 18708 7070 18760
rect 7190 18708 7196 18760
rect 7248 18708 7254 18760
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18748 9827 18751
rect 10134 18748 10140 18760
rect 9815 18720 10140 18748
rect 9815 18717 9827 18720
rect 9769 18711 9827 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10704 18757 10732 18788
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 10836 18788 11805 18816
rect 10836 18776 10842 18788
rect 10689 18751 10747 18757
rect 10689 18717 10701 18751
rect 10735 18748 10747 18751
rect 10962 18748 10968 18760
rect 10735 18720 10968 18748
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 11057 18751 11115 18757
rect 11057 18717 11069 18751
rect 11103 18717 11115 18751
rect 11057 18711 11115 18717
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18748 11207 18751
rect 11195 18720 11376 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 7208 18680 7236 18708
rect 6196 18652 7236 18680
rect 9674 18640 9680 18692
rect 9732 18640 9738 18692
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 10781 18683 10839 18689
rect 10781 18680 10793 18683
rect 10560 18652 10793 18680
rect 10560 18640 10566 18652
rect 10781 18649 10793 18652
rect 10827 18649 10839 18683
rect 10781 18643 10839 18649
rect 10870 18640 10876 18692
rect 10928 18640 10934 18692
rect 4338 18572 4344 18624
rect 4396 18572 4402 18624
rect 4709 18615 4767 18621
rect 4709 18581 4721 18615
rect 4755 18612 4767 18615
rect 4982 18612 4988 18624
rect 4755 18584 4988 18612
rect 4755 18581 4767 18584
rect 4709 18575 4767 18581
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 9692 18612 9720 18640
rect 6144 18584 9720 18612
rect 10321 18615 10379 18621
rect 6144 18572 6150 18584
rect 10321 18581 10333 18615
rect 10367 18612 10379 18615
rect 10410 18612 10416 18624
rect 10367 18584 10416 18612
rect 10367 18581 10379 18584
rect 10321 18575 10379 18581
rect 10410 18572 10416 18584
rect 10468 18612 10474 18624
rect 11072 18612 11100 18711
rect 11348 18624 11376 18720
rect 10468 18584 11100 18612
rect 10468 18572 10474 18584
rect 11330 18572 11336 18624
rect 11388 18572 11394 18624
rect 11440 18612 11468 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 12912 18816 12940 18856
rect 13740 18856 14372 18884
rect 13740 18825 13768 18856
rect 14366 18844 14372 18856
rect 14424 18884 14430 18896
rect 14461 18887 14519 18893
rect 14461 18884 14473 18887
rect 14424 18856 14473 18884
rect 14424 18844 14430 18856
rect 14461 18853 14473 18856
rect 14507 18853 14519 18887
rect 14461 18847 14519 18853
rect 17405 18887 17463 18893
rect 17405 18853 17417 18887
rect 17451 18853 17463 18887
rect 17405 18847 17463 18853
rect 17972 18856 19932 18884
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12912 18788 13553 18816
rect 11517 18751 11575 18757
rect 11517 18717 11529 18751
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11532 18680 11560 18711
rect 11606 18708 11612 18760
rect 11664 18708 11670 18760
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 12912 18757 12940 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 13725 18819 13783 18825
rect 13725 18785 13737 18819
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 15654 18816 15660 18828
rect 14240 18788 15660 18816
rect 14240 18776 14246 18788
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18717 12955 18751
rect 12897 18711 12955 18717
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18748 13231 18751
rect 13262 18748 13268 18760
rect 13219 18720 13268 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13262 18708 13268 18720
rect 13320 18748 13326 18760
rect 13449 18751 13507 18757
rect 13449 18748 13461 18751
rect 13320 18720 13461 18748
rect 13320 18708 13326 18720
rect 13449 18717 13461 18720
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 12526 18680 12532 18692
rect 11532 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 12676 18652 13001 18680
rect 12676 18640 12682 18652
rect 12989 18649 13001 18652
rect 13035 18680 13047 18683
rect 13648 18680 13676 18711
rect 14642 18708 14648 18760
rect 14700 18708 14706 18760
rect 14826 18708 14832 18760
rect 14884 18748 14890 18760
rect 15013 18751 15071 18757
rect 15013 18748 15025 18751
rect 14884 18720 15025 18748
rect 14884 18708 14890 18720
rect 15013 18717 15025 18720
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 13035 18652 13676 18680
rect 15672 18680 15700 18776
rect 16301 18751 16359 18757
rect 16301 18717 16313 18751
rect 16347 18748 16359 18751
rect 16390 18748 16396 18760
rect 16347 18720 16396 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17420 18748 17448 18847
rect 17972 18828 18000 18856
rect 17954 18776 17960 18828
rect 18012 18776 18018 18828
rect 19904 18816 19932 18856
rect 20070 18844 20076 18896
rect 20128 18884 20134 18896
rect 20128 18856 21128 18884
rect 20128 18844 20134 18856
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 19904 18788 19993 18816
rect 19981 18785 19993 18788
rect 20027 18816 20039 18819
rect 20898 18816 20904 18828
rect 20027 18788 20904 18816
rect 20027 18785 20039 18788
rect 19981 18779 20039 18785
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 20990 18776 20996 18828
rect 21048 18776 21054 18828
rect 21100 18816 21128 18856
rect 21450 18844 21456 18896
rect 21508 18844 21514 18896
rect 25222 18844 25228 18896
rect 25280 18844 25286 18896
rect 21100 18788 21496 18816
rect 17175 18720 17448 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 19242 18708 19248 18760
rect 19300 18748 19306 18760
rect 19300 18720 20576 18748
rect 19300 18708 19306 18720
rect 17773 18683 17831 18689
rect 17773 18680 17785 18683
rect 15672 18652 17785 18680
rect 13035 18649 13047 18652
rect 12989 18643 13047 18649
rect 17773 18649 17785 18652
rect 17819 18680 17831 18683
rect 18414 18680 18420 18692
rect 17819 18652 18420 18680
rect 17819 18649 17831 18652
rect 17773 18643 17831 18649
rect 18414 18640 18420 18652
rect 18472 18640 18478 18692
rect 19797 18683 19855 18689
rect 19797 18649 19809 18683
rect 19843 18680 19855 18683
rect 20441 18683 20499 18689
rect 20441 18680 20453 18683
rect 19843 18652 20453 18680
rect 19843 18649 19855 18652
rect 19797 18643 19855 18649
rect 20441 18649 20453 18652
rect 20487 18649 20499 18683
rect 20548 18680 20576 18720
rect 21082 18708 21088 18760
rect 21140 18748 21146 18760
rect 21468 18757 21496 18788
rect 22094 18776 22100 18828
rect 22152 18776 22158 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23492 18788 24041 18816
rect 21177 18751 21235 18757
rect 21177 18748 21189 18751
rect 21140 18720 21189 18748
rect 21140 18708 21146 18720
rect 21177 18717 21189 18720
rect 21223 18717 21235 18751
rect 21177 18711 21235 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 21729 18751 21787 18757
rect 21729 18717 21741 18751
rect 21775 18748 21787 18751
rect 21910 18748 21916 18760
rect 21775 18720 21916 18748
rect 21775 18717 21787 18720
rect 21729 18711 21787 18717
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 23492 18734 23520 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24029 18779 24087 18785
rect 24394 18776 24400 18828
rect 24452 18816 24458 18828
rect 24673 18819 24731 18825
rect 24452 18788 24624 18816
rect 24452 18776 24458 18788
rect 24121 18751 24179 18757
rect 24121 18748 24133 18751
rect 23768 18720 24133 18748
rect 20548 18652 21404 18680
rect 20441 18643 20499 18649
rect 15470 18612 15476 18624
rect 11440 18584 15476 18612
rect 15470 18572 15476 18584
rect 15528 18572 15534 18624
rect 16117 18615 16175 18621
rect 16117 18581 16129 18615
rect 16163 18612 16175 18615
rect 16482 18612 16488 18624
rect 16163 18584 16488 18612
rect 16163 18581 16175 18584
rect 16117 18575 16175 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 17865 18615 17923 18621
rect 17865 18581 17877 18615
rect 17911 18612 17923 18615
rect 18322 18612 18328 18624
rect 17911 18584 18328 18612
rect 17911 18581 17923 18584
rect 17865 18575 17923 18581
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 19886 18572 19892 18624
rect 19944 18572 19950 18624
rect 21266 18572 21272 18624
rect 21324 18572 21330 18624
rect 21376 18612 21404 18652
rect 22370 18640 22376 18692
rect 22428 18640 22434 18692
rect 23768 18612 23796 18720
rect 24121 18717 24133 18720
rect 24167 18748 24179 18751
rect 24596 18748 24624 18788
rect 24673 18785 24685 18819
rect 24719 18816 24731 18819
rect 24946 18816 24952 18828
rect 24719 18788 24952 18816
rect 24719 18785 24731 18788
rect 24673 18779 24731 18785
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25056 18788 25636 18816
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24167 18720 24532 18748
rect 24596 18720 24777 18748
rect 24167 18717 24179 18720
rect 24121 18711 24179 18717
rect 24504 18692 24532 18720
rect 24765 18717 24777 18720
rect 24811 18748 24823 18751
rect 25056 18748 25084 18788
rect 24811 18720 25084 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 25501 18751 25559 18757
rect 25501 18748 25513 18751
rect 25280 18720 25513 18748
rect 25280 18708 25286 18720
rect 25501 18717 25513 18720
rect 25547 18717 25559 18751
rect 25608 18748 25636 18788
rect 26234 18776 26240 18828
rect 26292 18776 26298 18828
rect 26602 18748 26608 18760
rect 25608 18720 26608 18748
rect 25501 18711 25559 18717
rect 26602 18708 26608 18720
rect 26660 18748 26666 18760
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26660 18720 26893 18748
rect 26660 18708 26666 18720
rect 26881 18717 26893 18720
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 24486 18640 24492 18692
rect 24544 18640 24550 18692
rect 24857 18683 24915 18689
rect 24596 18652 24808 18680
rect 21376 18584 23796 18612
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24596 18612 24624 18652
rect 23900 18584 24624 18612
rect 24780 18612 24808 18652
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 25593 18683 25651 18689
rect 25593 18680 25605 18683
rect 24903 18652 25605 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 25593 18649 25605 18652
rect 25639 18649 25651 18683
rect 30208 18680 30236 18711
rect 25593 18643 25651 18649
rect 25700 18652 30236 18680
rect 25700 18612 25728 18652
rect 24780 18584 25728 18612
rect 23900 18572 23906 18584
rect 26418 18572 26424 18624
rect 26476 18572 26482 18624
rect 30374 18572 30380 18624
rect 30432 18572 30438 18624
rect 1104 18522 30820 18544
rect 1104 18470 5324 18522
rect 5376 18470 5388 18522
rect 5440 18470 5452 18522
rect 5504 18470 5516 18522
rect 5568 18470 5580 18522
rect 5632 18470 12752 18522
rect 12804 18470 12816 18522
rect 12868 18470 12880 18522
rect 12932 18470 12944 18522
rect 12996 18470 13008 18522
rect 13060 18470 20180 18522
rect 20232 18470 20244 18522
rect 20296 18470 20308 18522
rect 20360 18470 20372 18522
rect 20424 18470 20436 18522
rect 20488 18470 27608 18522
rect 27660 18470 27672 18522
rect 27724 18470 27736 18522
rect 27788 18470 27800 18522
rect 27852 18470 27864 18522
rect 27916 18470 30820 18522
rect 1104 18448 30820 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 1627 18380 6500 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 5074 18300 5080 18352
rect 5132 18340 5138 18352
rect 5353 18343 5411 18349
rect 5353 18340 5365 18343
rect 5132 18312 5365 18340
rect 5132 18300 5138 18312
rect 5353 18309 5365 18312
rect 5399 18340 5411 18343
rect 5902 18340 5908 18352
rect 5399 18312 5908 18340
rect 5399 18309 5411 18312
rect 5353 18303 5411 18309
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 6472 18340 6500 18380
rect 6546 18368 6552 18420
rect 6604 18408 6610 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 6604 18380 7757 18408
rect 6604 18368 6610 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 7913 18411 7971 18417
rect 7913 18377 7925 18411
rect 7959 18408 7971 18411
rect 8573 18411 8631 18417
rect 8573 18408 8585 18411
rect 7959 18380 8585 18408
rect 7959 18377 7971 18380
rect 7913 18371 7971 18377
rect 8573 18377 8585 18380
rect 8619 18377 8631 18411
rect 8573 18371 8631 18377
rect 9309 18411 9367 18417
rect 9309 18377 9321 18411
rect 9355 18408 9367 18411
rect 9398 18408 9404 18420
rect 9355 18380 9404 18408
rect 9355 18377 9367 18380
rect 9309 18371 9367 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 11606 18408 11612 18420
rect 11563 18380 11612 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 12250 18408 12256 18420
rect 11756 18380 12256 18408
rect 11756 18368 11762 18380
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12618 18408 12624 18420
rect 12360 18380 12624 18408
rect 6730 18340 6736 18352
rect 6472 18312 6736 18340
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 7650 18340 7656 18352
rect 7024 18312 7656 18340
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 7024 18216 7052 18312
rect 7392 18281 7420 18312
rect 7650 18300 7656 18312
rect 7708 18340 7714 18352
rect 8018 18340 8024 18352
rect 7708 18312 8024 18340
rect 7708 18300 7714 18312
rect 8018 18300 8024 18312
rect 8076 18300 8082 18352
rect 8113 18343 8171 18349
rect 8113 18309 8125 18343
rect 8159 18340 8171 18343
rect 8662 18340 8668 18352
rect 8159 18312 8668 18340
rect 8159 18309 8171 18312
rect 8113 18303 8171 18309
rect 8662 18300 8668 18312
rect 8720 18340 8726 18352
rect 11882 18340 11888 18352
rect 8720 18312 11888 18340
rect 8720 18300 8726 18312
rect 11882 18300 11888 18312
rect 11940 18300 11946 18352
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7524 18244 8217 18272
rect 7524 18232 7530 18244
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8205 18235 8263 18241
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 10183 18275 10241 18281
rect 8536 18244 9720 18272
rect 8536 18232 8542 18244
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 7006 18204 7012 18216
rect 5859 18176 7012 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7392 18176 7665 18204
rect 7392 18148 7420 18176
rect 7653 18173 7665 18176
rect 7699 18204 7711 18207
rect 7742 18204 7748 18216
rect 7699 18176 7748 18204
rect 7699 18173 7711 18176
rect 7653 18167 7711 18173
rect 7742 18164 7748 18176
rect 7800 18204 7806 18216
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 7800 18176 8309 18204
rect 7800 18164 7806 18176
rect 8297 18173 8309 18176
rect 8343 18173 8355 18207
rect 8297 18167 8355 18173
rect 9490 18164 9496 18216
rect 9548 18164 9554 18216
rect 9692 18213 9720 18244
rect 10183 18241 10195 18275
rect 10229 18272 10241 18275
rect 10229 18244 10364 18272
rect 10229 18241 10241 18244
rect 10183 18235 10241 18241
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18173 9735 18207
rect 9677 18167 9735 18173
rect 9769 18207 9827 18213
rect 9769 18173 9781 18207
rect 9815 18173 9827 18207
rect 9769 18167 9827 18173
rect 5166 18096 5172 18148
rect 5224 18136 5230 18148
rect 5629 18139 5687 18145
rect 5629 18136 5641 18139
rect 5224 18108 5641 18136
rect 5224 18096 5230 18108
rect 5629 18105 5641 18108
rect 5675 18105 5687 18139
rect 5629 18099 5687 18105
rect 7374 18096 7380 18148
rect 7432 18096 7438 18148
rect 7561 18139 7619 18145
rect 7561 18105 7573 18139
rect 7607 18136 7619 18139
rect 9600 18136 9628 18167
rect 9784 18136 9812 18167
rect 9858 18164 9864 18216
rect 9916 18204 9922 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 9916 18176 10057 18204
rect 9916 18164 9922 18176
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10336 18204 10364 18244
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 10597 18275 10655 18281
rect 10597 18272 10609 18275
rect 10468 18244 10609 18272
rect 10468 18232 10474 18244
rect 10597 18241 10609 18244
rect 10643 18241 10655 18275
rect 10597 18235 10655 18241
rect 10873 18275 10931 18281
rect 10873 18241 10885 18275
rect 10919 18272 10931 18275
rect 10962 18272 10968 18284
rect 10919 18244 10968 18272
rect 10919 18241 10931 18244
rect 10873 18235 10931 18241
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18241 11207 18275
rect 11149 18235 11207 18241
rect 10502 18204 10508 18216
rect 10336 18176 10508 18204
rect 10045 18167 10103 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 11057 18207 11115 18213
rect 11057 18173 11069 18207
rect 11103 18204 11115 18207
rect 11164 18204 11192 18235
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11606 18272 11612 18284
rect 11388 18244 11612 18272
rect 11388 18232 11394 18244
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 12360 18281 12388 18380
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 13004 18380 13645 18408
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18272 12587 18275
rect 13004 18272 13032 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 13633 18371 13691 18377
rect 14366 18368 14372 18420
rect 14424 18368 14430 18420
rect 20070 18408 20076 18420
rect 17512 18380 20076 18408
rect 12575 18244 13032 18272
rect 13081 18275 13139 18281
rect 12575 18241 12587 18244
rect 12529 18235 12587 18241
rect 13081 18241 13093 18275
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 11103 18176 11192 18204
rect 11241 18207 11299 18213
rect 11103 18173 11115 18176
rect 11057 18167 11115 18173
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11287 18176 11713 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 10134 18136 10140 18148
rect 7607 18108 7972 18136
rect 9600 18108 9720 18136
rect 9784 18108 10140 18136
rect 7607 18105 7619 18108
rect 7561 18099 7619 18105
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7466 18068 7472 18080
rect 7340 18040 7472 18068
rect 7340 18028 7346 18040
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7944 18077 7972 18108
rect 7929 18071 7987 18077
rect 7929 18037 7941 18071
rect 7975 18037 7987 18071
rect 7929 18031 7987 18037
rect 8018 18028 8024 18080
rect 8076 18068 8082 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 8076 18040 8217 18068
rect 8076 18028 8082 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 9692 18068 9720 18108
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 10321 18139 10379 18145
rect 10321 18136 10333 18139
rect 10284 18108 10333 18136
rect 10284 18096 10290 18108
rect 10321 18105 10333 18108
rect 10367 18105 10379 18139
rect 10520 18136 10548 18164
rect 10796 18136 10824 18167
rect 11790 18164 11796 18216
rect 11848 18164 11854 18216
rect 11882 18164 11888 18216
rect 11940 18164 11946 18216
rect 11974 18164 11980 18216
rect 12032 18164 12038 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12176 18176 12449 18204
rect 10520 18108 10824 18136
rect 10321 18099 10379 18105
rect 10045 18071 10103 18077
rect 10045 18068 10057 18071
rect 9692 18040 10057 18068
rect 8205 18031 8263 18037
rect 10045 18037 10057 18040
rect 10091 18037 10103 18071
rect 10045 18031 10103 18037
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 12176 18068 12204 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 12250 18096 12256 18148
rect 12308 18136 12314 18148
rect 13096 18136 13124 18235
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 14384 18281 14412 18368
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 16942 18232 16948 18284
rect 17000 18232 17006 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17402 18272 17408 18284
rect 17359 18244 17408 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 17512 18281 17540 18380
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 20257 18411 20315 18417
rect 20257 18377 20269 18411
rect 20303 18408 20315 18411
rect 20346 18408 20352 18420
rect 20303 18380 20352 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 20346 18368 20352 18380
rect 20404 18408 20410 18420
rect 20993 18411 21051 18417
rect 20993 18408 21005 18411
rect 20404 18380 21005 18408
rect 20404 18368 20410 18380
rect 20993 18377 21005 18380
rect 21039 18408 21051 18411
rect 21266 18408 21272 18420
rect 21039 18380 21272 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 22370 18368 22376 18420
rect 22428 18368 22434 18420
rect 22830 18368 22836 18420
rect 22888 18368 22894 18420
rect 25777 18411 25835 18417
rect 25777 18377 25789 18411
rect 25823 18408 25835 18411
rect 25866 18408 25872 18420
rect 25823 18380 25872 18408
rect 25823 18377 25835 18380
rect 25777 18371 25835 18377
rect 25866 18368 25872 18380
rect 25924 18368 25930 18420
rect 19058 18340 19064 18352
rect 18800 18312 19064 18340
rect 18800 18281 18828 18312
rect 19058 18300 19064 18312
rect 19116 18340 19122 18352
rect 19242 18340 19248 18352
rect 19116 18312 19248 18340
rect 19116 18300 19122 18312
rect 19242 18300 19248 18312
rect 19300 18300 19306 18352
rect 21082 18300 21088 18352
rect 21140 18300 21146 18352
rect 21361 18343 21419 18349
rect 21361 18309 21373 18343
rect 21407 18340 21419 18343
rect 21407 18312 22692 18340
rect 21407 18309 21419 18312
rect 21361 18303 21419 18309
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 15194 18164 15200 18216
rect 15252 18204 15258 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 15252 18176 16681 18204
rect 15252 18164 15258 18176
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 16298 18136 16304 18148
rect 12308 18108 13308 18136
rect 12308 18096 12314 18108
rect 11664 18040 12204 18068
rect 11664 18028 11670 18040
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 12492 18040 12817 18068
rect 12492 18028 12498 18040
rect 12805 18037 12817 18040
rect 12851 18068 12863 18071
rect 13170 18068 13176 18080
rect 12851 18040 13176 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 13280 18077 13308 18108
rect 14476 18108 16304 18136
rect 13265 18071 13323 18077
rect 13265 18037 13277 18071
rect 13311 18037 13323 18071
rect 13265 18031 13323 18037
rect 14182 18028 14188 18080
rect 14240 18068 14246 18080
rect 14476 18077 14504 18108
rect 16298 18096 16304 18108
rect 16356 18136 16362 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 16356 18108 16865 18136
rect 16356 18096 16362 18108
rect 16853 18105 16865 18108
rect 16899 18136 16911 18139
rect 17512 18136 17540 18235
rect 19886 18232 19892 18284
rect 19944 18272 19950 18284
rect 20349 18275 20407 18281
rect 20349 18272 20361 18275
rect 19944 18244 20361 18272
rect 19944 18232 19950 18244
rect 20349 18241 20361 18244
rect 20395 18272 20407 18275
rect 20714 18272 20720 18284
rect 20395 18244 20720 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18272 20959 18275
rect 21100 18272 21128 18300
rect 20947 18244 21128 18272
rect 21177 18275 21235 18281
rect 20947 18241 20959 18244
rect 20901 18235 20959 18241
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18173 20039 18207
rect 19981 18167 20039 18173
rect 20809 18207 20867 18213
rect 20809 18173 20821 18207
rect 20855 18204 20867 18207
rect 21192 18204 21220 18235
rect 21266 18232 21272 18284
rect 21324 18272 21330 18284
rect 22204 18281 22232 18312
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21324 18244 22017 18272
rect 21324 18232 21330 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 22554 18232 22560 18284
rect 22612 18232 22618 18284
rect 22664 18281 22692 18312
rect 24486 18300 24492 18352
rect 24544 18340 24550 18352
rect 25409 18343 25467 18349
rect 25409 18340 25421 18343
rect 24544 18312 25421 18340
rect 24544 18300 24550 18312
rect 25409 18309 25421 18312
rect 25455 18340 25467 18343
rect 25958 18340 25964 18352
rect 25455 18312 25964 18340
rect 25455 18309 25467 18312
rect 25409 18303 25467 18309
rect 25958 18300 25964 18312
rect 26016 18340 26022 18352
rect 27430 18340 27436 18352
rect 26016 18312 27436 18340
rect 26016 18300 26022 18312
rect 27430 18300 27436 18312
rect 27488 18300 27494 18352
rect 22649 18275 22707 18281
rect 22649 18241 22661 18275
rect 22695 18241 22707 18275
rect 22649 18235 22707 18241
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18241 22891 18275
rect 22833 18235 22891 18241
rect 20855 18176 21220 18204
rect 22281 18207 22339 18213
rect 20855 18173 20867 18176
rect 20809 18167 20867 18173
rect 22281 18173 22293 18207
rect 22327 18204 22339 18207
rect 22848 18204 22876 18235
rect 23382 18232 23388 18284
rect 23440 18232 23446 18284
rect 25038 18232 25044 18284
rect 25096 18272 25102 18284
rect 25133 18275 25191 18281
rect 25133 18272 25145 18275
rect 25096 18244 25145 18272
rect 25096 18232 25102 18244
rect 25133 18241 25145 18244
rect 25179 18272 25191 18275
rect 25685 18275 25743 18281
rect 25685 18272 25697 18275
rect 25179 18244 25697 18272
rect 25179 18241 25191 18244
rect 25133 18235 25191 18241
rect 25685 18241 25697 18244
rect 25731 18241 25743 18275
rect 25685 18235 25743 18241
rect 30193 18275 30251 18281
rect 30193 18241 30205 18275
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 22327 18176 22876 18204
rect 22327 18173 22339 18176
rect 22281 18167 22339 18173
rect 16899 18108 17540 18136
rect 19996 18136 20024 18167
rect 20070 18136 20076 18148
rect 19996 18108 20076 18136
rect 16899 18105 16911 18108
rect 16853 18099 16911 18105
rect 20070 18096 20076 18108
rect 20128 18136 20134 18148
rect 20625 18139 20683 18145
rect 20625 18136 20637 18139
rect 20128 18108 20637 18136
rect 20128 18096 20134 18108
rect 20625 18105 20637 18108
rect 20671 18136 20683 18139
rect 22848 18136 22876 18176
rect 23477 18207 23535 18213
rect 23477 18173 23489 18207
rect 23523 18204 23535 18207
rect 23566 18204 23572 18216
rect 23523 18176 23572 18204
rect 23523 18173 23535 18176
rect 23477 18167 23535 18173
rect 23566 18164 23572 18176
rect 23624 18204 23630 18216
rect 23842 18204 23848 18216
rect 23624 18176 23848 18204
rect 23624 18164 23630 18176
rect 23842 18164 23848 18176
rect 23900 18164 23906 18216
rect 23017 18139 23075 18145
rect 23017 18136 23029 18139
rect 20671 18108 22784 18136
rect 22848 18108 23029 18136
rect 20671 18105 20683 18108
rect 20625 18099 20683 18105
rect 14461 18071 14519 18077
rect 14461 18068 14473 18071
rect 14240 18040 14473 18068
rect 14240 18028 14246 18040
rect 14461 18037 14473 18040
rect 14507 18037 14519 18071
rect 14461 18031 14519 18037
rect 16758 18028 16764 18080
rect 16816 18028 16822 18080
rect 17494 18028 17500 18080
rect 17552 18028 17558 18080
rect 18690 18028 18696 18080
rect 18748 18028 18754 18080
rect 21821 18071 21879 18077
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 22646 18068 22652 18080
rect 21867 18040 22652 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 22756 18068 22784 18108
rect 23017 18105 23029 18108
rect 23063 18105 23075 18139
rect 23017 18099 23075 18105
rect 30208 18068 30236 18235
rect 22756 18040 30236 18068
rect 30282 18028 30288 18080
rect 30340 18068 30346 18080
rect 30377 18071 30435 18077
rect 30377 18068 30389 18071
rect 30340 18040 30389 18068
rect 30340 18028 30346 18040
rect 30377 18037 30389 18040
rect 30423 18037 30435 18071
rect 30377 18031 30435 18037
rect 1104 17978 30820 18000
rect 1104 17926 4664 17978
rect 4716 17926 4728 17978
rect 4780 17926 4792 17978
rect 4844 17926 4856 17978
rect 4908 17926 4920 17978
rect 4972 17926 12092 17978
rect 12144 17926 12156 17978
rect 12208 17926 12220 17978
rect 12272 17926 12284 17978
rect 12336 17926 12348 17978
rect 12400 17926 19520 17978
rect 19572 17926 19584 17978
rect 19636 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 26948 17978
rect 27000 17926 27012 17978
rect 27064 17926 27076 17978
rect 27128 17926 27140 17978
rect 27192 17926 27204 17978
rect 27256 17926 30820 17978
rect 1104 17904 30820 17926
rect 4982 17824 4988 17876
rect 5040 17824 5046 17876
rect 5350 17824 5356 17876
rect 5408 17864 5414 17876
rect 6178 17864 6184 17876
rect 5408 17836 6184 17864
rect 5408 17824 5414 17836
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 6273 17867 6331 17873
rect 6273 17833 6285 17867
rect 6319 17864 6331 17867
rect 6454 17864 6460 17876
rect 6319 17836 6460 17864
rect 6319 17833 6331 17836
rect 6273 17827 6331 17833
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 9401 17867 9459 17873
rect 9401 17833 9413 17867
rect 9447 17864 9459 17867
rect 9490 17864 9496 17876
rect 9447 17836 9496 17864
rect 9447 17833 9459 17836
rect 9401 17827 9459 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 10686 17864 10692 17876
rect 9824 17836 10692 17864
rect 9824 17824 9830 17836
rect 10686 17824 10692 17836
rect 10744 17864 10750 17876
rect 10870 17864 10876 17876
rect 10744 17836 10876 17864
rect 10744 17824 10750 17836
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 17000 17836 18889 17864
rect 17000 17824 17006 17836
rect 18877 17833 18889 17836
rect 18923 17864 18935 17867
rect 19334 17864 19340 17876
rect 18923 17836 19340 17864
rect 18923 17833 18935 17836
rect 18877 17827 18935 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 19705 17867 19763 17873
rect 19705 17833 19717 17867
rect 19751 17864 19763 17867
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 19751 17836 20269 17864
rect 19751 17833 19763 17836
rect 19705 17827 19763 17833
rect 20257 17833 20269 17836
rect 20303 17864 20315 17867
rect 21082 17864 21088 17876
rect 20303 17836 21088 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 21450 17824 21456 17876
rect 21508 17824 21514 17876
rect 6638 17796 6644 17808
rect 5828 17768 6644 17796
rect 5718 17728 5724 17740
rect 5276 17700 5724 17728
rect 5166 17620 5172 17672
rect 5224 17620 5230 17672
rect 5276 17669 5304 17700
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17629 5319 17663
rect 5261 17623 5319 17629
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 5629 17663 5687 17669
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 5828 17660 5856 17768
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 6730 17756 6736 17808
rect 6788 17796 6794 17808
rect 6788 17768 10916 17796
rect 6788 17756 6794 17768
rect 10888 17740 10916 17768
rect 11238 17756 11244 17808
rect 11296 17796 11302 17808
rect 14182 17796 14188 17808
rect 11296 17768 14188 17796
rect 11296 17756 11302 17768
rect 14182 17756 14188 17768
rect 14240 17756 14246 17808
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 16724 17768 17264 17796
rect 16724 17756 16730 17768
rect 5994 17688 6000 17740
rect 6052 17728 6058 17740
rect 9122 17728 9128 17740
rect 6052 17700 9128 17728
rect 6052 17688 6058 17700
rect 5675 17632 5856 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5902 17620 5908 17672
rect 5960 17620 5966 17672
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 6656 17669 6684 17700
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 10502 17728 10508 17740
rect 9600 17700 10508 17728
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 6730 17620 6736 17672
rect 6788 17620 6794 17672
rect 6914 17620 6920 17672
rect 6972 17660 6978 17672
rect 7101 17663 7159 17669
rect 7101 17660 7113 17663
rect 6972 17632 7113 17660
rect 6972 17620 6978 17632
rect 7101 17629 7113 17632
rect 7147 17660 7159 17663
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 7147 17632 7665 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 7837 17663 7895 17669
rect 7837 17660 7849 17663
rect 7800 17632 7849 17660
rect 7800 17620 7806 17632
rect 7837 17629 7849 17632
rect 7883 17629 7895 17663
rect 7837 17623 7895 17629
rect 8662 17620 8668 17672
rect 8720 17660 8726 17672
rect 9600 17669 9628 17700
rect 10502 17688 10508 17700
rect 10560 17688 10566 17740
rect 10870 17688 10876 17740
rect 10928 17728 10934 17740
rect 11974 17728 11980 17740
rect 10928 17700 11980 17728
rect 10928 17688 10934 17700
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 14274 17688 14280 17740
rect 14332 17688 14338 17740
rect 17034 17688 17040 17740
rect 17092 17728 17098 17740
rect 17129 17731 17187 17737
rect 17129 17728 17141 17731
rect 17092 17700 17141 17728
rect 17092 17688 17098 17700
rect 17129 17697 17141 17700
rect 17175 17697 17187 17731
rect 17236 17728 17264 17768
rect 18966 17756 18972 17808
rect 19024 17756 19030 17808
rect 21468 17796 21496 17824
rect 20088 17768 21496 17796
rect 17402 17728 17408 17740
rect 17236 17700 17408 17728
rect 17129 17691 17187 17697
rect 17402 17688 17408 17700
rect 17460 17728 17466 17740
rect 18984 17728 19012 17756
rect 17460 17700 19012 17728
rect 17460 17688 17466 17700
rect 9585 17663 9643 17669
rect 9585 17660 9597 17663
rect 8720 17632 9597 17660
rect 8720 17620 8726 17632
rect 9585 17629 9597 17632
rect 9631 17629 9643 17663
rect 9585 17623 9643 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17660 9735 17663
rect 9766 17660 9772 17672
rect 9723 17632 9772 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10410 17660 10416 17672
rect 9999 17632 10416 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 5471 17595 5529 17601
rect 5471 17561 5483 17595
rect 5517 17561 5529 17595
rect 5471 17555 5529 17561
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5486 17524 5514 17555
rect 5040 17496 5514 17524
rect 5920 17524 5948 17620
rect 6089 17595 6147 17601
rect 6089 17561 6101 17595
rect 6135 17592 6147 17595
rect 6270 17592 6276 17604
rect 6135 17564 6276 17592
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 6270 17552 6276 17564
rect 6328 17552 6334 17604
rect 6564 17592 6592 17620
rect 9490 17592 9496 17604
rect 6564 17564 9496 17592
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 9876 17592 9904 17623
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 13722 17620 13728 17672
rect 13780 17620 13786 17672
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 16264 17632 16528 17660
rect 16264 17620 16270 17632
rect 10226 17592 10232 17604
rect 9876 17564 10232 17592
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 14553 17595 14611 17601
rect 14553 17592 14565 17595
rect 13924 17564 14565 17592
rect 6822 17524 6828 17536
rect 5920 17496 6828 17524
rect 5040 17484 5046 17496
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7006 17484 7012 17536
rect 7064 17484 7070 17536
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17524 7895 17527
rect 8294 17524 8300 17536
rect 7883 17496 8300 17524
rect 7883 17493 7895 17496
rect 7837 17487 7895 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 13630 17524 13636 17536
rect 9088 17496 13636 17524
rect 9088 17484 9094 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13924 17533 13952 17564
rect 14553 17561 14565 17564
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 15286 17552 15292 17604
rect 15344 17552 15350 17604
rect 16301 17595 16359 17601
rect 16301 17561 16313 17595
rect 16347 17561 16359 17595
rect 16500 17592 16528 17632
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16666 17620 16672 17672
rect 16724 17620 16730 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17629 16819 17663
rect 16761 17623 16819 17629
rect 16776 17592 16804 17623
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 18690 17660 18696 17672
rect 18538 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 18984 17660 19012 17700
rect 20088 17669 20116 17768
rect 20346 17688 20352 17740
rect 20404 17688 20410 17740
rect 24762 17688 24768 17740
rect 24820 17728 24826 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24820 17700 24869 17728
rect 24820 17688 24826 17700
rect 24857 17697 24869 17700
rect 24903 17697 24915 17731
rect 24857 17691 24915 17697
rect 26605 17731 26663 17737
rect 26605 17697 26617 17731
rect 26651 17728 26663 17731
rect 26651 17700 27384 17728
rect 26651 17697 26663 17700
rect 26605 17691 26663 17697
rect 27356 17672 27384 17700
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18984 17632 19257 17660
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 17392 17595 17450 17601
rect 17392 17592 17404 17595
rect 16500 17564 16804 17592
rect 17052 17564 17404 17592
rect 16301 17555 16359 17561
rect 13909 17527 13967 17533
rect 13909 17493 13921 17527
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15838 17524 15844 17536
rect 14792 17496 15844 17524
rect 14792 17484 14798 17496
rect 15838 17484 15844 17496
rect 15896 17524 15902 17536
rect 16316 17524 16344 17555
rect 17052 17533 17080 17564
rect 17392 17561 17404 17564
rect 17438 17561 17450 17595
rect 19260 17592 19288 17623
rect 27338 17620 27344 17672
rect 27396 17620 27402 17672
rect 27430 17620 27436 17672
rect 27488 17620 27494 17672
rect 20990 17592 20996 17604
rect 19260 17564 20996 17592
rect 17392 17555 17450 17561
rect 20990 17552 20996 17564
rect 21048 17552 21054 17604
rect 25130 17552 25136 17604
rect 25188 17552 25194 17604
rect 27525 17595 27583 17601
rect 27525 17592 27537 17595
rect 26358 17564 27537 17592
rect 27525 17561 27537 17564
rect 27571 17561 27583 17595
rect 27525 17555 27583 17561
rect 15896 17496 16344 17524
rect 17037 17527 17095 17533
rect 15896 17484 15902 17496
rect 17037 17493 17049 17527
rect 17083 17493 17095 17527
rect 17037 17487 17095 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 19794 17524 19800 17536
rect 17644 17496 19800 17524
rect 17644 17484 17650 17496
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 19886 17484 19892 17536
rect 19944 17484 19950 17536
rect 26694 17484 26700 17536
rect 26752 17484 26758 17536
rect 1104 17434 30820 17456
rect 1104 17382 5324 17434
rect 5376 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 12752 17434
rect 12804 17382 12816 17434
rect 12868 17382 12880 17434
rect 12932 17382 12944 17434
rect 12996 17382 13008 17434
rect 13060 17382 20180 17434
rect 20232 17382 20244 17434
rect 20296 17382 20308 17434
rect 20360 17382 20372 17434
rect 20424 17382 20436 17434
rect 20488 17382 27608 17434
rect 27660 17382 27672 17434
rect 27724 17382 27736 17434
rect 27788 17382 27800 17434
rect 27852 17382 27864 17434
rect 27916 17382 30820 17434
rect 1104 17360 30820 17382
rect 4982 17280 4988 17332
rect 5040 17280 5046 17332
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5224 17292 5457 17320
rect 5224 17280 5230 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6454 17320 6460 17332
rect 6227 17292 6460 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6604 17292 6837 17320
rect 6604 17280 6610 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 6825 17283 6883 17289
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 7248 17292 7788 17320
rect 7248 17280 7254 17292
rect 7006 17252 7012 17264
rect 4632 17224 7012 17252
rect 4632 17193 4660 17224
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 7760 17261 7788 17292
rect 8662 17280 8668 17332
rect 8720 17280 8726 17332
rect 8956 17292 9628 17320
rect 7745 17255 7803 17261
rect 7745 17221 7757 17255
rect 7791 17221 7803 17255
rect 7745 17215 7803 17221
rect 7929 17255 7987 17261
rect 7929 17221 7941 17255
rect 7975 17252 7987 17255
rect 7975 17224 8248 17252
rect 7975 17221 7987 17224
rect 7929 17215 7987 17221
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17153 4675 17187
rect 4617 17147 4675 17153
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 5132 17156 5457 17184
rect 5132 17144 5138 17156
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 5445 17147 5503 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 5718 17184 5724 17196
rect 5675 17156 5724 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 5997 17187 6055 17193
rect 5997 17184 6009 17187
rect 5960 17156 6009 17184
rect 5960 17144 5966 17156
rect 5997 17153 6009 17156
rect 6043 17153 6055 17187
rect 5997 17147 6055 17153
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1397 17119 1455 17125
rect 1397 17116 1409 17119
rect 992 17088 1409 17116
rect 992 17076 998 17088
rect 1397 17085 1409 17088
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1670 17076 1676 17128
rect 1728 17076 1734 17128
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17116 4767 17119
rect 4755 17088 6132 17116
rect 4755 17085 4767 17088
rect 4709 17079 4767 17085
rect 6104 16980 6132 17088
rect 6196 17048 6224 17147
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 6328 17156 6377 17184
rect 6328 17144 6334 17156
rect 6365 17153 6377 17156
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6641 17187 6699 17193
rect 6641 17153 6653 17187
rect 6687 17153 6699 17187
rect 7024 17184 7052 17212
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 7024 17156 7389 17184
rect 6641 17147 6699 17153
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7377 17147 7435 17153
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 6656 17116 6684 17147
rect 7466 17144 7472 17196
rect 7524 17144 7530 17196
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 8021 17187 8079 17193
rect 8021 17184 8033 17187
rect 7699 17182 7788 17184
rect 7852 17182 8033 17184
rect 7699 17156 8033 17182
rect 7699 17153 7711 17156
rect 7760 17154 7880 17156
rect 7653 17147 7711 17153
rect 8021 17153 8033 17156
rect 8067 17184 8079 17187
rect 8110 17184 8116 17196
rect 8067 17156 8116 17184
rect 8067 17153 8079 17156
rect 8021 17147 8079 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 6822 17116 6828 17128
rect 6656 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7248 17088 7297 17116
rect 7248 17076 7254 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7484 17116 7512 17144
rect 8220 17116 8248 17224
rect 8389 17187 8447 17193
rect 8389 17153 8401 17187
rect 8435 17184 8447 17187
rect 8573 17187 8631 17193
rect 8435 17156 8524 17184
rect 8435 17153 8447 17156
rect 8389 17147 8447 17153
rect 7484 17088 8248 17116
rect 8496 17116 8524 17156
rect 8573 17153 8585 17187
rect 8619 17184 8631 17187
rect 8680 17184 8708 17280
rect 8619 17156 8708 17184
rect 8619 17153 8631 17156
rect 8573 17147 8631 17153
rect 8754 17144 8760 17196
rect 8812 17184 8818 17196
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 8812 17156 8861 17184
rect 8812 17144 8818 17156
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 8956 17128 8984 17292
rect 9214 17212 9220 17264
rect 9272 17252 9278 17264
rect 9309 17255 9367 17261
rect 9309 17252 9321 17255
rect 9272 17224 9321 17252
rect 9272 17212 9278 17224
rect 9309 17221 9321 17224
rect 9355 17221 9367 17255
rect 9309 17215 9367 17221
rect 9490 17212 9496 17264
rect 9548 17212 9554 17264
rect 9600 17261 9628 17292
rect 9692 17292 10732 17320
rect 9692 17264 9720 17292
rect 9585 17255 9643 17261
rect 9585 17221 9597 17255
rect 9631 17221 9643 17255
rect 9585 17215 9643 17221
rect 9674 17212 9680 17264
rect 9732 17212 9738 17264
rect 9950 17212 9956 17264
rect 10008 17212 10014 17264
rect 10704 17261 10732 17292
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11606 17320 11612 17332
rect 11204 17292 11612 17320
rect 11204 17280 11210 17292
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 13078 17320 13084 17332
rect 12943 17292 13084 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 13780 17292 14381 17320
rect 13780 17280 13786 17292
rect 14369 17289 14381 17292
rect 14415 17289 14427 17323
rect 14369 17283 14427 17289
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 15381 17323 15439 17329
rect 15381 17320 15393 17323
rect 15344 17292 15393 17320
rect 15344 17280 15350 17292
rect 15381 17289 15393 17292
rect 15427 17289 15439 17323
rect 15381 17283 15439 17289
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 16206 17320 16212 17332
rect 15528 17292 16212 17320
rect 15528 17280 15534 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16574 17280 16580 17332
rect 16632 17320 16638 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16632 17292 17141 17320
rect 16632 17280 16638 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 17129 17283 17187 17289
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 20070 17280 20076 17332
rect 20128 17280 20134 17332
rect 22554 17280 22560 17332
rect 22612 17280 22618 17332
rect 24765 17323 24823 17329
rect 24765 17289 24777 17323
rect 24811 17320 24823 17323
rect 25130 17320 25136 17332
rect 24811 17292 25136 17320
rect 24811 17289 24823 17292
rect 24765 17283 24823 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 26694 17280 26700 17332
rect 26752 17280 26758 17332
rect 10689 17255 10747 17261
rect 10689 17221 10701 17255
rect 10735 17252 10747 17255
rect 11330 17252 11336 17264
rect 10735 17224 11336 17252
rect 10735 17221 10747 17224
rect 10689 17215 10747 17221
rect 11330 17212 11336 17224
rect 11388 17252 11394 17264
rect 12253 17255 12311 17261
rect 12253 17252 12265 17255
rect 11388 17224 12265 17252
rect 11388 17212 11394 17224
rect 12253 17221 12265 17224
rect 12299 17252 12311 17255
rect 12526 17252 12532 17264
rect 12299 17224 12532 17252
rect 12299 17221 12311 17224
rect 12253 17215 12311 17221
rect 12526 17212 12532 17224
rect 12584 17252 12590 17264
rect 14001 17255 14059 17261
rect 12584 17224 13308 17252
rect 12584 17212 12590 17224
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9508 17184 9536 17212
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9171 17156 9873 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9968 17184 9996 17212
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 9968 17156 10885 17184
rect 9861 17147 9919 17153
rect 10873 17153 10885 17156
rect 10919 17184 10931 17187
rect 10962 17184 10968 17196
rect 10919 17156 10968 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 11057 17187 11115 17193
rect 11057 17153 11069 17187
rect 11103 17184 11115 17187
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11103 17156 11529 17184
rect 11103 17153 11115 17156
rect 11057 17147 11115 17153
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 8662 17116 8668 17128
rect 8496 17088 8668 17116
rect 7285 17079 7343 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8938 17076 8944 17128
rect 8996 17076 9002 17128
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17116 9091 17119
rect 9306 17116 9312 17128
rect 9079 17088 9312 17116
rect 9079 17085 9091 17088
rect 9033 17079 9091 17085
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 6270 17048 6276 17060
rect 6196 17020 6276 17048
rect 6270 17008 6276 17020
rect 6328 17008 6334 17060
rect 7745 17051 7803 17057
rect 7745 17048 7757 17051
rect 6396 17020 7757 17048
rect 6396 16980 6424 17020
rect 7745 17017 7757 17020
rect 7791 17017 7803 17051
rect 7745 17011 7803 17017
rect 8481 17051 8539 17057
rect 8481 17017 8493 17051
rect 8527 17048 8539 17051
rect 9416 17048 9444 17079
rect 8527 17020 9444 17048
rect 8527 17017 8539 17020
rect 8481 17011 8539 17017
rect 6104 16952 6424 16980
rect 7282 16940 7288 16992
rect 7340 16940 7346 16992
rect 8754 16940 8760 16992
rect 8812 16980 8818 16992
rect 9508 16980 9536 17079
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 10134 17076 10140 17128
rect 10192 17076 10198 17128
rect 10778 17076 10784 17128
rect 10836 17116 10842 17128
rect 11072 17116 11100 17147
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 12434 17193 12440 17196
rect 12400 17187 12440 17193
rect 12400 17153 12412 17187
rect 12492 17184 12498 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12492 17156 13093 17184
rect 12400 17147 12440 17153
rect 12434 17144 12440 17147
rect 12492 17144 12498 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 13170 17144 13176 17196
rect 13228 17144 13234 17196
rect 13280 17193 13308 17224
rect 14001 17221 14013 17255
rect 14047 17252 14059 17255
rect 15746 17252 15752 17264
rect 14047 17224 15752 17252
rect 14047 17221 14059 17224
rect 14001 17215 14059 17221
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 13265 17147 13323 17153
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 10836 17088 11100 17116
rect 10836 17076 10842 17088
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12032 17088 12633 17116
rect 12032 17076 12038 17088
rect 12621 17085 12633 17088
rect 12667 17116 12679 17119
rect 13556 17116 13584 17147
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 13725 17187 13783 17193
rect 13725 17184 13737 17187
rect 13688 17156 13737 17184
rect 13688 17144 13694 17156
rect 13725 17153 13737 17156
rect 13771 17153 13783 17187
rect 13725 17147 13783 17153
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 15304 17193 15332 17224
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 15838 17212 15844 17264
rect 15896 17252 15902 17264
rect 16482 17252 16488 17264
rect 15896 17224 16488 17252
rect 15896 17212 15902 17224
rect 16482 17212 16488 17224
rect 16540 17252 16546 17264
rect 18984 17252 19012 17280
rect 16540 17224 19012 17252
rect 16540 17212 16546 17224
rect 19334 17212 19340 17264
rect 19392 17212 19398 17264
rect 15289 17187 15347 17193
rect 14516 17156 14964 17184
rect 14516 17144 14522 17156
rect 12667 17088 13584 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 14936 17125 14964 17156
rect 15289 17153 15301 17187
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 16022 17144 16028 17196
rect 16080 17184 16086 17196
rect 16117 17187 16175 17193
rect 16117 17184 16129 17187
rect 16080 17156 16129 17184
rect 16080 17144 16086 17156
rect 16117 17153 16129 17156
rect 16163 17184 16175 17187
rect 16390 17184 16396 17196
rect 16163 17156 16396 17184
rect 16163 17153 16175 17156
rect 16117 17147 16175 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17313 17187 17371 17193
rect 17313 17184 17325 17187
rect 17000 17156 17325 17184
rect 17000 17144 17006 17156
rect 17313 17153 17325 17156
rect 17359 17153 17371 17187
rect 17313 17147 17371 17153
rect 17494 17144 17500 17196
rect 17552 17144 17558 17196
rect 20088 17184 20116 17280
rect 24118 17212 24124 17264
rect 24176 17252 24182 17264
rect 24176 17224 25084 17252
rect 24176 17212 24182 17224
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20088 17156 20729 17184
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14608 17088 14841 17116
rect 14608 17076 14614 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17085 17647 17119
rect 17589 17079 17647 17085
rect 18325 17119 18383 17125
rect 18325 17085 18337 17119
rect 18371 17085 18383 17119
rect 18325 17079 18383 17085
rect 10152 17048 10180 17076
rect 11793 17051 11851 17057
rect 11793 17048 11805 17051
rect 10152 17020 11805 17048
rect 11793 17017 11805 17020
rect 11839 17017 11851 17051
rect 11793 17011 11851 17017
rect 12066 17008 12072 17060
rect 12124 17048 12130 17060
rect 17604 17048 17632 17079
rect 18230 17048 18236 17060
rect 12124 17020 18236 17048
rect 12124 17008 12130 17020
rect 18230 17008 18236 17020
rect 18288 17008 18294 17060
rect 8812 16952 9536 16980
rect 8812 16940 8818 16952
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12434 16980 12440 16992
rect 11664 16952 12440 16980
rect 11664 16940 11670 16952
rect 12434 16940 12440 16952
rect 12492 16980 12498 16992
rect 12529 16983 12587 16989
rect 12529 16980 12541 16983
rect 12492 16952 12541 16980
rect 12492 16940 12498 16952
rect 12529 16949 12541 16952
rect 12575 16980 12587 16983
rect 13403 16983 13461 16989
rect 13403 16980 13415 16983
rect 12575 16952 13415 16980
rect 12575 16949 12587 16952
rect 12529 16943 12587 16949
rect 13403 16949 13415 16952
rect 13449 16949 13461 16983
rect 13403 16943 13461 16949
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18340 16980 18368 17079
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 18966 17076 18972 17128
rect 19024 17116 19030 17128
rect 21266 17116 21272 17128
rect 19024 17088 21272 17116
rect 19024 17076 19030 17088
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 22002 17076 22008 17128
rect 22060 17076 22066 17128
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17085 22155 17119
rect 22204 17116 22232 17147
rect 22278 17144 22284 17196
rect 22336 17184 22342 17196
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 22336 17156 22661 17184
rect 22336 17144 22342 17156
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 22738 17144 22744 17196
rect 22796 17184 22802 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 22796 17156 22845 17184
rect 22796 17144 22802 17156
rect 22833 17153 22845 17156
rect 22879 17184 22891 17187
rect 23382 17184 23388 17196
rect 22879 17156 23388 17184
rect 22879 17153 22891 17156
rect 22833 17147 22891 17153
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 23566 17144 23572 17196
rect 23624 17144 23630 17196
rect 24946 17144 24952 17196
rect 25004 17144 25010 17196
rect 25056 17193 25084 17224
rect 25041 17187 25099 17193
rect 25041 17153 25053 17187
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17184 25375 17187
rect 26712 17184 26740 17280
rect 25363 17156 26740 17184
rect 25363 17153 25375 17156
rect 25317 17147 25375 17153
rect 27338 17144 27344 17196
rect 27396 17184 27402 17196
rect 30193 17187 30251 17193
rect 30193 17184 30205 17187
rect 27396 17156 30205 17184
rect 27396 17144 27402 17156
rect 30193 17153 30205 17156
rect 30239 17153 30251 17187
rect 30193 17147 30251 17153
rect 23584 17116 23612 17144
rect 22204 17088 23612 17116
rect 22097 17079 22155 17085
rect 22112 17048 22140 17079
rect 22186 17048 22192 17060
rect 22112 17020 22192 17048
rect 22186 17008 22192 17020
rect 22244 17008 22250 17060
rect 25225 17051 25283 17057
rect 25225 17048 25237 17051
rect 22296 17020 25237 17048
rect 19150 16980 19156 16992
rect 18012 16952 19156 16980
rect 18012 16940 18018 16952
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 20162 16940 20168 16992
rect 20220 16940 20226 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21542 16980 21548 16992
rect 20956 16952 21548 16980
rect 20956 16940 20962 16952
rect 21542 16940 21548 16952
rect 21600 16980 21606 16992
rect 22296 16980 22324 17020
rect 25225 17017 25237 17020
rect 25271 17048 25283 17051
rect 26142 17048 26148 17060
rect 25271 17020 26148 17048
rect 25271 17017 25283 17020
rect 25225 17011 25283 17017
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 30374 17008 30380 17060
rect 30432 17008 30438 17060
rect 21600 16952 22324 16980
rect 21600 16940 21606 16952
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 22741 16983 22799 16989
rect 22741 16980 22753 16983
rect 22428 16952 22753 16980
rect 22428 16940 22434 16952
rect 22741 16949 22753 16952
rect 22787 16949 22799 16983
rect 22741 16943 22799 16949
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 23661 16983 23719 16989
rect 23661 16980 23673 16983
rect 23440 16952 23673 16980
rect 23440 16940 23446 16952
rect 23661 16949 23673 16952
rect 23707 16949 23719 16983
rect 23661 16943 23719 16949
rect 24029 16983 24087 16989
rect 24029 16949 24041 16983
rect 24075 16980 24087 16983
rect 25038 16980 25044 16992
rect 24075 16952 25044 16980
rect 24075 16949 24087 16952
rect 24029 16943 24087 16949
rect 25038 16940 25044 16952
rect 25096 16980 25102 16992
rect 25498 16980 25504 16992
rect 25096 16952 25504 16980
rect 25096 16940 25102 16952
rect 25498 16940 25504 16952
rect 25556 16980 25562 16992
rect 25958 16980 25964 16992
rect 25556 16952 25964 16980
rect 25556 16940 25562 16952
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 1104 16890 30820 16912
rect 1104 16838 4664 16890
rect 4716 16838 4728 16890
rect 4780 16838 4792 16890
rect 4844 16838 4856 16890
rect 4908 16838 4920 16890
rect 4972 16838 12092 16890
rect 12144 16838 12156 16890
rect 12208 16838 12220 16890
rect 12272 16838 12284 16890
rect 12336 16838 12348 16890
rect 12400 16838 19520 16890
rect 19572 16838 19584 16890
rect 19636 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 26948 16890
rect 27000 16838 27012 16890
rect 27064 16838 27076 16890
rect 27128 16838 27140 16890
rect 27192 16838 27204 16890
rect 27256 16838 30820 16890
rect 1104 16816 30820 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1728 16748 2774 16776
rect 1728 16736 1734 16748
rect 2746 16708 2774 16748
rect 6454 16736 6460 16788
rect 6512 16776 6518 16788
rect 6730 16776 6736 16788
rect 6512 16748 6736 16776
rect 6512 16736 6518 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7248 16748 7849 16776
rect 7248 16736 7254 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 8205 16779 8263 16785
rect 8205 16745 8217 16779
rect 8251 16776 8263 16779
rect 8938 16776 8944 16788
rect 8251 16748 8944 16776
rect 8251 16745 8263 16748
rect 8205 16739 8263 16745
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 9030 16736 9036 16788
rect 9088 16736 9094 16788
rect 9122 16736 9128 16788
rect 9180 16736 9186 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 9585 16779 9643 16785
rect 9585 16776 9597 16779
rect 9548 16748 9597 16776
rect 9548 16736 9554 16748
rect 9585 16745 9597 16748
rect 9631 16745 9643 16779
rect 9585 16739 9643 16745
rect 11790 16736 11796 16788
rect 11848 16776 11854 16788
rect 11848 16748 12480 16776
rect 11848 16736 11854 16748
rect 9048 16708 9076 16736
rect 2746 16680 9076 16708
rect 9140 16708 9168 16736
rect 11146 16708 11152 16720
rect 9140 16680 11152 16708
rect 4522 16600 4528 16652
rect 4580 16640 4586 16652
rect 7929 16643 7987 16649
rect 4580 16612 5396 16640
rect 4580 16600 4586 16612
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 5166 16572 5172 16584
rect 1719 16544 5172 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5368 16581 5396 16612
rect 7929 16609 7941 16643
rect 7975 16640 7987 16643
rect 8294 16640 8300 16652
rect 7975 16612 8300 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 8294 16600 8300 16612
rect 8352 16640 8358 16652
rect 9122 16640 9128 16652
rect 8352 16612 9128 16640
rect 8352 16600 8358 16612
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9766 16640 9772 16652
rect 9508 16612 9772 16640
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 9508 16581 9536 16612
rect 9766 16600 9772 16612
rect 9824 16640 9830 16652
rect 10318 16640 10324 16652
rect 9824 16612 10324 16640
rect 9824 16600 9830 16612
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10888 16649 10916 16680
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 12452 16717 12480 16748
rect 12618 16736 12624 16788
rect 12676 16776 12682 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12676 16748 12909 16776
rect 12676 16736 12682 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 13078 16736 13084 16788
rect 13136 16736 13142 16788
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 19242 16776 19248 16788
rect 15620 16748 19248 16776
rect 15620 16736 15626 16748
rect 19242 16736 19248 16748
rect 19300 16736 19306 16788
rect 19334 16736 19340 16788
rect 19392 16736 19398 16788
rect 19886 16776 19892 16788
rect 19720 16748 19892 16776
rect 12437 16711 12495 16717
rect 12437 16677 12449 16711
rect 12483 16677 12495 16711
rect 12437 16671 12495 16677
rect 18598 16668 18604 16720
rect 18656 16708 18662 16720
rect 19521 16711 19579 16717
rect 19521 16708 19533 16711
rect 18656 16680 19533 16708
rect 18656 16668 18662 16680
rect 19521 16677 19533 16680
rect 19567 16677 19579 16711
rect 19521 16671 19579 16677
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10612 16612 10701 16640
rect 7837 16575 7895 16581
rect 7837 16572 7849 16575
rect 7524 16544 7849 16572
rect 7524 16532 7530 16544
rect 7837 16541 7849 16544
rect 7883 16541 7895 16575
rect 7837 16535 7895 16541
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 9677 16575 9735 16581
rect 9677 16541 9689 16575
rect 9723 16572 9735 16575
rect 10410 16572 10416 16584
rect 9723 16544 10416 16572
rect 9723 16541 9735 16544
rect 9677 16535 9735 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 10502 16532 10508 16584
rect 10560 16532 10566 16584
rect 3418 16464 3424 16516
rect 3476 16504 3482 16516
rect 10520 16504 10548 16532
rect 3476 16476 10548 16504
rect 10612 16504 10640 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16609 10931 16643
rect 10873 16603 10931 16609
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 17957 16643 18015 16649
rect 11112 16612 12020 16640
rect 11112 16600 11118 16612
rect 10778 16581 10784 16584
rect 10770 16575 10784 16581
rect 10770 16541 10782 16575
rect 10836 16572 10842 16584
rect 11072 16572 11100 16600
rect 11992 16584 12020 16612
rect 17957 16609 17969 16643
rect 18003 16609 18015 16643
rect 18690 16640 18696 16652
rect 17957 16603 18015 16609
rect 18432 16612 18696 16640
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10836 16544 10870 16572
rect 11072 16544 11161 16572
rect 10770 16535 10784 16541
rect 10778 16532 10784 16535
rect 10836 16532 10842 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 11241 16507 11299 16513
rect 11241 16504 11253 16507
rect 10612 16476 11253 16504
rect 3476 16464 3482 16476
rect 11241 16473 11253 16476
rect 11287 16473 11299 16507
rect 11241 16467 11299 16473
rect 11348 16448 11376 16535
rect 11974 16532 11980 16584
rect 12032 16532 12038 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12434 16572 12440 16584
rect 12391 16544 12440 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 12434 16532 12440 16544
rect 12492 16532 12498 16584
rect 12526 16532 12532 16584
rect 12584 16532 12590 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 15344 16544 16957 16572
rect 15344 16532 15350 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 17865 16535 17923 16541
rect 12805 16507 12863 16513
rect 12805 16473 12817 16507
rect 12851 16473 12863 16507
rect 12805 16467 12863 16473
rect 13065 16507 13123 16513
rect 13065 16473 13077 16507
rect 13111 16504 13123 16507
rect 13170 16504 13176 16516
rect 13111 16476 13176 16504
rect 13111 16473 13123 16476
rect 13065 16467 13123 16473
rect 934 16396 940 16448
rect 992 16436 998 16448
rect 1489 16439 1547 16445
rect 1489 16436 1501 16439
rect 992 16408 1501 16436
rect 992 16396 998 16408
rect 1489 16405 1501 16408
rect 1535 16405 1547 16439
rect 1489 16399 1547 16405
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 4488 16408 5273 16436
rect 4488 16396 4494 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 10502 16396 10508 16448
rect 10560 16396 10566 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 12820 16436 12848 16467
rect 13170 16464 13176 16476
rect 13228 16464 13234 16516
rect 13265 16507 13323 16513
rect 13265 16473 13277 16507
rect 13311 16504 13323 16507
rect 13722 16504 13728 16516
rect 13311 16476 13728 16504
rect 13311 16473 13323 16476
rect 13265 16467 13323 16473
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 13814 16464 13820 16516
rect 13872 16464 13878 16516
rect 14274 16464 14280 16516
rect 14332 16464 14338 16516
rect 14826 16464 14832 16516
rect 14884 16504 14890 16516
rect 15010 16504 15016 16516
rect 14884 16476 15016 16504
rect 14884 16464 14890 16476
rect 15010 16464 15016 16476
rect 15068 16504 15074 16516
rect 17880 16504 17908 16535
rect 15068 16476 17908 16504
rect 17972 16504 18000 16603
rect 18432 16581 18460 16612
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 18966 16640 18972 16652
rect 18800 16612 18972 16640
rect 18800 16581 18828 16612
rect 18966 16600 18972 16612
rect 19024 16600 19030 16652
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19116 16612 19288 16640
rect 19116 16600 19122 16612
rect 19260 16581 19288 16612
rect 19720 16581 19748 16748
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 21499 16779 21557 16785
rect 21499 16776 21511 16779
rect 20772 16748 21511 16776
rect 20772 16736 20778 16748
rect 21499 16745 21511 16748
rect 21545 16745 21557 16779
rect 21499 16739 21557 16745
rect 21637 16779 21695 16785
rect 21637 16745 21649 16779
rect 21683 16776 21695 16779
rect 22738 16776 22744 16788
rect 21683 16748 22744 16776
rect 21683 16745 21695 16748
rect 21637 16739 21695 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 22888 16748 24900 16776
rect 22888 16736 22894 16748
rect 20349 16711 20407 16717
rect 20349 16708 20361 16711
rect 19812 16680 20361 16708
rect 19812 16581 19840 16680
rect 20349 16677 20361 16680
rect 20395 16677 20407 16711
rect 20898 16708 20904 16720
rect 20349 16671 20407 16677
rect 20548 16680 20904 16708
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20548 16640 20576 16680
rect 20898 16668 20904 16680
rect 20956 16668 20962 16720
rect 20990 16668 20996 16720
rect 21048 16668 21054 16720
rect 23385 16711 23443 16717
rect 21100 16680 23060 16708
rect 20036 16612 20576 16640
rect 20036 16600 20042 16612
rect 20622 16600 20628 16652
rect 20680 16600 20686 16652
rect 20717 16643 20775 16649
rect 20717 16609 20729 16643
rect 20763 16640 20775 16643
rect 21100 16640 21128 16680
rect 20763 16612 21128 16640
rect 20763 16609 20775 16612
rect 20717 16603 20775 16609
rect 20916 16584 20944 16612
rect 21726 16600 21732 16652
rect 21784 16600 21790 16652
rect 22097 16643 22155 16649
rect 22097 16609 22109 16643
rect 22143 16640 22155 16643
rect 22922 16640 22928 16652
rect 22143 16612 22928 16640
rect 22143 16609 22155 16612
rect 22097 16603 22155 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 23032 16640 23060 16680
rect 23385 16677 23397 16711
rect 23431 16708 23443 16711
rect 23431 16680 23888 16708
rect 23431 16677 23443 16680
rect 23385 16671 23443 16677
rect 23860 16649 23888 16680
rect 24118 16668 24124 16720
rect 24176 16668 24182 16720
rect 24872 16708 24900 16748
rect 25590 16736 25596 16788
rect 25648 16736 25654 16788
rect 26326 16776 26332 16788
rect 26160 16748 26332 16776
rect 24872 16680 25176 16708
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23032 16612 23765 16640
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23845 16643 23903 16649
rect 23845 16609 23857 16643
rect 23891 16609 23903 16643
rect 23845 16603 23903 16609
rect 24872 16584 24900 16680
rect 25038 16640 25044 16652
rect 24964 16612 25044 16640
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16541 18475 16575
rect 18417 16535 18475 16541
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 20073 16575 20131 16581
rect 20073 16541 20085 16575
rect 20119 16572 20131 16575
rect 20162 16572 20168 16584
rect 20119 16544 20168 16572
rect 20119 16541 20131 16544
rect 20073 16535 20131 16541
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20530 16532 20536 16584
rect 20588 16532 20594 16584
rect 20806 16532 20812 16584
rect 20864 16532 20870 16584
rect 20898 16532 20904 16584
rect 20956 16532 20962 16584
rect 22186 16532 22192 16584
rect 22244 16532 22250 16584
rect 22370 16532 22376 16584
rect 22428 16532 22434 16584
rect 22646 16532 22652 16584
rect 22704 16581 22710 16584
rect 22704 16575 22733 16581
rect 22721 16541 22733 16575
rect 22704 16535 22733 16541
rect 22704 16532 22710 16535
rect 22830 16532 22836 16584
rect 22888 16532 22894 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 23934 16532 23940 16584
rect 23992 16532 23998 16584
rect 24670 16572 24676 16584
rect 24044 16544 24676 16572
rect 19058 16504 19064 16516
rect 17972 16476 19064 16504
rect 15068 16464 15074 16476
rect 19058 16464 19064 16476
rect 19116 16504 19122 16516
rect 20824 16504 20852 16532
rect 19116 16476 20852 16504
rect 21177 16507 21235 16513
rect 19116 16464 19122 16476
rect 21177 16473 21189 16507
rect 21223 16504 21235 16507
rect 21361 16507 21419 16513
rect 21361 16504 21373 16507
rect 21223 16476 21373 16504
rect 21223 16473 21235 16476
rect 21177 16467 21235 16473
rect 21361 16473 21373 16476
rect 21407 16473 21419 16507
rect 21361 16467 21419 16473
rect 13354 16436 13360 16448
rect 12820 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16436 13418 16448
rect 13541 16439 13599 16445
rect 13541 16436 13553 16439
rect 13412 16408 13553 16436
rect 13412 16396 13418 16408
rect 13541 16405 13553 16408
rect 13587 16405 13599 16439
rect 13541 16399 13599 16405
rect 17034 16396 17040 16448
rect 17092 16396 17098 16448
rect 21376 16436 21404 16467
rect 22462 16464 22468 16516
rect 22520 16464 22526 16516
rect 22554 16464 22560 16516
rect 22612 16464 22618 16516
rect 24044 16436 24072 16544
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 24854 16532 24860 16584
rect 24912 16532 24918 16584
rect 24964 16581 24992 16612
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 25148 16640 25176 16680
rect 25682 16668 25688 16720
rect 25740 16708 25746 16720
rect 26160 16717 26188 16748
rect 26326 16736 26332 16748
rect 26384 16776 26390 16788
rect 26384 16748 27016 16776
rect 26384 16736 26390 16748
rect 26145 16711 26203 16717
rect 25740 16680 26096 16708
rect 25740 16668 25746 16680
rect 25409 16643 25467 16649
rect 25409 16640 25421 16643
rect 25148 16612 25421 16640
rect 25409 16609 25421 16612
rect 25455 16609 25467 16643
rect 25409 16603 25467 16609
rect 25498 16600 25504 16652
rect 25556 16600 25562 16652
rect 25961 16643 26019 16649
rect 25961 16640 25973 16643
rect 25792 16612 25973 16640
rect 25792 16584 25820 16612
rect 25961 16609 25973 16612
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 25130 16532 25136 16584
rect 25188 16532 25194 16584
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 25774 16532 25780 16584
rect 25832 16532 25838 16584
rect 26068 16572 26096 16680
rect 26145 16677 26157 16711
rect 26191 16677 26203 16711
rect 26605 16711 26663 16717
rect 26605 16708 26617 16711
rect 26145 16671 26203 16677
rect 26436 16680 26617 16708
rect 26436 16652 26464 16680
rect 26605 16677 26617 16680
rect 26651 16677 26663 16711
rect 26605 16671 26663 16677
rect 26418 16600 26424 16652
rect 26476 16600 26482 16652
rect 26988 16649 27016 16748
rect 26513 16643 26571 16649
rect 26513 16609 26525 16643
rect 26559 16609 26571 16643
rect 26513 16603 26571 16609
rect 26973 16643 27031 16649
rect 26973 16609 26985 16643
rect 27019 16640 27031 16643
rect 27338 16640 27344 16652
rect 27019 16612 27344 16640
rect 27019 16609 27031 16612
rect 26973 16603 27031 16609
rect 26528 16572 26556 16603
rect 27338 16600 27344 16612
rect 27396 16600 27402 16652
rect 26068 16544 26556 16572
rect 30469 16575 30527 16581
rect 30469 16541 30481 16575
rect 30515 16572 30527 16575
rect 30515 16544 30972 16572
rect 30515 16541 30527 16544
rect 30469 16535 30527 16541
rect 30944 16516 30972 16544
rect 25884 16476 30328 16504
rect 21376 16408 24072 16436
rect 24670 16396 24676 16448
rect 24728 16396 24734 16448
rect 24762 16396 24768 16448
rect 24820 16436 24826 16448
rect 25884 16436 25912 16476
rect 30300 16445 30328 16476
rect 30926 16464 30932 16516
rect 30984 16464 30990 16516
rect 24820 16408 25912 16436
rect 30285 16439 30343 16445
rect 24820 16396 24826 16408
rect 30285 16405 30297 16439
rect 30331 16405 30343 16439
rect 30285 16399 30343 16405
rect 1104 16346 30820 16368
rect 1104 16294 5324 16346
rect 5376 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 12752 16346
rect 12804 16294 12816 16346
rect 12868 16294 12880 16346
rect 12932 16294 12944 16346
rect 12996 16294 13008 16346
rect 13060 16294 20180 16346
rect 20232 16294 20244 16346
rect 20296 16294 20308 16346
rect 20360 16294 20372 16346
rect 20424 16294 20436 16346
rect 20488 16294 27608 16346
rect 27660 16294 27672 16346
rect 27724 16294 27736 16346
rect 27788 16294 27800 16346
rect 27852 16294 27864 16346
rect 27916 16294 30820 16346
rect 1104 16272 30820 16294
rect 4430 16192 4436 16244
rect 4488 16192 4494 16244
rect 5166 16192 5172 16244
rect 5224 16192 5230 16244
rect 5442 16192 5448 16244
rect 5500 16232 5506 16244
rect 6086 16232 6092 16244
rect 5500 16204 6092 16232
rect 5500 16192 5506 16204
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 7466 16192 7472 16244
rect 7524 16192 7530 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 9272 16204 9536 16232
rect 9272 16192 9278 16204
rect 4448 16164 4476 16192
rect 4370 16136 4476 16164
rect 5184 16164 5212 16192
rect 5184 16136 9260 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1688 16028 1716 16059
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6086 16056 6092 16108
rect 6144 16056 6150 16108
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16065 7067 16099
rect 7009 16059 7067 16065
rect 3329 16031 3387 16037
rect 3329 16028 3341 16031
rect 1688 16000 3341 16028
rect 3329 15997 3341 16000
rect 3375 15997 3387 16031
rect 3329 15991 3387 15997
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 1489 15895 1547 15901
rect 1489 15892 1501 15895
rect 992 15864 1501 15892
rect 992 15852 998 15864
rect 1489 15861 1501 15864
rect 1535 15861 1547 15895
rect 3344 15892 3372 15991
rect 4430 15988 4436 16040
rect 4488 16028 4494 16040
rect 4801 16031 4859 16037
rect 4801 16028 4813 16031
rect 4488 16000 4813 16028
rect 4488 15988 4494 16000
rect 4801 15997 4813 16000
rect 4847 15997 4859 16031
rect 4801 15991 4859 15997
rect 5074 15988 5080 16040
rect 5132 15988 5138 16040
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 6270 16028 6276 16040
rect 5767 16000 6276 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 5736 15960 5764 15991
rect 6270 15988 6276 16000
rect 6328 16028 6334 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 6328 16000 6377 16028
rect 6328 15988 6334 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 7024 15972 7052 16059
rect 9232 16028 9260 16136
rect 9508 16105 9536 16204
rect 10502 16192 10508 16244
rect 10560 16192 10566 16244
rect 11974 16192 11980 16244
rect 12032 16192 12038 16244
rect 17862 16232 17868 16244
rect 16684 16204 17868 16232
rect 10520 16164 10548 16192
rect 9600 16136 10548 16164
rect 9600 16105 9628 16136
rect 11422 16124 11428 16176
rect 11480 16164 11486 16176
rect 11606 16164 11612 16176
rect 11480 16136 11612 16164
rect 11480 16124 11486 16136
rect 11606 16124 11612 16136
rect 11664 16164 11670 16176
rect 11664 16136 11928 16164
rect 11664 16124 11670 16136
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9907 16068 10333 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10468 16068 11560 16096
rect 10468 16056 10474 16068
rect 10778 16028 10784 16040
rect 9232 16000 10784 16028
rect 10778 15988 10784 16000
rect 10836 16028 10842 16040
rect 11532 16037 11560 16068
rect 10873 16031 10931 16037
rect 10873 16028 10885 16031
rect 10836 16000 10885 16028
rect 10836 15988 10842 16000
rect 10873 15997 10885 16000
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 15997 11575 16031
rect 11900 16028 11928 16136
rect 11992 16105 12020 16192
rect 13909 16167 13967 16173
rect 13909 16164 13921 16167
rect 12406 16136 13921 16164
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12406 16028 12434 16136
rect 13909 16133 13921 16136
rect 13955 16133 13967 16167
rect 13909 16127 13967 16133
rect 14200 16136 15056 16164
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 13630 16096 13636 16108
rect 13587 16068 13636 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 13630 16056 13636 16068
rect 13688 16096 13694 16108
rect 14200 16105 14228 16136
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13688 16068 14197 16096
rect 13688 16056 13694 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16096 14703 16099
rect 14826 16096 14832 16108
rect 14691 16068 14832 16096
rect 14691 16065 14703 16068
rect 14645 16059 14703 16065
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 15028 16105 15056 16136
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16065 15071 16099
rect 15838 16096 15844 16108
rect 15013 16059 15071 16065
rect 15120 16068 15844 16096
rect 11900 16000 12434 16028
rect 11517 15991 11575 15997
rect 5092 15932 5764 15960
rect 5092 15892 5120 15932
rect 5902 15920 5908 15972
rect 5960 15960 5966 15972
rect 6641 15963 6699 15969
rect 6641 15960 6653 15963
rect 5960 15932 6653 15960
rect 5960 15920 5966 15932
rect 6641 15929 6653 15932
rect 6687 15929 6699 15963
rect 6641 15923 6699 15929
rect 7006 15920 7012 15972
rect 7064 15920 7070 15972
rect 7377 15963 7435 15969
rect 7377 15929 7389 15963
rect 7423 15960 7435 15963
rect 7466 15960 7472 15972
rect 7423 15932 7472 15960
rect 7423 15929 7435 15932
rect 7377 15923 7435 15929
rect 7466 15920 7472 15932
rect 7524 15920 7530 15972
rect 9769 15963 9827 15969
rect 9769 15929 9781 15963
rect 9815 15960 9827 15963
rect 10686 15960 10692 15972
rect 9815 15932 10692 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 3344 15864 5120 15892
rect 5169 15895 5227 15901
rect 1489 15855 1547 15861
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5350 15892 5356 15904
rect 5215 15864 5356 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 5994 15852 6000 15904
rect 6052 15852 6058 15904
rect 6825 15895 6883 15901
rect 6825 15861 6837 15895
rect 6871 15892 6883 15895
rect 7190 15892 7196 15904
rect 6871 15864 7196 15892
rect 6871 15861 6883 15864
rect 6825 15855 6883 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 9306 15852 9312 15904
rect 9364 15852 9370 15904
rect 10888 15892 10916 15991
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 14936 16028 14964 16059
rect 15120 16028 15148 16068
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 16022 16056 16028 16108
rect 16080 16056 16086 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16574 16096 16580 16108
rect 16163 16068 16580 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 16684 16105 16712 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 18693 16235 18751 16241
rect 18693 16232 18705 16235
rect 18288 16204 18705 16232
rect 18288 16192 18294 16204
rect 18693 16201 18705 16204
rect 18739 16201 18751 16235
rect 18693 16195 18751 16201
rect 20530 16192 20536 16244
rect 20588 16192 20594 16244
rect 20714 16192 20720 16244
rect 20772 16192 20778 16244
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21140 16204 22324 16232
rect 21140 16192 21146 16204
rect 17034 16124 17040 16176
rect 17092 16164 17098 16176
rect 20732 16164 20760 16192
rect 22296 16176 22324 16204
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 22741 16235 22799 16241
rect 22741 16232 22753 16235
rect 22520 16204 22753 16232
rect 22520 16192 22526 16204
rect 22741 16201 22753 16204
rect 22787 16201 22799 16235
rect 22741 16195 22799 16201
rect 23569 16235 23627 16241
rect 23569 16201 23581 16235
rect 23615 16232 23627 16235
rect 23934 16232 23940 16244
rect 23615 16204 23940 16232
rect 23615 16201 23627 16204
rect 23569 16195 23627 16201
rect 20901 16167 20959 16173
rect 20901 16164 20913 16167
rect 17092 16136 17434 16164
rect 20548 16136 20913 16164
rect 17092 16124 17098 16136
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 18969 16099 19027 16105
rect 18969 16065 18981 16099
rect 19015 16096 19027 16099
rect 19058 16096 19064 16108
rect 19015 16068 19064 16096
rect 19015 16065 19027 16068
rect 18969 16059 19027 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20548 16105 20576 16136
rect 20901 16133 20913 16136
rect 20947 16133 20959 16167
rect 20901 16127 20959 16133
rect 20990 16124 20996 16176
rect 21048 16124 21054 16176
rect 21726 16124 21732 16176
rect 21784 16124 21790 16176
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 22373 16167 22431 16173
rect 22373 16164 22385 16167
rect 22336 16136 22385 16164
rect 22336 16124 22342 16136
rect 22373 16133 22385 16136
rect 22419 16133 22431 16167
rect 22373 16127 22431 16133
rect 22557 16167 22615 16173
rect 22557 16133 22569 16167
rect 22603 16164 22615 16167
rect 22646 16164 22652 16176
rect 22603 16136 22652 16164
rect 22603 16133 22615 16136
rect 22557 16127 22615 16133
rect 22646 16124 22652 16136
rect 22704 16124 22710 16176
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16096 20775 16099
rect 21008 16096 21036 16124
rect 20763 16068 21036 16096
rect 20763 16065 20775 16068
rect 20717 16059 20775 16065
rect 14936 16000 15148 16028
rect 15286 15988 15292 16040
rect 15344 15988 15350 16040
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15488 16000 16221 16028
rect 11422 15920 11428 15972
rect 11480 15960 11486 15972
rect 13814 15960 13820 15972
rect 11480 15932 13820 15960
rect 11480 15920 11486 15932
rect 13814 15920 13820 15932
rect 13872 15960 13878 15972
rect 14829 15963 14887 15969
rect 14829 15960 14841 15963
rect 13872 15932 14841 15960
rect 13872 15920 13878 15932
rect 14829 15929 14841 15932
rect 14875 15960 14887 15963
rect 14918 15960 14924 15972
rect 14875 15932 14924 15960
rect 14875 15929 14887 15932
rect 14829 15923 14887 15929
rect 14918 15920 14924 15932
rect 14976 15960 14982 15972
rect 15378 15960 15384 15972
rect 14976 15932 15384 15960
rect 14976 15920 14982 15932
rect 15378 15920 15384 15932
rect 15436 15920 15442 15972
rect 11701 15895 11759 15901
rect 11701 15892 11713 15895
rect 10888 15864 11713 15892
rect 11701 15861 11713 15864
rect 11747 15861 11759 15895
rect 11701 15855 11759 15861
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 13688 15864 14473 15892
rect 13688 15852 13694 15864
rect 14461 15861 14473 15864
rect 14507 15892 14519 15895
rect 15488 15892 15516 16000
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 14507 15864 15516 15892
rect 14507 15861 14519 15864
rect 14461 15855 14519 15861
rect 15654 15852 15660 15904
rect 15712 15852 15718 15904
rect 16224 15892 16252 15991
rect 16942 15988 16948 16040
rect 17000 15988 17006 16040
rect 20364 16028 20392 16059
rect 20732 16028 20760 16059
rect 20364 16000 20760 16028
rect 21744 16028 21772 16124
rect 22756 16096 22784 16195
rect 23934 16192 23940 16204
rect 23992 16192 23998 16244
rect 24486 16192 24492 16244
rect 24544 16192 24550 16244
rect 24791 16235 24849 16241
rect 24791 16201 24803 16235
rect 24837 16232 24849 16235
rect 25590 16232 25596 16244
rect 24837 16204 25596 16232
rect 24837 16201 24849 16204
rect 24791 16195 24849 16201
rect 25590 16192 25596 16204
rect 25648 16192 25654 16244
rect 25774 16192 25780 16244
rect 25832 16192 25838 16244
rect 26326 16192 26332 16244
rect 26384 16192 26390 16244
rect 24394 16164 24400 16176
rect 23584 16136 24400 16164
rect 23584 16105 23612 16136
rect 24394 16124 24400 16136
rect 24452 16124 24458 16176
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22756 16068 23397 16096
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 24504 16096 24532 16192
rect 24581 16167 24639 16173
rect 24581 16133 24593 16167
rect 24627 16164 24639 16167
rect 24627 16136 24808 16164
rect 24627 16133 24639 16136
rect 24581 16127 24639 16133
rect 24780 16108 24808 16136
rect 25130 16124 25136 16176
rect 25188 16164 25194 16176
rect 25792 16164 25820 16192
rect 25188 16136 25820 16164
rect 25188 16124 25194 16136
rect 23891 16068 24532 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 23584 16028 23612 16059
rect 24762 16056 24768 16108
rect 24820 16056 24826 16108
rect 25222 16056 25228 16108
rect 25280 16096 25286 16108
rect 25682 16096 25688 16108
rect 25280 16068 25688 16096
rect 25280 16056 25286 16068
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 26344 16105 26372 16192
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 30193 16099 30251 16105
rect 30193 16065 30205 16099
rect 30239 16065 30251 16099
rect 30193 16059 30251 16065
rect 30208 16028 30236 16059
rect 21744 16000 23612 16028
rect 24136 16000 30236 16028
rect 18414 15920 18420 15972
rect 18472 15960 18478 15972
rect 24136 15960 24164 16000
rect 18472 15932 24164 15960
rect 18472 15920 18478 15932
rect 24946 15920 24952 15972
rect 25004 15920 25010 15972
rect 17678 15892 17684 15904
rect 16224 15864 17684 15892
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 21082 15892 21088 15904
rect 20772 15864 21088 15892
rect 20772 15852 20778 15864
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 23750 15852 23756 15904
rect 23808 15852 23814 15904
rect 24670 15852 24676 15904
rect 24728 15892 24734 15904
rect 24765 15895 24823 15901
rect 24765 15892 24777 15895
rect 24728 15864 24777 15892
rect 24728 15852 24734 15864
rect 24765 15861 24777 15864
rect 24811 15861 24823 15895
rect 24765 15855 24823 15861
rect 25130 15852 25136 15904
rect 25188 15892 25194 15904
rect 25774 15892 25780 15904
rect 25188 15864 25780 15892
rect 25188 15852 25194 15864
rect 25774 15852 25780 15864
rect 25832 15852 25838 15904
rect 25866 15852 25872 15904
rect 25924 15852 25930 15904
rect 26237 15895 26295 15901
rect 26237 15861 26249 15895
rect 26283 15892 26295 15895
rect 26418 15892 26424 15904
rect 26283 15864 26424 15892
rect 26283 15861 26295 15864
rect 26237 15855 26295 15861
rect 26418 15852 26424 15864
rect 26476 15852 26482 15904
rect 30374 15852 30380 15904
rect 30432 15852 30438 15904
rect 1104 15802 30820 15824
rect 1104 15750 4664 15802
rect 4716 15750 4728 15802
rect 4780 15750 4792 15802
rect 4844 15750 4856 15802
rect 4908 15750 4920 15802
rect 4972 15750 12092 15802
rect 12144 15750 12156 15802
rect 12208 15750 12220 15802
rect 12272 15750 12284 15802
rect 12336 15750 12348 15802
rect 12400 15750 19520 15802
rect 19572 15750 19584 15802
rect 19636 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 26948 15802
rect 27000 15750 27012 15802
rect 27064 15750 27076 15802
rect 27128 15750 27140 15802
rect 27192 15750 27204 15802
rect 27256 15750 30820 15802
rect 1104 15728 30820 15750
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4488 15660 4721 15688
rect 4488 15648 4494 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 5169 15691 5227 15697
rect 5169 15688 5181 15691
rect 4948 15660 5181 15688
rect 4948 15648 4954 15660
rect 5169 15657 5181 15660
rect 5215 15688 5227 15691
rect 5442 15688 5448 15700
rect 5215 15660 5448 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5994 15688 6000 15700
rect 5552 15660 6000 15688
rect 1581 15623 1639 15629
rect 1581 15589 1593 15623
rect 1627 15620 1639 15623
rect 1627 15592 5488 15620
rect 1627 15589 1639 15592
rect 1581 15583 1639 15589
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 4893 15447 4951 15453
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 4908 15348 4936 15447
rect 5000 15416 5028 15447
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 5368 15416 5396 15515
rect 5000 15388 5396 15416
rect 5460 15416 5488 15592
rect 5552 15561 5580 15660
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6270 15648 6276 15700
rect 6328 15648 6334 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 9306 15697 9312 15700
rect 9296 15691 9312 15697
rect 7984 15660 8156 15688
rect 7984 15648 7990 15660
rect 5810 15580 5816 15632
rect 5868 15580 5874 15632
rect 6288 15620 6316 15648
rect 6365 15623 6423 15629
rect 6365 15620 6377 15623
rect 6288 15592 6377 15620
rect 6365 15589 6377 15592
rect 6411 15589 6423 15623
rect 6365 15583 6423 15589
rect 7561 15623 7619 15629
rect 7561 15589 7573 15623
rect 7607 15620 7619 15623
rect 7607 15592 8064 15620
rect 7607 15589 7619 15592
rect 7561 15583 7619 15589
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15521 5595 15555
rect 5828 15552 5856 15580
rect 5537 15515 5595 15521
rect 5736 15524 5856 15552
rect 6457 15555 6515 15561
rect 5626 15444 5632 15496
rect 5684 15444 5690 15496
rect 5736 15493 5764 15524
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 6457 15515 6515 15521
rect 6932 15524 7665 15552
rect 5721 15487 5779 15493
rect 5721 15453 5733 15487
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5859 15456 6408 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 6380 15428 6408 15456
rect 5994 15416 6000 15428
rect 5460 15388 6000 15416
rect 5994 15376 6000 15388
rect 6052 15376 6058 15428
rect 6362 15376 6368 15428
rect 6420 15376 6426 15428
rect 6472 15416 6500 15515
rect 6932 15493 6960 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7653 15515 7711 15521
rect 7760 15524 7941 15552
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 6917 15447 6975 15453
rect 7006 15444 7012 15496
rect 7064 15444 7070 15496
rect 7098 15444 7104 15496
rect 7156 15444 7162 15496
rect 7190 15444 7196 15496
rect 7248 15444 7254 15496
rect 7466 15444 7472 15496
rect 7524 15484 7530 15496
rect 7760 15484 7788 15524
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8036 15496 8064 15592
rect 7524 15456 7788 15484
rect 7837 15487 7895 15493
rect 7524 15444 7530 15456
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7024 15416 7052 15444
rect 7377 15419 7435 15425
rect 7377 15416 7389 15419
rect 6472 15388 7389 15416
rect 7377 15385 7389 15388
rect 7423 15385 7435 15419
rect 7852 15416 7880 15447
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8128 15493 8156 15660
rect 9296 15657 9308 15691
rect 9296 15651 9312 15657
rect 9306 15648 9312 15651
rect 9364 15648 9370 15700
rect 10318 15648 10324 15700
rect 10376 15688 10382 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 10376 15660 10885 15688
rect 10376 15648 10382 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 10873 15651 10931 15657
rect 11054 15648 11060 15700
rect 11112 15648 11118 15700
rect 15654 15648 15660 15700
rect 15712 15648 15718 15700
rect 18414 15648 18420 15700
rect 18472 15648 18478 15700
rect 24854 15648 24860 15700
rect 24912 15688 24918 15700
rect 25130 15688 25136 15700
rect 24912 15660 25136 15688
rect 24912 15648 24918 15660
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 25314 15648 25320 15700
rect 25372 15688 25378 15700
rect 25685 15691 25743 15697
rect 25685 15688 25697 15691
rect 25372 15660 25697 15688
rect 25372 15648 25378 15660
rect 25685 15657 25697 15660
rect 25731 15657 25743 15691
rect 25685 15651 25743 15657
rect 25866 15648 25872 15700
rect 25924 15648 25930 15700
rect 10778 15580 10784 15632
rect 10836 15580 10842 15632
rect 13722 15620 13728 15632
rect 13096 15592 13728 15620
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15552 9091 15555
rect 9306 15552 9312 15564
rect 9079 15524 9312 15552
rect 9079 15521 9091 15524
rect 9033 15515 9091 15521
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 10796 15484 10824 15580
rect 11793 15555 11851 15561
rect 11793 15552 11805 15555
rect 11532 15524 11805 15552
rect 11532 15496 11560 15524
rect 11793 15521 11805 15524
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 13096 15552 13124 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 14185 15555 14243 15561
rect 14185 15552 14197 15555
rect 12584 15524 13124 15552
rect 13556 15524 14197 15552
rect 12584 15512 12590 15524
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 8159 15456 9076 15484
rect 10796 15456 11345 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 7852 15388 8156 15416
rect 7377 15379 7435 15385
rect 8128 15360 8156 15388
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 4908 15320 7021 15348
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 8110 15308 8116 15360
rect 8168 15308 8174 15360
rect 9048 15348 9076 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11514 15444 11520 15496
rect 11572 15444 11578 15496
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 10534 15388 11376 15416
rect 11238 15348 11244 15360
rect 9048 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 11348 15348 11376 15388
rect 12066 15376 12072 15428
rect 12124 15376 12130 15428
rect 12618 15376 12624 15428
rect 12676 15376 12682 15428
rect 13556 15360 13584 15524
rect 14185 15521 14197 15524
rect 14231 15521 14243 15555
rect 14185 15515 14243 15521
rect 14642 15512 14648 15564
rect 14700 15512 14706 15564
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15484 14335 15487
rect 14734 15484 14740 15496
rect 14323 15456 14740 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 14734 15444 14740 15456
rect 14792 15484 14798 15496
rect 15102 15484 15108 15496
rect 14792 15456 15108 15484
rect 14792 15444 14798 15456
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 15672 15484 15700 15648
rect 16022 15580 16028 15632
rect 16080 15620 16086 15632
rect 18432 15620 18460 15648
rect 16080 15592 18460 15620
rect 16080 15580 16086 15592
rect 17052 15561 17080 15592
rect 23750 15580 23756 15632
rect 23808 15580 23814 15632
rect 25884 15620 25912 15648
rect 25608 15592 25912 15620
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17310 15512 17316 15564
rect 17368 15512 17374 15564
rect 15427 15456 15700 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 16666 15444 16672 15496
rect 16724 15484 16730 15496
rect 16945 15487 17003 15493
rect 16945 15484 16957 15487
rect 16724 15456 16957 15484
rect 16724 15444 16730 15456
rect 16945 15453 16957 15456
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 18874 15444 18880 15496
rect 18932 15444 18938 15496
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21266 15484 21272 15496
rect 21039 15456 21272 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 22278 15444 22284 15496
rect 22336 15444 22342 15496
rect 23768 15484 23796 15580
rect 25608 15552 25636 15592
rect 25056 15524 25268 15552
rect 25056 15496 25084 15524
rect 23690 15456 23796 15484
rect 25038 15444 25044 15496
rect 25096 15444 25102 15496
rect 25130 15444 25136 15496
rect 25188 15444 25194 15496
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 20898 15416 20904 15428
rect 13780 15388 20904 15416
rect 13780 15376 13786 15388
rect 20898 15376 20904 15388
rect 20956 15376 20962 15428
rect 22557 15419 22615 15425
rect 22557 15416 22569 15419
rect 22204 15388 22569 15416
rect 11517 15351 11575 15357
rect 11517 15348 11529 15351
rect 11348 15320 11529 15348
rect 11517 15317 11529 15320
rect 11563 15317 11575 15351
rect 11517 15311 11575 15317
rect 13538 15308 13544 15360
rect 13596 15308 13602 15360
rect 15565 15351 15623 15357
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 16942 15348 16948 15360
rect 15611 15320 16948 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 19061 15351 19119 15357
rect 19061 15317 19073 15351
rect 19107 15348 19119 15351
rect 19334 15348 19340 15360
rect 19107 15320 19340 15348
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 22204 15357 22232 15388
rect 22557 15385 22569 15388
rect 22603 15385 22615 15419
rect 24486 15416 24492 15428
rect 22557 15379 22615 15385
rect 24044 15388 24492 15416
rect 24044 15357 24072 15388
rect 24486 15376 24492 15388
rect 24544 15416 24550 15428
rect 25240 15425 25268 15524
rect 25332 15524 25636 15552
rect 25332 15493 25360 15524
rect 25682 15512 25688 15564
rect 25740 15512 25746 15564
rect 25774 15512 25780 15564
rect 25832 15512 25838 15564
rect 25884 15552 25912 15592
rect 26053 15555 26111 15561
rect 26053 15552 26065 15555
rect 25884 15524 26065 15552
rect 26053 15521 26065 15524
rect 26099 15521 26111 15555
rect 26053 15515 26111 15521
rect 25317 15487 25375 15493
rect 25317 15453 25329 15487
rect 25363 15453 25375 15487
rect 25317 15447 25375 15453
rect 25498 15444 25504 15496
rect 25556 15444 25562 15496
rect 25593 15487 25651 15493
rect 25593 15453 25605 15487
rect 25639 15484 25651 15487
rect 25700 15484 25728 15512
rect 25639 15456 25728 15484
rect 25792 15484 25820 15512
rect 25869 15487 25927 15493
rect 25869 15484 25881 15487
rect 25792 15456 25881 15484
rect 25639 15453 25651 15456
rect 25593 15447 25651 15453
rect 25225 15419 25283 15425
rect 24544 15388 25084 15416
rect 24544 15376 24550 15388
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 20864 15320 21097 15348
rect 20864 15308 20870 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21085 15311 21143 15317
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15317 22247 15351
rect 22189 15311 22247 15317
rect 24029 15351 24087 15357
rect 24029 15317 24041 15351
rect 24075 15317 24087 15351
rect 24029 15311 24087 15317
rect 24946 15308 24952 15360
rect 25004 15308 25010 15360
rect 25056 15348 25084 15388
rect 25225 15385 25237 15419
rect 25271 15385 25283 15419
rect 25700 15416 25728 15456
rect 25869 15453 25881 15456
rect 25915 15453 25927 15487
rect 25869 15447 25927 15453
rect 25958 15444 25964 15496
rect 26016 15444 26022 15496
rect 26145 15487 26203 15493
rect 26145 15453 26157 15487
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 30193 15487 30251 15493
rect 30193 15453 30205 15487
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 26160 15416 26188 15447
rect 25700 15388 26188 15416
rect 25225 15379 25283 15385
rect 30208 15348 30236 15447
rect 25056 15320 30236 15348
rect 30282 15308 30288 15360
rect 30340 15348 30346 15360
rect 30377 15351 30435 15357
rect 30377 15348 30389 15351
rect 30340 15320 30389 15348
rect 30340 15308 30346 15320
rect 30377 15317 30389 15320
rect 30423 15317 30435 15351
rect 30377 15311 30435 15317
rect 1104 15258 30820 15280
rect 1104 15206 5324 15258
rect 5376 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 12752 15258
rect 12804 15206 12816 15258
rect 12868 15206 12880 15258
rect 12932 15206 12944 15258
rect 12996 15206 13008 15258
rect 13060 15206 20180 15258
rect 20232 15206 20244 15258
rect 20296 15206 20308 15258
rect 20360 15206 20372 15258
rect 20424 15206 20436 15258
rect 20488 15206 27608 15258
rect 27660 15206 27672 15258
rect 27724 15206 27736 15258
rect 27788 15206 27800 15258
rect 27852 15206 27864 15258
rect 27916 15206 30820 15258
rect 1104 15184 30820 15206
rect 5629 15147 5687 15153
rect 5629 15113 5641 15147
rect 5675 15144 5687 15147
rect 5718 15144 5724 15156
rect 5675 15116 5724 15144
rect 5675 15113 5687 15116
rect 5629 15107 5687 15113
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 11701 15147 11759 15153
rect 6236 15116 11008 15144
rect 6236 15104 6242 15116
rect 6362 15076 6368 15088
rect 4816 15048 6368 15076
rect 4816 15017 4844 15048
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 7377 15079 7435 15085
rect 7377 15045 7389 15079
rect 7423 15076 7435 15079
rect 8018 15076 8024 15088
rect 7423 15048 8024 15076
rect 7423 15045 7435 15048
rect 7377 15039 7435 15045
rect 8018 15036 8024 15048
rect 8076 15076 8082 15088
rect 8076 15048 9260 15076
rect 8076 15036 8082 15048
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 15008 4951 15011
rect 5074 15008 5080 15020
rect 4939 14980 5080 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 4890 14832 4896 14884
rect 4948 14872 4954 14884
rect 5077 14875 5135 14881
rect 5077 14872 5089 14875
rect 4948 14844 5089 14872
rect 4948 14832 4954 14844
rect 5077 14841 5089 14844
rect 5123 14841 5135 14875
rect 5077 14835 5135 14841
rect 5184 14816 5212 14971
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5316 14980 5825 15008
rect 5316 14968 5322 14980
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 5813 14971 5871 14977
rect 5994 14968 6000 15020
rect 6052 14968 6058 15020
rect 6089 15011 6147 15017
rect 6089 14977 6101 15011
rect 6135 15008 6147 15011
rect 6270 15008 6276 15020
rect 6135 14980 6276 15008
rect 6135 14977 6147 14980
rect 6089 14971 6147 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 7524 14980 7573 15008
rect 7524 14968 7530 14980
rect 7561 14977 7573 14980
rect 7607 14977 7619 15011
rect 7561 14971 7619 14977
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 8205 15011 8263 15017
rect 7699 14980 8156 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 8128 14952 8156 14980
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8294 15008 8300 15020
rect 8251 14980 8300 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 8389 15011 8447 15017
rect 8389 14977 8401 15011
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 7098 14900 7104 14952
rect 7156 14900 7162 14952
rect 8110 14900 8116 14952
rect 8168 14900 8174 14952
rect 8404 14940 8432 14971
rect 9232 14952 9260 15048
rect 10594 15036 10600 15088
rect 10652 15036 10658 15088
rect 10980 15085 11008 15116
rect 11701 15113 11713 15147
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 10965 15079 11023 15085
rect 10965 15045 10977 15079
rect 11011 15076 11023 15079
rect 11716 15076 11744 15107
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 12124 15116 12265 15144
rect 12124 15104 12130 15116
rect 12253 15113 12265 15116
rect 12299 15113 12311 15147
rect 12253 15107 12311 15113
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 13541 15147 13599 15153
rect 13541 15113 13553 15147
rect 13587 15144 13599 15147
rect 15381 15147 15439 15153
rect 15381 15144 15393 15147
rect 13587 15116 15393 15144
rect 13587 15113 13599 15116
rect 13541 15107 13599 15113
rect 15381 15113 15393 15116
rect 15427 15113 15439 15147
rect 15381 15107 15439 15113
rect 13096 15076 13124 15107
rect 18874 15104 18880 15156
rect 18932 15144 18938 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 18932 15116 19073 15144
rect 18932 15104 18938 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 21453 15147 21511 15153
rect 21453 15113 21465 15147
rect 21499 15144 21511 15147
rect 21542 15144 21548 15156
rect 21499 15116 21548 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 21821 15147 21879 15153
rect 21821 15113 21833 15147
rect 21867 15144 21879 15147
rect 22002 15144 22008 15156
rect 21867 15116 22008 15144
rect 21867 15113 21879 15116
rect 21821 15107 21879 15113
rect 22002 15104 22008 15116
rect 22060 15104 22066 15156
rect 22094 15104 22100 15156
rect 22152 15104 22158 15156
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 22235 15116 24077 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 16301 15079 16359 15085
rect 16301 15076 16313 15079
rect 11011 15048 11744 15076
rect 11011 15045 11023 15048
rect 10965 15039 11023 15045
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 11422 15008 11428 15020
rect 10376 14980 11428 15008
rect 10376 14968 10382 14980
rect 11422 14968 11428 14980
rect 11480 15008 11486 15020
rect 11609 15011 11667 15017
rect 11609 15008 11621 15011
rect 11480 14980 11621 15008
rect 11480 14968 11486 14980
rect 11609 14977 11621 14980
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 8570 14940 8576 14952
rect 8404 14912 8576 14940
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 11716 14940 11744 15048
rect 12452 15048 13124 15076
rect 15028 15048 16313 15076
rect 12452 15017 12480 15048
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 15008 12771 15011
rect 13262 15008 13268 15020
rect 12759 14980 13268 15008
rect 12759 14977 12771 14980
rect 12713 14971 12771 14977
rect 12526 14940 12532 14952
rect 11716 14912 12532 14940
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12728 14940 12756 14971
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13538 15008 13544 15020
rect 13495 14980 13544 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 12676 14912 12756 14940
rect 12676 14900 12682 14912
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 6086 14872 6092 14884
rect 5684 14844 6092 14872
rect 5684 14832 5690 14844
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 7116 14872 7144 14900
rect 7377 14875 7435 14881
rect 7377 14872 7389 14875
rect 7116 14844 7389 14872
rect 7377 14841 7389 14844
rect 7423 14841 7435 14875
rect 13464 14872 13492 14971
rect 13538 14968 13544 14980
rect 13596 15008 13602 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13596 14980 14197 15008
rect 13596 14968 13602 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 14700 14980 14933 15008
rect 14700 14968 14706 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15028 14949 15056 15048
rect 16301 15045 16313 15048
rect 16347 15045 16359 15079
rect 17310 15076 17316 15088
rect 16301 15039 16359 15045
rect 16776 15048 17316 15076
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 14977 15715 15011
rect 15657 14971 15715 14977
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 13556 14912 13645 14940
rect 13556 14884 13584 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14909 15071 14943
rect 15013 14903 15071 14909
rect 7377 14835 7435 14841
rect 7484 14844 13492 14872
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4580 14776 4629 14804
rect 4580 14764 4586 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 5902 14764 5908 14816
rect 5960 14804 5966 14816
rect 7484 14804 7512 14844
rect 13538 14832 13544 14884
rect 13596 14832 13602 14884
rect 14550 14832 14556 14884
rect 14608 14832 14614 14884
rect 15289 14875 15347 14881
rect 15289 14841 15301 14875
rect 15335 14872 15347 14875
rect 15580 14872 15608 14971
rect 15672 14940 15700 14971
rect 15746 14968 15752 15020
rect 15804 14968 15810 15020
rect 15838 14968 15844 15020
rect 15896 14968 15902 15020
rect 15930 14968 15936 15020
rect 15988 14968 15994 15020
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16666 15008 16672 15020
rect 16071 14980 16672 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 15856 14940 15884 14968
rect 16040 14940 16068 14971
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16776 15017 16804 15048
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 19334 15036 19340 15088
rect 19392 15076 19398 15088
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 19392 15048 19441 15076
rect 19392 15036 19398 15048
rect 19429 15045 19441 15048
rect 19475 15045 19487 15079
rect 19429 15039 19487 15045
rect 22112 15076 22140 15104
rect 24049 15076 24077 15116
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 25038 15144 25044 15156
rect 24820 15116 25044 15144
rect 24820 15104 24826 15116
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 24486 15076 24492 15088
rect 22112 15048 22416 15076
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 15672 14912 15884 14940
rect 15948 14912 16068 14940
rect 15335 14844 15608 14872
rect 15335 14841 15347 14844
rect 15289 14835 15347 14841
rect 5960 14776 7512 14804
rect 5960 14764 5966 14776
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 8260 14776 8309 14804
rect 8260 14764 8266 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 9306 14764 9312 14816
rect 9364 14764 9370 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 11204 14776 11253 14804
rect 11204 14764 11210 14776
rect 11241 14773 11253 14776
rect 11287 14804 11299 14807
rect 13630 14804 13636 14816
rect 11287 14776 13636 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 14274 14764 14280 14816
rect 14332 14764 14338 14816
rect 14568 14804 14596 14832
rect 15948 14804 15976 14912
rect 16298 14900 16304 14952
rect 16356 14900 16362 14952
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 17736 14912 18429 14940
rect 17736 14900 17742 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 14568 14776 15976 14804
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 16080 14776 16129 14804
rect 16080 14764 16086 14776
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 16117 14767 16175 14773
rect 16850 14764 16856 14816
rect 16908 14764 16914 14816
rect 18432 14804 18460 14903
rect 18598 14900 18604 14952
rect 18656 14900 18662 14952
rect 18708 14940 18736 14971
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20772 14980 21189 15008
rect 20772 14968 20778 14980
rect 21177 14977 21189 14980
rect 21223 15008 21235 15011
rect 22112 15008 22140 15048
rect 21223 14980 22140 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 18708 14912 20484 14940
rect 20456 14884 20484 14912
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22388 14949 22416 15048
rect 24049 15048 24492 15076
rect 24049 15017 24077 15048
rect 24486 15036 24492 15048
rect 24544 15036 24550 15088
rect 24029 15011 24087 15017
rect 24029 14977 24041 15011
rect 24075 14977 24087 15011
rect 24029 14971 24087 14977
rect 24228 14980 30236 15008
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 22152 14912 22293 14940
rect 22152 14900 22158 14912
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 22373 14943 22431 14949
rect 22373 14909 22385 14943
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 20438 14832 20444 14884
rect 20496 14872 20502 14884
rect 20901 14875 20959 14881
rect 20901 14872 20913 14875
rect 20496 14844 20913 14872
rect 20496 14832 20502 14844
rect 20901 14841 20913 14844
rect 20947 14872 20959 14875
rect 24228 14872 24256 14980
rect 20947 14844 24256 14872
rect 24320 14844 24900 14872
rect 20947 14841 20959 14844
rect 20901 14835 20959 14841
rect 20714 14804 20720 14816
rect 18432 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 21910 14764 21916 14816
rect 21968 14804 21974 14816
rect 22278 14804 22284 14816
rect 21968 14776 22284 14804
rect 21968 14764 21974 14776
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 22738 14764 22744 14816
rect 22796 14804 22802 14816
rect 24320 14813 24348 14844
rect 24872 14816 24900 14844
rect 30208 14816 30236 14980
rect 24305 14807 24363 14813
rect 24305 14804 24317 14807
rect 22796 14776 24317 14804
rect 22796 14764 22802 14776
rect 24305 14773 24317 14776
rect 24351 14773 24363 14807
rect 24305 14767 24363 14773
rect 24489 14807 24547 14813
rect 24489 14773 24501 14807
rect 24535 14804 24547 14807
rect 24762 14804 24768 14816
rect 24535 14776 24768 14804
rect 24535 14773 24547 14776
rect 24489 14767 24547 14773
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 24854 14764 24860 14816
rect 24912 14804 24918 14816
rect 25222 14804 25228 14816
rect 24912 14776 25228 14804
rect 24912 14764 24918 14776
rect 25222 14764 25228 14776
rect 25280 14764 25286 14816
rect 30190 14764 30196 14816
rect 30248 14764 30254 14816
rect 1104 14714 30820 14736
rect 1104 14662 4664 14714
rect 4716 14662 4728 14714
rect 4780 14662 4792 14714
rect 4844 14662 4856 14714
rect 4908 14662 4920 14714
rect 4972 14662 12092 14714
rect 12144 14662 12156 14714
rect 12208 14662 12220 14714
rect 12272 14662 12284 14714
rect 12336 14662 12348 14714
rect 12400 14662 19520 14714
rect 19572 14662 19584 14714
rect 19636 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 26948 14714
rect 27000 14662 27012 14714
rect 27064 14662 27076 14714
rect 27128 14662 27140 14714
rect 27192 14662 27204 14714
rect 27256 14662 30820 14714
rect 1104 14640 30820 14662
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14600 4951 14603
rect 5166 14600 5172 14612
rect 4939 14572 5172 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5902 14560 5908 14612
rect 5960 14560 5966 14612
rect 5997 14603 6055 14609
rect 5997 14569 6009 14603
rect 6043 14600 6055 14603
rect 6086 14600 6092 14612
rect 6043 14572 6092 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6604 14572 6653 14600
rect 6604 14560 6610 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6641 14563 6699 14569
rect 6748 14572 7205 14600
rect 5074 14492 5080 14544
rect 5132 14532 5138 14544
rect 5353 14535 5411 14541
rect 5353 14532 5365 14535
rect 5132 14504 5365 14532
rect 5132 14492 5138 14504
rect 5353 14501 5365 14504
rect 5399 14501 5411 14535
rect 5920 14532 5948 14560
rect 6748 14532 6776 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 13722 14600 13728 14612
rect 11020 14572 13728 14600
rect 11020 14560 11026 14572
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14332 14572 14657 14600
rect 14332 14560 14338 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 16298 14560 16304 14612
rect 16356 14560 16362 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 16632 14572 16773 14600
rect 16632 14560 16638 14572
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 16761 14563 16819 14569
rect 16850 14560 16856 14612
rect 16908 14560 16914 14612
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17957 14603 18015 14609
rect 17957 14600 17969 14603
rect 17000 14572 17969 14600
rect 17000 14560 17006 14572
rect 17957 14569 17969 14572
rect 18003 14569 18015 14603
rect 17957 14563 18015 14569
rect 19150 14560 19156 14612
rect 19208 14600 19214 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 19208 14572 20545 14600
rect 19208 14560 19214 14572
rect 20533 14569 20545 14572
rect 20579 14600 20591 14603
rect 21910 14600 21916 14612
rect 20579 14572 21916 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 22005 14603 22063 14609
rect 22005 14569 22017 14603
rect 22051 14600 22063 14603
rect 22094 14600 22100 14612
rect 22051 14572 22100 14600
rect 22051 14569 22063 14572
rect 22005 14563 22063 14569
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 24486 14560 24492 14612
rect 24544 14600 24550 14612
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 24544 14572 24593 14600
rect 24544 14560 24550 14572
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 24581 14563 24639 14569
rect 25038 14560 25044 14612
rect 25096 14560 25102 14612
rect 25314 14560 25320 14612
rect 25372 14560 25378 14612
rect 25498 14560 25504 14612
rect 25556 14600 25562 14612
rect 26053 14603 26111 14609
rect 26053 14600 26065 14603
rect 25556 14572 26065 14600
rect 25556 14560 25562 14572
rect 26053 14569 26065 14572
rect 26099 14569 26111 14603
rect 26053 14563 26111 14569
rect 5353 14495 5411 14501
rect 5460 14504 5948 14532
rect 6564 14504 6776 14532
rect 7009 14535 7067 14541
rect 5460 14464 5488 14504
rect 2746 14436 5488 14464
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1688 14328 1716 14359
rect 2746 14328 2774 14436
rect 5626 14424 5632 14476
rect 5684 14424 5690 14476
rect 6454 14464 6460 14476
rect 5920 14436 6460 14464
rect 5920 14430 5948 14436
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 3292 14368 4261 14396
rect 3292 14356 3298 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 1688 14300 2774 14328
rect 4264 14328 4292 14359
rect 5534 14356 5540 14408
rect 5592 14356 5598 14408
rect 5718 14356 5724 14408
rect 5776 14356 5782 14408
rect 5828 14405 5948 14430
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6564 14405 6592 14504
rect 7009 14501 7021 14535
rect 7055 14532 7067 14535
rect 7466 14532 7472 14544
rect 7055 14504 7472 14532
rect 7055 14501 7067 14504
rect 7009 14495 7067 14501
rect 7466 14492 7472 14504
rect 7524 14532 7530 14544
rect 7524 14504 7880 14532
rect 7524 14492 7530 14504
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 5813 14402 5948 14405
rect 5813 14399 5871 14402
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 5813 14359 5871 14365
rect 6012 14368 6561 14396
rect 6012 14328 6040 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14365 7159 14399
rect 7576 14396 7604 14427
rect 7852 14405 7880 14504
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7576 14368 7665 14396
rect 7101 14359 7159 14365
rect 7653 14365 7665 14368
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8312 14396 8340 14560
rect 8570 14532 8576 14544
rect 8159 14368 8340 14396
rect 8496 14504 8576 14532
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 4264 14300 6040 14328
rect 6086 14288 6092 14340
rect 6144 14328 6150 14340
rect 6181 14331 6239 14337
rect 6181 14328 6193 14331
rect 6144 14300 6193 14328
rect 6144 14288 6150 14300
rect 6181 14297 6193 14300
rect 6227 14297 6239 14331
rect 6181 14291 6239 14297
rect 934 14220 940 14272
rect 992 14260 998 14272
rect 1489 14263 1547 14269
rect 1489 14260 1501 14263
rect 992 14232 1501 14260
rect 992 14220 998 14232
rect 1489 14229 1501 14232
rect 1535 14229 1547 14263
rect 6196 14260 6224 14291
rect 6270 14288 6276 14340
rect 6328 14328 6334 14340
rect 6365 14331 6423 14337
rect 6365 14328 6377 14331
rect 6328 14300 6377 14328
rect 6328 14288 6334 14300
rect 6365 14297 6377 14300
rect 6411 14297 6423 14331
rect 7116 14328 7144 14359
rect 6365 14291 6423 14297
rect 6564 14300 7144 14328
rect 7745 14331 7803 14337
rect 6564 14272 6592 14300
rect 7745 14297 7757 14331
rect 7791 14328 7803 14331
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 7791 14300 8309 14328
rect 7791 14297 7803 14300
rect 7745 14291 7803 14297
rect 8297 14297 8309 14300
rect 8343 14328 8355 14331
rect 8496 14328 8524 14504
rect 8570 14492 8576 14504
rect 8628 14532 8634 14544
rect 9401 14535 9459 14541
rect 9401 14532 9413 14535
rect 8628 14504 9413 14532
rect 8628 14492 8634 14504
rect 9401 14501 9413 14504
rect 9447 14501 9459 14535
rect 9401 14495 9459 14501
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14464 8815 14467
rect 8803 14436 9076 14464
rect 8803 14433 8815 14436
rect 8757 14427 8815 14433
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8343 14300 8524 14328
rect 8588 14328 8616 14359
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 8956 14328 8984 14356
rect 8588 14300 8984 14328
rect 8343 14297 8355 14300
rect 8297 14291 8355 14297
rect 6546 14260 6552 14272
rect 6196 14232 6552 14260
rect 1489 14223 1547 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14260 7987 14263
rect 8110 14260 8116 14272
rect 7975 14232 8116 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 9048 14269 9076 14436
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9180 14436 9229 14464
rect 9180 14424 9186 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 16022 14464 16028 14476
rect 9217 14427 9275 14433
rect 14384 14436 16028 14464
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 10551 14368 12265 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 12253 14365 12265 14368
rect 12299 14396 12311 14399
rect 12618 14396 12624 14408
rect 12299 14368 12624 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 14384 14405 14412 14436
rect 16022 14424 16028 14436
rect 16080 14424 16086 14476
rect 16316 14464 16344 14560
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 16316 14436 16497 14464
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 16485 14427 16543 14433
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 16868 14464 16896 14560
rect 16623 14436 16896 14464
rect 16960 14504 18276 14532
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 14550 14396 14556 14408
rect 14507 14368 14556 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 14734 14356 14740 14408
rect 14792 14356 14798 14408
rect 16114 14356 16120 14408
rect 16172 14356 16178 14408
rect 16298 14356 16304 14408
rect 16356 14356 16362 14408
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14365 16451 14399
rect 16500 14396 16528 14427
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 16500 14368 16865 14396
rect 16393 14359 16451 14365
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 13464 14328 13492 14356
rect 16408 14328 16436 14359
rect 16960 14328 16988 14504
rect 18248 14464 18276 14504
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 18417 14535 18475 14541
rect 18417 14532 18429 14535
rect 18380 14504 18429 14532
rect 18380 14492 18386 14504
rect 18417 14501 18429 14504
rect 18463 14501 18475 14535
rect 18417 14495 18475 14501
rect 20438 14492 20444 14544
rect 20496 14492 20502 14544
rect 25056 14532 25084 14560
rect 22066 14504 25084 14532
rect 25332 14532 25360 14560
rect 25332 14504 25452 14532
rect 18785 14467 18843 14473
rect 17420 14436 17816 14464
rect 18248 14436 18736 14464
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17129 14399 17187 14405
rect 17129 14365 17141 14399
rect 17175 14365 17187 14399
rect 17129 14359 17187 14365
rect 13464 14300 16988 14328
rect 17052 14272 17080 14359
rect 17144 14328 17172 14359
rect 17310 14356 17316 14408
rect 17368 14356 17374 14408
rect 17420 14405 17448 14436
rect 17788 14405 17816 14436
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 17773 14399 17831 14405
rect 17543 14368 17724 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 17586 14328 17592 14340
rect 17144 14300 17592 14328
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 9033 14263 9091 14269
rect 9033 14229 9045 14263
rect 9079 14260 9091 14263
rect 9214 14260 9220 14272
rect 9079 14232 9220 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 10502 14220 10508 14272
rect 10560 14260 10566 14272
rect 10597 14263 10655 14269
rect 10597 14260 10609 14263
rect 10560 14232 10609 14260
rect 10560 14220 10566 14232
rect 10597 14229 10609 14232
rect 10643 14229 10655 14263
rect 10597 14223 10655 14229
rect 12342 14220 12348 14272
rect 12400 14220 12406 14272
rect 14182 14220 14188 14272
rect 14240 14220 14246 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17696 14260 17724 14368
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 17819 14368 18368 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18340 14269 18368 14368
rect 18708 14328 18736 14436
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 19426 14464 19432 14476
rect 18831 14436 19432 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 19076 14405 19104 14436
rect 19426 14424 19432 14436
rect 19484 14464 19490 14476
rect 20456 14464 20484 14492
rect 19484 14436 20484 14464
rect 19484 14424 19490 14436
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19242 14356 19248 14408
rect 19300 14356 19306 14408
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 21082 14396 21088 14408
rect 20772 14368 21088 14396
rect 20772 14356 20778 14368
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21266 14356 21272 14408
rect 21324 14396 21330 14408
rect 21913 14399 21971 14405
rect 21913 14396 21925 14399
rect 21324 14368 21925 14396
rect 21324 14356 21330 14368
rect 21913 14365 21925 14368
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 19334 14328 19340 14340
rect 18708 14300 19340 14328
rect 19334 14288 19340 14300
rect 19392 14328 19398 14340
rect 20806 14328 20812 14340
rect 19392 14300 20812 14328
rect 19392 14288 19398 14300
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 21361 14331 21419 14337
rect 21361 14297 21373 14331
rect 21407 14328 21419 14331
rect 21450 14328 21456 14340
rect 21407 14300 21456 14328
rect 21407 14297 21419 14300
rect 21361 14291 21419 14297
rect 21450 14288 21456 14300
rect 21508 14288 21514 14340
rect 17092 14232 17724 14260
rect 18325 14263 18383 14269
rect 17092 14220 17098 14232
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 18782 14260 18788 14272
rect 18371 14232 18788 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 18966 14220 18972 14272
rect 19024 14220 19030 14272
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21729 14263 21787 14269
rect 21729 14260 21741 14263
rect 20772 14232 21741 14260
rect 20772 14220 20778 14232
rect 21729 14229 21741 14232
rect 21775 14260 21787 14263
rect 22066 14260 22094 14504
rect 22833 14467 22891 14473
rect 22833 14464 22845 14467
rect 22204 14436 22845 14464
rect 22204 14405 22232 14436
rect 22833 14433 22845 14436
rect 22879 14433 22891 14467
rect 22833 14427 22891 14433
rect 25041 14467 25099 14473
rect 25041 14433 25053 14467
rect 25087 14433 25099 14467
rect 25041 14427 25099 14433
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22370 14356 22376 14408
rect 22428 14356 22434 14408
rect 22646 14356 22652 14408
rect 22704 14356 22710 14408
rect 22738 14356 22744 14408
rect 22796 14356 22802 14408
rect 22922 14356 22928 14408
rect 22980 14356 22986 14408
rect 24854 14356 24860 14408
rect 24912 14356 24918 14408
rect 22278 14288 22284 14340
rect 22336 14288 22342 14340
rect 22511 14331 22569 14337
rect 22511 14297 22523 14331
rect 22557 14328 22569 14331
rect 25056 14328 25084 14427
rect 25222 14424 25228 14476
rect 25280 14464 25286 14476
rect 25317 14467 25375 14473
rect 25317 14464 25329 14467
rect 25280 14436 25329 14464
rect 25280 14424 25286 14436
rect 25317 14433 25329 14436
rect 25363 14433 25375 14467
rect 25317 14427 25375 14433
rect 22557 14300 25084 14328
rect 25332 14328 25360 14427
rect 25424 14405 25452 14504
rect 30374 14492 30380 14544
rect 30432 14492 30438 14544
rect 25409 14399 25467 14405
rect 25409 14365 25421 14399
rect 25455 14365 25467 14399
rect 25409 14359 25467 14365
rect 30190 14356 30196 14408
rect 30248 14356 30254 14408
rect 25685 14331 25743 14337
rect 25685 14328 25697 14331
rect 25332 14300 25697 14328
rect 22557 14297 22569 14300
rect 22511 14291 22569 14297
rect 25685 14297 25697 14300
rect 25731 14297 25743 14331
rect 25685 14291 25743 14297
rect 25866 14288 25872 14340
rect 25924 14288 25930 14340
rect 21775 14232 22094 14260
rect 21775 14229 21787 14232
rect 21729 14223 21787 14229
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 1104 14170 30820 14192
rect 1104 14118 5324 14170
rect 5376 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 12752 14170
rect 12804 14118 12816 14170
rect 12868 14118 12880 14170
rect 12932 14118 12944 14170
rect 12996 14118 13008 14170
rect 13060 14118 20180 14170
rect 20232 14118 20244 14170
rect 20296 14118 20308 14170
rect 20360 14118 20372 14170
rect 20424 14118 20436 14170
rect 20488 14118 27608 14170
rect 27660 14118 27672 14170
rect 27724 14118 27736 14170
rect 27788 14118 27800 14170
rect 27852 14118 27864 14170
rect 27916 14118 30820 14170
rect 1104 14096 30820 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 5166 14056 5172 14068
rect 1627 14028 5172 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 5166 14016 5172 14028
rect 5224 14056 5230 14068
rect 5629 14059 5687 14065
rect 5224 14028 5580 14056
rect 5224 14016 5230 14028
rect 4246 13948 4252 14000
rect 4304 13948 4310 14000
rect 4614 13948 4620 14000
rect 4672 13988 4678 14000
rect 4709 13991 4767 13997
rect 4709 13988 4721 13991
rect 4672 13960 4721 13988
rect 4672 13948 4678 13960
rect 4709 13957 4721 13960
rect 4755 13957 4767 13991
rect 4709 13951 4767 13957
rect 5552 13988 5580 14028
rect 5629 14025 5641 14059
rect 5675 14056 5687 14059
rect 5718 14056 5724 14068
rect 5675 14028 5724 14056
rect 5675 14025 5687 14028
rect 5629 14019 5687 14025
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6178 14016 6184 14068
rect 6236 14016 6242 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 6420 14028 7941 14056
rect 6420 14016 6426 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 8097 14059 8155 14065
rect 8097 14025 8109 14059
rect 8143 14056 8155 14059
rect 8202 14056 8208 14068
rect 8143 14028 8208 14056
rect 8143 14025 8155 14028
rect 8097 14019 8155 14025
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9364 14028 11560 14056
rect 9364 14016 9370 14028
rect 6086 13988 6092 14000
rect 5552 13960 6092 13988
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 5552 13929 5580 13960
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 6196 13988 6224 14016
rect 6454 13988 6460 14000
rect 6196 13960 6460 13988
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 8297 13991 8355 13997
rect 8297 13957 8309 13991
rect 8343 13988 8355 13991
rect 8662 13988 8668 14000
rect 8343 13960 8668 13988
rect 8343 13957 8355 13960
rect 8297 13951 8355 13957
rect 8662 13948 8668 13960
rect 8720 13988 8726 14000
rect 9122 13988 9128 14000
rect 8720 13960 9128 13988
rect 8720 13948 8726 13960
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 6270 13920 6276 13932
rect 5767 13892 6276 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 9508 13929 9536 14028
rect 10502 13948 10508 14000
rect 10560 13948 10566 14000
rect 9493 13923 9551 13929
rect 9493 13889 9505 13923
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 9508 13852 9536 13883
rect 11532 13864 11560 14028
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 14274 14016 14280 14068
rect 14332 14016 14338 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14734 14056 14740 14068
rect 14415 14028 14740 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15746 14056 15752 14068
rect 15059 14028 15752 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 17310 14016 17316 14068
rect 17368 14016 17374 14068
rect 17586 14056 17592 14068
rect 17420 14028 17592 14056
rect 12342 13948 12348 14000
rect 12400 13948 12406 14000
rect 14200 13929 14228 14016
rect 14292 13988 14320 14016
rect 14292 13960 14504 13988
rect 14476 13929 14504 13960
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14752 13920 14780 14016
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14752 13892 14933 13920
rect 14461 13883 14519 13889
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15470 13920 15476 13932
rect 15151 13892 15476 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17328 13920 17356 14016
rect 17420 13997 17448 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18966 14056 18972 14068
rect 17972 14028 18972 14056
rect 17405 13991 17463 13997
rect 17405 13957 17417 13991
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 17175 13892 17356 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17770 13880 17776 13932
rect 17828 13880 17834 13932
rect 17972 13929 18000 14028
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 20349 14059 20407 14065
rect 20349 14025 20361 14059
rect 20395 14056 20407 14059
rect 20530 14056 20536 14068
rect 20395 14028 20536 14056
rect 20395 14025 20407 14028
rect 20349 14019 20407 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 22646 14056 22652 14068
rect 22066 14028 22652 14056
rect 18782 13948 18788 14000
rect 18840 13948 18846 14000
rect 19705 13991 19763 13997
rect 19705 13988 19717 13991
rect 18892 13960 19717 13988
rect 18892 13932 18920 13960
rect 19705 13957 19717 13960
rect 19751 13957 19763 13991
rect 19705 13951 19763 13957
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18230 13920 18236 13932
rect 18095 13892 18236 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18230 13880 18236 13892
rect 18288 13920 18294 13932
rect 18874 13920 18880 13932
rect 18288 13892 18880 13920
rect 18288 13880 18294 13892
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13920 19027 13923
rect 19015 13892 19288 13920
rect 19015 13889 19027 13892
rect 18969 13883 19027 13889
rect 5040 13824 9536 13852
rect 5040 13812 5046 13824
rect 9766 13812 9772 13864
rect 9824 13812 9830 13864
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 14001 13855 14059 13861
rect 14001 13821 14013 13855
rect 14047 13852 14059 13855
rect 16022 13852 16028 13864
rect 14047 13824 16028 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 17313 13855 17371 13861
rect 17313 13821 17325 13855
rect 17359 13852 17371 13855
rect 18782 13852 18788 13864
rect 17359 13824 18788 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 19260 13861 19288 13892
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13821 19303 13855
rect 19720 13852 19748 13951
rect 20806 13948 20812 14000
rect 20864 13988 20870 14000
rect 22066 13988 22094 14028
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 24394 14016 24400 14068
rect 24452 14016 24458 14068
rect 25314 14016 25320 14068
rect 25372 14016 25378 14068
rect 20864 13960 22094 13988
rect 20864 13948 20870 13960
rect 22738 13948 22744 14000
rect 22796 13948 22802 14000
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 22922 13988 22928 14000
rect 22879 13960 22928 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20487 13892 20913 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20901 13889 20913 13892
rect 20947 13920 20959 13923
rect 22094 13920 22100 13932
rect 20947 13892 22100 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 22649 13923 22707 13929
rect 22649 13889 22661 13923
rect 22695 13920 22707 13923
rect 22756 13920 22784 13948
rect 22695 13892 22784 13920
rect 24412 13920 24440 14016
rect 25041 13991 25099 13997
rect 25041 13957 25053 13991
rect 25087 13988 25099 13991
rect 25130 13988 25136 14000
rect 25087 13960 25136 13988
rect 25087 13957 25099 13960
rect 25041 13951 25099 13957
rect 25130 13948 25136 13960
rect 25188 13948 25194 14000
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24412 13892 24593 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 24762 13880 24768 13932
rect 24820 13880 24826 13932
rect 25332 13929 25360 14016
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13889 25375 13923
rect 25317 13883 25375 13889
rect 30469 13923 30527 13929
rect 30469 13889 30481 13923
rect 30515 13889 30527 13923
rect 30469 13883 30527 13889
rect 19720 13824 24440 13852
rect 19245 13815 19303 13821
rect 14660 13756 17172 13784
rect 14660 13728 14688 13756
rect 17144 13728 17172 13756
rect 19426 13744 19432 13796
rect 19484 13744 19490 13796
rect 24412 13784 24440 13824
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24780 13852 24808 13880
rect 25041 13855 25099 13861
rect 25041 13852 25053 13855
rect 24544 13824 25053 13852
rect 24544 13812 24550 13824
rect 25041 13821 25053 13824
rect 25087 13821 25099 13855
rect 30190 13852 30196 13864
rect 25041 13815 25099 13821
rect 25148 13824 30196 13852
rect 25148 13784 25176 13824
rect 30190 13812 30196 13824
rect 30248 13812 30254 13864
rect 30282 13812 30288 13864
rect 30340 13852 30346 13864
rect 30484 13852 30512 13883
rect 30340 13824 30512 13852
rect 30340 13812 30346 13824
rect 24412 13756 25176 13784
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 3234 13716 3240 13728
rect 1728 13688 3240 13716
rect 1728 13676 1734 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 8110 13676 8116 13728
rect 8168 13676 8174 13728
rect 11241 13719 11299 13725
rect 11241 13685 11253 13719
rect 11287 13716 11299 13719
rect 11606 13716 11612 13728
rect 11287 13688 11612 13716
rect 11287 13685 11299 13688
rect 11241 13679 11299 13685
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 13262 13676 13268 13728
rect 13320 13676 13326 13728
rect 14642 13676 14648 13728
rect 14700 13676 14706 13728
rect 16942 13676 16948 13728
rect 17000 13676 17006 13728
rect 17126 13676 17132 13728
rect 17184 13676 17190 13728
rect 19150 13676 19156 13728
rect 19208 13676 19214 13728
rect 20990 13676 20996 13728
rect 21048 13676 21054 13728
rect 22278 13676 22284 13728
rect 22336 13716 22342 13728
rect 22462 13716 22468 13728
rect 22336 13688 22468 13716
rect 22336 13676 22342 13688
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 24673 13719 24731 13725
rect 24673 13685 24685 13719
rect 24719 13716 24731 13719
rect 25222 13716 25228 13728
rect 24719 13688 25228 13716
rect 24719 13685 24731 13688
rect 24673 13679 24731 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 28994 13676 29000 13728
rect 29052 13716 29058 13728
rect 30285 13719 30343 13725
rect 30285 13716 30297 13719
rect 29052 13688 30297 13716
rect 29052 13676 29058 13688
rect 30285 13685 30297 13688
rect 30331 13685 30343 13719
rect 30285 13679 30343 13685
rect 1104 13626 30820 13648
rect 1104 13574 4664 13626
rect 4716 13574 4728 13626
rect 4780 13574 4792 13626
rect 4844 13574 4856 13626
rect 4908 13574 4920 13626
rect 4972 13574 12092 13626
rect 12144 13574 12156 13626
rect 12208 13574 12220 13626
rect 12272 13574 12284 13626
rect 12336 13574 12348 13626
rect 12400 13574 19520 13626
rect 19572 13574 19584 13626
rect 19636 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 26948 13626
rect 27000 13574 27012 13626
rect 27064 13574 27076 13626
rect 27128 13574 27140 13626
rect 27192 13574 27204 13626
rect 27256 13574 30820 13626
rect 1104 13552 30820 13574
rect 4246 13472 4252 13524
rect 4304 13472 4310 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 6270 13512 6276 13524
rect 6227 13484 6276 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 8938 13472 8944 13524
rect 8996 13472 9002 13524
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 10321 13515 10379 13521
rect 10321 13512 10333 13515
rect 9824 13484 10333 13512
rect 9824 13472 9830 13484
rect 10321 13481 10333 13484
rect 10367 13481 10379 13515
rect 10321 13475 10379 13481
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 10744 13484 10824 13512
rect 10744 13472 10750 13484
rect 5184 13416 7880 13444
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 5184 13385 5212 13416
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4120 13348 5181 13376
rect 4120 13336 4126 13348
rect 5169 13345 5181 13348
rect 5215 13345 5227 13379
rect 5169 13339 5227 13345
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 6730 13376 6736 13388
rect 5767 13348 6736 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 7852 13320 7880 13416
rect 9030 13404 9036 13456
rect 9088 13404 9094 13456
rect 10796 13453 10824 13484
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11885 13515 11943 13521
rect 11885 13512 11897 13515
rect 11848 13484 11897 13512
rect 11848 13472 11854 13484
rect 11885 13481 11897 13484
rect 11931 13481 11943 13515
rect 11885 13475 11943 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15528 13484 15577 13512
rect 15528 13472 15534 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 16298 13512 16304 13524
rect 15795 13484 16304 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 10781 13447 10839 13453
rect 10781 13413 10793 13447
rect 10827 13413 10839 13447
rect 15580 13444 15608 13475
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 17313 13515 17371 13521
rect 17313 13512 17325 13515
rect 17184 13484 17325 13512
rect 17184 13472 17190 13484
rect 17313 13481 17325 13484
rect 17359 13481 17371 13515
rect 17313 13475 17371 13481
rect 17420 13484 19104 13512
rect 15841 13447 15899 13453
rect 15841 13444 15853 13447
rect 15580 13416 15853 13444
rect 10781 13407 10839 13413
rect 15841 13413 15853 13416
rect 15887 13413 15899 13447
rect 15841 13407 15899 13413
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 10796 13376 10824 13407
rect 8168 13348 10824 13376
rect 13081 13379 13139 13385
rect 8168 13336 8174 13348
rect 13081 13345 13093 13379
rect 13127 13376 13139 13379
rect 13538 13376 13544 13388
rect 13127 13348 13544 13376
rect 13127 13345 13139 13348
rect 13081 13339 13139 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 17420 13376 17448 13484
rect 19076 13388 19104 13484
rect 23492 13484 30236 13512
rect 21266 13404 21272 13456
rect 21324 13444 21330 13456
rect 21729 13447 21787 13453
rect 21729 13444 21741 13447
rect 21324 13416 21741 13444
rect 21324 13404 21330 13416
rect 21729 13413 21741 13416
rect 21775 13444 21787 13447
rect 23492 13444 23520 13484
rect 21775 13416 23520 13444
rect 21775 13413 21787 13416
rect 21729 13407 21787 13413
rect 15120 13348 17448 13376
rect 17773 13379 17831 13385
rect 15120 13320 15148 13348
rect 1670 13268 1676 13320
rect 1728 13268 1734 13320
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4172 13280 4353 13308
rect 4172 13184 4200 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6144 13280 6469 13308
rect 6144 13268 6150 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 7006 13308 7012 13320
rect 6687 13280 7012 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 7834 13268 7840 13320
rect 7892 13268 7898 13320
rect 10502 13268 10508 13320
rect 10560 13268 10566 13320
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13308 10931 13311
rect 11057 13311 11115 13317
rect 11057 13308 11069 13311
rect 10919 13280 11069 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 11057 13277 11069 13280
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 5994 13200 6000 13252
rect 6052 13200 6058 13252
rect 6213 13243 6271 13249
rect 6213 13209 6225 13243
rect 6259 13240 6271 13243
rect 6549 13243 6607 13249
rect 6549 13240 6561 13243
rect 6259 13212 6561 13240
rect 6259 13209 6271 13212
rect 6213 13203 6271 13209
rect 6549 13209 6561 13212
rect 6595 13209 6607 13243
rect 6549 13203 6607 13209
rect 9398 13200 9404 13252
rect 9456 13200 9462 13252
rect 10612 13240 10640 13271
rect 11606 13268 11612 13320
rect 11664 13268 11670 13320
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 12805 13311 12863 13317
rect 12115 13280 12480 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 10612 13212 11468 13240
rect 11440 13184 11468 13212
rect 934 13132 940 13184
rect 992 13172 998 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 992 13144 1501 13172
rect 992 13132 998 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1489 13135 1547 13141
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 11422 13132 11428 13184
rect 11480 13132 11486 13184
rect 12452 13181 12480 13280
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 13262 13308 13268 13320
rect 12851 13280 13268 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 14829 13311 14887 13317
rect 14829 13308 14841 13311
rect 14792 13280 14841 13308
rect 14792 13268 14798 13280
rect 14829 13277 14841 13280
rect 14875 13277 14887 13311
rect 14829 13271 14887 13277
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15335 13280 16037 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 16025 13277 16037 13280
rect 16071 13308 16083 13311
rect 16114 13308 16120 13320
rect 16071 13280 16120 13308
rect 16071 13277 16083 13280
rect 16025 13271 16083 13277
rect 14568 13240 14596 13268
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 14568 13212 15025 13240
rect 15013 13209 15025 13212
rect 15059 13240 15071 13243
rect 15304 13240 15332 13271
rect 16114 13268 16120 13280
rect 16172 13268 16178 13320
rect 16224 13317 16252 13348
rect 17773 13345 17785 13379
rect 17819 13376 17831 13379
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 17819 13348 18521 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 18509 13345 18521 13348
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 19058 13336 19064 13388
rect 19116 13336 19122 13388
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13376 20039 13379
rect 21910 13376 21916 13388
rect 20027 13348 21916 13376
rect 20027 13345 20039 13348
rect 19981 13339 20039 13345
rect 21910 13336 21916 13348
rect 21968 13336 21974 13388
rect 22370 13336 22376 13388
rect 22428 13336 22434 13388
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13376 22615 13379
rect 22646 13376 22652 13388
rect 22603 13348 22652 13376
rect 22603 13345 22615 13348
rect 22557 13339 22615 13345
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13376 23351 13379
rect 23382 13376 23388 13388
rect 23339 13348 23388 13376
rect 23339 13345 23351 13348
rect 23293 13339 23351 13345
rect 23382 13336 23388 13348
rect 23440 13376 23446 13388
rect 23492 13376 23520 13416
rect 23661 13447 23719 13453
rect 23661 13413 23673 13447
rect 23707 13444 23719 13447
rect 28994 13444 29000 13456
rect 23707 13416 29000 13444
rect 23707 13413 23719 13416
rect 23661 13407 23719 13413
rect 23440 13348 23520 13376
rect 23440 13336 23446 13348
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 17310 13268 17316 13320
rect 17368 13268 17374 13320
rect 17402 13268 17408 13320
rect 17460 13268 17466 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17512 13280 17693 13308
rect 15059 13212 15332 13240
rect 15059 13209 15071 13212
rect 15013 13203 15071 13209
rect 15378 13200 15384 13252
rect 15436 13200 15442 13252
rect 17034 13200 17040 13252
rect 17092 13240 17098 13252
rect 17512 13240 17540 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17681 13271 17739 13277
rect 17788 13280 17877 13308
rect 17788 13252 17816 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 17865 13271 17923 13277
rect 17972 13280 18613 13308
rect 17092 13212 17540 13240
rect 17589 13243 17647 13249
rect 17092 13200 17098 13212
rect 17589 13209 17601 13243
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 12437 13175 12495 13181
rect 12437 13141 12449 13175
rect 12483 13141 12495 13175
rect 12437 13135 12495 13141
rect 12897 13175 12955 13181
rect 12897 13141 12909 13175
rect 12943 13172 12955 13175
rect 13078 13172 13084 13184
rect 12943 13144 13084 13172
rect 12943 13141 12955 13144
rect 12897 13135 12955 13141
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15581 13175 15639 13181
rect 15581 13172 15593 13175
rect 15335 13144 15593 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15581 13141 15593 13144
rect 15627 13141 15639 13175
rect 15581 13135 15639 13141
rect 17126 13132 17132 13184
rect 17184 13132 17190 13184
rect 17604 13172 17632 13203
rect 17770 13200 17776 13252
rect 17828 13200 17834 13252
rect 17972 13172 18000 13280
rect 18601 13277 18613 13280
rect 18647 13308 18659 13311
rect 19150 13308 19156 13320
rect 18647 13280 19156 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 19150 13268 19156 13280
rect 19208 13268 19214 13320
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 22189 13311 22247 13317
rect 22189 13277 22201 13311
rect 22235 13308 22247 13311
rect 22388 13308 22416 13336
rect 22235 13280 22416 13308
rect 22235 13277 22247 13280
rect 22189 13271 22247 13277
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 20257 13243 20315 13249
rect 18196 13212 20208 13240
rect 18196 13200 18202 13212
rect 17604 13144 18000 13172
rect 18966 13132 18972 13184
rect 19024 13132 19030 13184
rect 20180 13172 20208 13212
rect 20257 13209 20269 13243
rect 20303 13240 20315 13243
rect 20530 13240 20536 13252
rect 20303 13212 20536 13240
rect 20303 13209 20315 13212
rect 20257 13203 20315 13209
rect 20530 13200 20536 13212
rect 20588 13200 20594 13252
rect 20990 13200 20996 13252
rect 21048 13200 21054 13252
rect 20622 13172 20628 13184
rect 20180 13144 20628 13172
rect 20622 13132 20628 13144
rect 20680 13132 20686 13184
rect 21818 13132 21824 13184
rect 21876 13172 21882 13184
rect 21913 13175 21971 13181
rect 21913 13172 21925 13175
rect 21876 13144 21925 13172
rect 21876 13132 21882 13144
rect 21913 13141 21925 13144
rect 21959 13141 21971 13175
rect 22112 13172 22140 13271
rect 22738 13268 22744 13320
rect 22796 13308 22802 13320
rect 22833 13311 22891 13317
rect 22833 13308 22845 13311
rect 22796 13280 22845 13308
rect 22796 13268 22802 13280
rect 22833 13277 22845 13280
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23676 13308 23704 13407
rect 28994 13404 29000 13416
rect 29052 13404 29058 13456
rect 23753 13379 23811 13385
rect 23753 13345 23765 13379
rect 23799 13376 23811 13379
rect 23799 13348 24716 13376
rect 23799 13345 23811 13348
rect 23753 13339 23811 13345
rect 24688 13320 24716 13348
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25409 13379 25467 13385
rect 25409 13376 25421 13379
rect 25188 13348 25421 13376
rect 25188 13336 25194 13348
rect 25409 13345 25421 13348
rect 25455 13345 25467 13379
rect 25409 13339 25467 13345
rect 23072 13280 23704 13308
rect 24397 13311 24455 13317
rect 23072 13268 23078 13280
rect 24397 13277 24409 13311
rect 24443 13308 24455 13311
rect 24486 13308 24492 13320
rect 24443 13280 24492 13308
rect 24443 13277 24455 13280
rect 24397 13271 24455 13277
rect 24486 13268 24492 13280
rect 24544 13268 24550 13320
rect 24670 13268 24676 13320
rect 24728 13268 24734 13320
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13308 25559 13311
rect 25866 13308 25872 13320
rect 25547 13280 25872 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 30208 13317 30236 13484
rect 30193 13311 30251 13317
rect 30193 13277 30205 13311
rect 30239 13277 30251 13311
rect 30193 13271 30251 13277
rect 22278 13200 22284 13252
rect 22336 13200 22342 13252
rect 22419 13243 22477 13249
rect 22419 13209 22431 13243
rect 22465 13240 22477 13243
rect 22465 13212 22784 13240
rect 22465 13209 22477 13212
rect 22419 13203 22477 13209
rect 22554 13172 22560 13184
rect 22112 13144 22560 13172
rect 21913 13135 21971 13141
rect 22554 13132 22560 13144
rect 22612 13132 22618 13184
rect 22646 13132 22652 13184
rect 22704 13132 22710 13184
rect 22756 13172 22784 13212
rect 23400 13212 25176 13240
rect 23400 13172 23428 13212
rect 22756 13144 23428 13172
rect 24486 13132 24492 13184
rect 24544 13132 24550 13184
rect 24854 13132 24860 13184
rect 24912 13132 24918 13184
rect 25148 13181 25176 13212
rect 25133 13175 25191 13181
rect 25133 13141 25145 13175
rect 25179 13141 25191 13175
rect 25133 13135 25191 13141
rect 30374 13132 30380 13184
rect 30432 13132 30438 13184
rect 1104 13082 30820 13104
rect 1104 13030 5324 13082
rect 5376 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 12752 13082
rect 12804 13030 12816 13082
rect 12868 13030 12880 13082
rect 12932 13030 12944 13082
rect 12996 13030 13008 13082
rect 13060 13030 20180 13082
rect 20232 13030 20244 13082
rect 20296 13030 20308 13082
rect 20360 13030 20372 13082
rect 20424 13030 20436 13082
rect 20488 13030 27608 13082
rect 27660 13030 27672 13082
rect 27724 13030 27736 13082
rect 27788 13030 27800 13082
rect 27852 13030 27864 13082
rect 27916 13030 30820 13082
rect 1104 13008 30820 13030
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 2746 12940 3249 12968
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2746 12832 2774 12940
rect 3237 12937 3249 12940
rect 3283 12968 3295 12971
rect 4062 12968 4068 12980
rect 3283 12940 4068 12968
rect 3283 12937 3295 12940
rect 3237 12931 3295 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4338 12928 4344 12980
rect 4396 12968 4402 12980
rect 5353 12971 5411 12977
rect 4396 12940 5304 12968
rect 4396 12928 4402 12940
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 4278 12872 5181 12900
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 1719 12804 2774 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5276 12841 5304 12940
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 6086 12968 6092 12980
rect 5399 12940 6092 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6362 12928 6368 12980
rect 6420 12928 6426 12980
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 6788 12940 7788 12968
rect 6788 12928 6794 12940
rect 6380 12900 6408 12928
rect 6380 12872 7420 12900
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5534 12792 5540 12844
rect 5592 12792 5598 12844
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 5810 12832 5816 12844
rect 5767 12804 5816 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 5810 12792 5816 12804
rect 5868 12832 5874 12844
rect 5868 12804 6224 12832
rect 5868 12792 5874 12804
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 6196 12764 6224 12804
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6328 12804 6377 12832
rect 6328 12792 6334 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6512 12804 6837 12832
rect 6512 12792 6518 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7392 12841 7420 12872
rect 7760 12841 7788 12940
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 11480 12940 13277 12968
rect 11480 12928 11486 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 13354 12928 13360 12980
rect 13412 12968 13418 12980
rect 15105 12971 15163 12977
rect 13412 12940 14964 12968
rect 13412 12928 13418 12940
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9033 12903 9091 12909
rect 9033 12900 9045 12903
rect 8352 12872 9045 12900
rect 8352 12860 8358 12872
rect 9033 12869 9045 12872
rect 9079 12900 9091 12903
rect 9398 12900 9404 12912
rect 9079 12872 9404 12900
rect 9079 12869 9091 12872
rect 9033 12863 9091 12869
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 10410 12860 10416 12912
rect 10468 12860 10474 12912
rect 13909 12903 13967 12909
rect 13909 12900 13921 12903
rect 13464 12872 13921 12900
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12801 7159 12835
rect 7101 12795 7159 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 8386 12832 8392 12844
rect 7745 12795 7803 12801
rect 7852 12804 8392 12832
rect 7116 12764 7144 12795
rect 4755 12736 5948 12764
rect 6196 12736 7144 12764
rect 7484 12764 7512 12795
rect 7852 12764 7880 12804
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 8849 12835 8907 12841
rect 8849 12832 8861 12835
rect 8772 12804 8861 12832
rect 7484 12736 7880 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 5920 12696 5948 12736
rect 7926 12724 7932 12776
rect 7984 12764 7990 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7984 12736 8309 12764
rect 7984 12724 7990 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 5920 12668 7205 12696
rect 7193 12665 7205 12668
rect 7239 12665 7251 12699
rect 7193 12659 7251 12665
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 7800 12668 8585 12696
rect 7800 12656 7806 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 6270 12628 6276 12640
rect 6144 12600 6276 12628
rect 6144 12588 6150 12600
rect 6270 12588 6276 12600
rect 6328 12588 6334 12640
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7524 12600 7665 12628
rect 7524 12588 7530 12600
rect 7653 12597 7665 12600
rect 7699 12628 7711 12631
rect 8110 12628 8116 12640
rect 7699 12600 8116 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 8110 12588 8116 12600
rect 8168 12588 8174 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 8772 12637 8800 12804
rect 8849 12801 8861 12804
rect 8895 12801 8907 12835
rect 8849 12795 8907 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11606 12832 11612 12844
rect 11563 12804 11612 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11532 12764 11560 12795
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 13464 12841 13492 12872
rect 13909 12869 13921 12872
rect 13955 12869 13967 12903
rect 14642 12900 14648 12912
rect 13909 12863 13967 12869
rect 14108 12872 14648 12900
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 14108 12841 14136 12872
rect 14642 12860 14648 12872
rect 14700 12900 14706 12912
rect 14700 12872 14780 12900
rect 14700 12860 14706 12872
rect 14752 12841 14780 12872
rect 14936 12844 14964 12940
rect 15105 12937 15117 12971
rect 15151 12968 15163 12971
rect 15930 12968 15936 12980
rect 15151 12940 15936 12968
rect 15151 12937 15163 12940
rect 15105 12931 15163 12937
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16080 12940 17448 12968
rect 16080 12928 16086 12940
rect 16853 12903 16911 12909
rect 16853 12869 16865 12903
rect 16899 12869 16911 12903
rect 16853 12863 16911 12869
rect 14093 12835 14151 12841
rect 13832 12804 14044 12832
rect 11204 12736 11560 12764
rect 11204 12724 11210 12736
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13832 12764 13860 12804
rect 14016 12776 14044 12804
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 14185 12835 14243 12841
rect 14185 12801 14197 12835
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 13688 12736 13860 12764
rect 13688 12724 13694 12736
rect 13906 12724 13912 12776
rect 13964 12724 13970 12776
rect 13998 12724 14004 12776
rect 14056 12724 14062 12776
rect 14200 12764 14228 12795
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15102 12792 15108 12844
rect 15160 12792 15166 12844
rect 14550 12764 14556 12776
rect 14200 12736 14556 12764
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14608 12736 14657 12764
rect 14608 12724 14614 12736
rect 14645 12733 14657 12736
rect 14691 12764 14703 12767
rect 15120 12764 15148 12792
rect 16868 12764 16896 12863
rect 16942 12860 16948 12912
rect 17000 12900 17006 12912
rect 17000 12872 17356 12900
rect 17000 12860 17006 12872
rect 17126 12792 17132 12844
rect 17184 12792 17190 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17328 12841 17356 12872
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12801 17371 12835
rect 17420 12832 17448 12940
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 18785 12971 18843 12977
rect 18785 12968 18797 12971
rect 18656 12940 18797 12968
rect 18656 12928 18662 12940
rect 18785 12937 18797 12940
rect 18831 12937 18843 12971
rect 18785 12931 18843 12937
rect 18966 12928 18972 12980
rect 19024 12928 19030 12980
rect 19426 12928 19432 12980
rect 19484 12928 19490 12980
rect 20530 12928 20536 12980
rect 20588 12928 20594 12980
rect 20901 12971 20959 12977
rect 20901 12937 20913 12971
rect 20947 12937 20959 12971
rect 20901 12931 20959 12937
rect 18984 12900 19012 12928
rect 19271 12903 19329 12909
rect 19271 12900 19283 12903
rect 18984 12872 19283 12900
rect 19271 12869 19283 12872
rect 19317 12869 19329 12903
rect 19271 12863 19329 12869
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17420 12804 17509 12832
rect 17313 12795 17371 12801
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 14691 12736 15148 12764
rect 15212 12736 16896 12764
rect 17144 12764 17172 12792
rect 18064 12764 18092 12792
rect 17144 12736 18092 12764
rect 18984 12764 19012 12795
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 19444 12841 19472 12928
rect 19429 12835 19487 12841
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 20916 12832 20944 12931
rect 21266 12928 21272 12980
rect 21324 12928 21330 12980
rect 21361 12971 21419 12977
rect 21361 12937 21373 12971
rect 21407 12968 21419 12971
rect 21818 12968 21824 12980
rect 21407 12940 21824 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22646 12968 22652 12980
rect 22204 12940 22652 12968
rect 22204 12912 22232 12940
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 23014 12928 23020 12980
rect 23072 12928 23078 12980
rect 23382 12928 23388 12980
rect 23440 12928 23446 12980
rect 23845 12971 23903 12977
rect 23845 12937 23857 12971
rect 23891 12968 23903 12971
rect 24486 12968 24492 12980
rect 23891 12940 24492 12968
rect 23891 12937 23903 12940
rect 23845 12931 23903 12937
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25314 12968 25320 12980
rect 25004 12940 25320 12968
rect 25004 12928 25010 12940
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 30190 12928 30196 12980
rect 30248 12968 30254 12980
rect 30285 12971 30343 12977
rect 30285 12968 30297 12971
rect 30248 12940 30297 12968
rect 30248 12928 30254 12940
rect 30285 12937 30297 12940
rect 30331 12937 30343 12971
rect 30285 12931 30343 12937
rect 22186 12860 22192 12912
rect 22244 12860 22250 12912
rect 22554 12860 22560 12912
rect 22612 12900 22618 12912
rect 22741 12903 22799 12909
rect 22741 12900 22753 12903
rect 22612 12872 22753 12900
rect 22612 12860 22618 12872
rect 22741 12869 22753 12872
rect 22787 12869 22799 12903
rect 22741 12863 22799 12869
rect 20763 12804 20944 12832
rect 22373 12835 22431 12841
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 22373 12801 22385 12835
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 19334 12764 19340 12776
rect 18984 12736 19340 12764
rect 14691 12733 14703 12736
rect 14645 12727 14703 12733
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9180 12668 9674 12696
rect 9180 12656 9186 12668
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8720 12600 8769 12628
rect 8720 12588 8726 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 8757 12591 8815 12597
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9646 12628 9674 12668
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 15212 12696 15240 12736
rect 19334 12724 19340 12736
rect 19392 12724 19398 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 21140 12736 21465 12764
rect 21140 12724 21146 12736
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 22388 12764 22416 12795
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 22649 12835 22707 12841
rect 22649 12832 22661 12835
rect 22520 12804 22661 12832
rect 22520 12792 22526 12804
rect 22649 12801 22661 12804
rect 22695 12801 22707 12835
rect 22649 12795 22707 12801
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12832 22891 12835
rect 23032 12832 23060 12928
rect 23400 12841 23428 12928
rect 22879 12804 23060 12832
rect 22879 12801 22891 12804
rect 22833 12795 22891 12801
rect 22554 12764 22560 12776
rect 22388 12736 22560 12764
rect 21453 12727 21511 12733
rect 22554 12724 22560 12736
rect 22612 12764 22618 12776
rect 22922 12764 22928 12776
rect 22612 12736 22928 12764
rect 22612 12724 22618 12736
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 11020 12668 15240 12696
rect 11020 12656 11026 12668
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 20070 12696 20076 12708
rect 19484 12668 20076 12696
rect 19484 12656 19490 12668
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21174 12696 21180 12708
rect 20864 12668 21180 12696
rect 20864 12656 20870 12668
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 23032 12696 23060 12804
rect 23385 12835 23443 12841
rect 23385 12801 23397 12835
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 24305 12835 24363 12841
rect 24305 12801 24317 12835
rect 24351 12832 24363 12835
rect 24504 12832 24532 12928
rect 24351 12804 24532 12832
rect 24351 12801 24363 12804
rect 24305 12795 24363 12801
rect 24854 12792 24860 12844
rect 24912 12792 24918 12844
rect 25133 12835 25191 12841
rect 25133 12801 25145 12835
rect 25179 12832 25191 12835
rect 25682 12832 25688 12844
rect 25179 12804 25688 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 30282 12792 30288 12844
rect 30340 12832 30346 12844
rect 30377 12835 30435 12841
rect 30377 12832 30389 12835
rect 30340 12804 30389 12832
rect 30340 12792 30346 12804
rect 30377 12801 30389 12804
rect 30423 12801 30435 12835
rect 30377 12795 30435 12801
rect 24670 12724 24676 12776
rect 24728 12724 24734 12776
rect 24765 12767 24823 12773
rect 24765 12733 24777 12767
rect 24811 12764 24823 12767
rect 25866 12764 25872 12776
rect 24811 12736 25872 12764
rect 24811 12733 24823 12736
rect 24765 12727 24823 12733
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 23032 12668 23520 12696
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 9646 12600 10425 12628
rect 10413 12597 10425 12600
rect 10459 12628 10471 12631
rect 11054 12628 11060 12640
rect 10459 12600 11060 12628
rect 10459 12597 10471 12600
rect 10413 12591 10471 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11388 12600 11621 12628
rect 11388 12588 11394 12600
rect 11609 12597 11621 12600
rect 11655 12597 11667 12631
rect 11609 12591 11667 12597
rect 11974 12588 11980 12640
rect 12032 12588 12038 12640
rect 12894 12588 12900 12640
rect 12952 12628 12958 12640
rect 13354 12628 13360 12640
rect 12952 12600 13360 12628
rect 12952 12588 12958 12600
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 16298 12588 16304 12640
rect 16356 12628 16362 12640
rect 18138 12628 18144 12640
rect 16356 12600 18144 12628
rect 16356 12588 16362 12600
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19150 12628 19156 12640
rect 18748 12600 19156 12628
rect 18748 12588 18754 12600
rect 19150 12588 19156 12600
rect 19208 12628 19214 12640
rect 22278 12628 22284 12640
rect 19208 12600 22284 12628
rect 19208 12588 19214 12600
rect 22278 12588 22284 12600
rect 22336 12588 22342 12640
rect 22370 12588 22376 12640
rect 22428 12628 22434 12640
rect 22465 12631 22523 12637
rect 22465 12628 22477 12631
rect 22428 12600 22477 12628
rect 22428 12588 22434 12600
rect 22465 12597 22477 12600
rect 22511 12628 22523 12631
rect 23014 12628 23020 12640
rect 22511 12600 23020 12628
rect 22511 12597 22523 12600
rect 22465 12591 22523 12597
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 23492 12637 23520 12668
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12597 23535 12631
rect 23477 12591 23535 12597
rect 24581 12631 24639 12637
rect 24581 12597 24593 12631
rect 24627 12628 24639 12631
rect 24688 12628 24716 12724
rect 24627 12600 24716 12628
rect 24627 12597 24639 12600
rect 24581 12591 24639 12597
rect 25038 12588 25044 12640
rect 25096 12628 25102 12640
rect 25317 12631 25375 12637
rect 25317 12628 25329 12631
rect 25096 12600 25329 12628
rect 25096 12588 25102 12600
rect 25317 12597 25329 12600
rect 25363 12597 25375 12631
rect 25317 12591 25375 12597
rect 1104 12538 30820 12560
rect 1104 12486 4664 12538
rect 4716 12486 4728 12538
rect 4780 12486 4792 12538
rect 4844 12486 4856 12538
rect 4908 12486 4920 12538
rect 4972 12486 12092 12538
rect 12144 12486 12156 12538
rect 12208 12486 12220 12538
rect 12272 12486 12284 12538
rect 12336 12486 12348 12538
rect 12400 12486 19520 12538
rect 19572 12486 19584 12538
rect 19636 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 26948 12538
rect 27000 12486 27012 12538
rect 27064 12486 27076 12538
rect 27128 12486 27140 12538
rect 27192 12486 27204 12538
rect 27256 12486 30820 12538
rect 1104 12464 30820 12486
rect 6362 12384 6368 12436
rect 6420 12384 6426 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 8205 12427 8263 12433
rect 6696 12396 8156 12424
rect 6696 12384 6702 12396
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 8021 12359 8079 12365
rect 8021 12356 8033 12359
rect 7892 12328 8033 12356
rect 7892 12316 7898 12328
rect 8021 12325 8033 12328
rect 8067 12325 8079 12359
rect 8128 12356 8156 12396
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8294 12424 8300 12436
rect 8251 12396 8300 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 8444 12396 8493 12424
rect 8444 12384 8450 12396
rect 8481 12393 8493 12396
rect 8527 12393 8539 12427
rect 8481 12387 8539 12393
rect 9306 12384 9312 12436
rect 9364 12384 9370 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10505 12427 10563 12433
rect 10505 12424 10517 12427
rect 10100 12396 10517 12424
rect 10100 12384 10106 12396
rect 10505 12393 10517 12396
rect 10551 12393 10563 12427
rect 10505 12387 10563 12393
rect 10689 12427 10747 12433
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 10962 12424 10968 12436
rect 10735 12396 10968 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 8128 12328 8248 12356
rect 8021 12319 8079 12325
rect 8220 12300 8248 12328
rect 10410 12316 10416 12368
rect 10468 12316 10474 12368
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 7006 12288 7012 12300
rect 4028 12260 7012 12288
rect 4028 12248 4034 12260
rect 7006 12248 7012 12260
rect 7064 12288 7070 12300
rect 7742 12288 7748 12300
rect 7064 12260 7748 12288
rect 7064 12248 7070 12260
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9306 12288 9312 12300
rect 8619 12260 9312 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 10704 12288 10732 12387
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11146 12384 11152 12436
rect 11204 12384 11210 12436
rect 12805 12427 12863 12433
rect 12805 12393 12817 12427
rect 12851 12424 12863 12427
rect 13078 12424 13084 12436
rect 12851 12396 13084 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 13538 12384 13544 12436
rect 13596 12384 13602 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 14458 12424 14464 12436
rect 13955 12396 14464 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 14458 12384 14464 12396
rect 14516 12424 14522 12436
rect 14664 12427 14722 12433
rect 14664 12424 14676 12427
rect 14516 12396 14676 12424
rect 14516 12384 14522 12396
rect 14664 12393 14676 12396
rect 14710 12393 14722 12427
rect 14664 12387 14722 12393
rect 16209 12427 16267 12433
rect 16209 12393 16221 12427
rect 16255 12424 16267 12427
rect 16298 12424 16304 12436
rect 16255 12396 16304 12424
rect 16255 12393 16267 12396
rect 16209 12387 16267 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 17034 12384 17040 12436
rect 17092 12384 17098 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17770 12424 17776 12436
rect 17276 12396 17776 12424
rect 17276 12384 17282 12396
rect 17770 12384 17776 12396
rect 17828 12384 17834 12436
rect 17880 12396 20392 12424
rect 14553 12359 14611 12365
rect 14553 12356 14565 12359
rect 9508 12260 10732 12288
rect 10980 12328 13584 12356
rect 5718 12180 5724 12232
rect 5776 12180 5782 12232
rect 5810 12180 5816 12232
rect 5868 12180 5874 12232
rect 5997 12223 6055 12229
rect 5997 12189 6009 12223
rect 6043 12220 6055 12223
rect 6454 12220 6460 12232
rect 6043 12192 6460 12220
rect 6043 12189 6055 12192
rect 5997 12183 6055 12189
rect 5736 12152 5764 12180
rect 6012 12152 6040 12183
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 7616 12192 8309 12220
rect 7616 12180 7622 12192
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 9508 12229 9536 12260
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12189 9551 12223
rect 9493 12183 9551 12189
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 5736 12124 6040 12152
rect 6181 12155 6239 12161
rect 6181 12121 6193 12155
rect 6227 12152 6239 12155
rect 9600 12152 9628 12183
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9732 12192 9781 12220
rect 9732 12180 9738 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9858 12180 9864 12232
rect 9916 12180 9922 12232
rect 9968 12229 9996 12260
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12220 10287 12223
rect 10686 12220 10692 12232
rect 10275 12192 10692 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10045 12155 10103 12161
rect 10045 12152 10057 12155
rect 6227 12124 7696 12152
rect 9600 12124 10057 12152
rect 6227 12121 6239 12124
rect 6181 12115 6239 12121
rect 5997 12087 6055 12093
rect 5997 12053 6009 12087
rect 6043 12084 6055 12087
rect 6381 12087 6439 12093
rect 6381 12084 6393 12087
rect 6043 12056 6393 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6381 12053 6393 12056
rect 6427 12053 6439 12087
rect 6381 12047 6439 12053
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6822 12084 6828 12096
rect 6595 12056 6828 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7668 12084 7696 12124
rect 10045 12121 10057 12124
rect 10091 12152 10103 12155
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10091 12124 10885 12152
rect 10091 12121 10103 12124
rect 10045 12115 10103 12121
rect 10873 12121 10885 12124
rect 10919 12152 10931 12155
rect 10980 12152 11008 12328
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12288 12127 12291
rect 12529 12291 12587 12297
rect 12529 12288 12541 12291
rect 12115 12260 12541 12288
rect 12115 12257 12127 12260
rect 12069 12251 12127 12257
rect 12529 12257 12541 12260
rect 12575 12257 12587 12291
rect 12529 12251 12587 12257
rect 13446 12248 13452 12300
rect 13504 12248 13510 12300
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12220 11115 12223
rect 11330 12220 11336 12232
rect 11103 12192 11336 12220
rect 11103 12189 11115 12192
rect 11057 12183 11115 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11940 12192 11989 12220
rect 11940 12180 11946 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12452 12152 12480 12183
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13081 12223 13139 12229
rect 13081 12189 13093 12223
rect 13127 12222 13139 12223
rect 13127 12220 13308 12222
rect 13127 12194 13492 12220
rect 13127 12189 13139 12194
rect 13280 12192 13492 12194
rect 13081 12183 13139 12189
rect 10919 12124 11008 12152
rect 11992 12124 12480 12152
rect 10919 12121 10931 12124
rect 10873 12115 10931 12121
rect 11992 12096 12020 12124
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13173 12155 13231 12161
rect 13173 12152 13185 12155
rect 12952 12124 13185 12152
rect 12952 12112 12958 12124
rect 13173 12121 13185 12124
rect 13219 12121 13231 12155
rect 13291 12155 13349 12161
rect 13291 12152 13303 12155
rect 13173 12115 13231 12121
rect 13280 12121 13303 12152
rect 13337 12121 13349 12155
rect 13280 12115 13349 12121
rect 10318 12084 10324 12096
rect 7668 12056 10324 12084
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10686 12093 10692 12096
rect 10673 12087 10692 12093
rect 10673 12053 10685 12087
rect 10673 12047 10692 12053
rect 10686 12044 10692 12047
rect 10744 12044 10750 12096
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11606 12084 11612 12096
rect 11563 12056 11612 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11974 12044 11980 12096
rect 12032 12044 12038 12096
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 13280 12084 13308 12115
rect 12391 12056 13308 12084
rect 13464 12084 13492 12192
rect 13556 12152 13584 12328
rect 13648 12328 14565 12356
rect 13648 12232 13676 12328
rect 14553 12325 14565 12328
rect 14599 12325 14611 12359
rect 14553 12319 14611 12325
rect 15841 12359 15899 12365
rect 15841 12325 15853 12359
rect 15887 12356 15899 12359
rect 17589 12359 17647 12365
rect 17589 12356 17601 12359
rect 15887 12328 17601 12356
rect 15887 12325 15899 12328
rect 15841 12319 15899 12325
rect 17589 12325 17601 12328
rect 17635 12325 17647 12359
rect 17589 12319 17647 12325
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 13832 12260 14473 12288
rect 13832 12232 13860 12260
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 17880 12288 17908 12396
rect 18046 12316 18052 12368
rect 18104 12356 18110 12368
rect 20364 12365 20392 12396
rect 20990 12384 20996 12436
rect 21048 12384 21054 12436
rect 25038 12384 25044 12436
rect 25096 12424 25102 12436
rect 25133 12427 25191 12433
rect 25133 12424 25145 12427
rect 25096 12396 25145 12424
rect 25096 12384 25102 12396
rect 25133 12393 25145 12396
rect 25179 12393 25191 12427
rect 25133 12387 25191 12393
rect 20349 12359 20407 12365
rect 18104 12328 19932 12356
rect 18104 12316 18110 12328
rect 14461 12251 14519 12257
rect 14936 12260 17908 12288
rect 13630 12180 13636 12232
rect 13688 12180 13694 12232
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12220 13967 12223
rect 14642 12220 14648 12232
rect 13955 12192 14648 12220
rect 13955 12189 13967 12192
rect 13909 12183 13967 12189
rect 14642 12180 14648 12192
rect 14700 12220 14706 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14700 12192 14841 12220
rect 14700 12180 14706 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14936 12152 14964 12260
rect 18874 12248 18880 12300
rect 18932 12248 18938 12300
rect 19334 12248 19340 12300
rect 19392 12248 19398 12300
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12220 17279 12223
rect 17402 12220 17408 12232
rect 17267 12192 17408 12220
rect 17267 12189 17279 12192
rect 17221 12183 17279 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17497 12223 17555 12229
rect 17497 12189 17509 12223
rect 17543 12220 17555 12223
rect 18892 12220 18920 12248
rect 19904 12229 19932 12328
rect 20349 12325 20361 12359
rect 20395 12325 20407 12359
rect 23753 12359 23811 12365
rect 20349 12319 20407 12325
rect 20456 12328 21128 12356
rect 20257 12291 20315 12297
rect 20257 12257 20269 12291
rect 20303 12288 20315 12291
rect 20456 12288 20484 12328
rect 20303 12260 20484 12288
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 17543 12192 18092 12220
rect 18892 12192 19257 12220
rect 17543 12189 17555 12192
rect 17497 12183 17555 12189
rect 13556 12124 14964 12152
rect 16209 12155 16267 12161
rect 16209 12121 16221 12155
rect 16255 12152 16267 12155
rect 17034 12152 17040 12164
rect 16255 12124 17040 12152
rect 16255 12121 16267 12124
rect 16209 12115 16267 12121
rect 17034 12112 17040 12124
rect 17092 12112 17098 12164
rect 17420 12152 17448 12180
rect 17862 12152 17868 12164
rect 17420 12124 17868 12152
rect 17862 12112 17868 12124
rect 17920 12152 17926 12164
rect 17957 12155 18015 12161
rect 17957 12152 17969 12155
rect 17920 12124 17969 12152
rect 17920 12112 17926 12124
rect 17957 12121 17969 12124
rect 18003 12121 18015 12155
rect 17957 12115 18015 12121
rect 13906 12084 13912 12096
rect 13464 12056 13912 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 13906 12044 13912 12056
rect 13964 12084 13970 12096
rect 14185 12087 14243 12093
rect 14185 12084 14197 12087
rect 13964 12056 14197 12084
rect 13964 12044 13970 12056
rect 14185 12053 14197 12056
rect 14231 12053 14243 12087
rect 14185 12047 14243 12053
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 16356 12056 16405 12084
rect 16356 12044 16362 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17276 12056 17417 12084
rect 17276 12044 17282 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 17757 12087 17815 12093
rect 17757 12053 17769 12087
rect 17803 12084 17815 12087
rect 18064 12084 18092 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19245 12183 19303 12189
rect 19352 12192 19441 12220
rect 19352 12096 19380 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 19889 12183 19947 12189
rect 20456 12192 20545 12220
rect 20456 12164 20484 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 20625 12223 20683 12229
rect 20625 12189 20637 12223
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20073 12155 20131 12161
rect 20073 12152 20085 12155
rect 19904 12124 20085 12152
rect 19904 12096 19932 12124
rect 20073 12121 20085 12124
rect 20119 12121 20131 12155
rect 20073 12115 20131 12121
rect 20438 12112 20444 12164
rect 20496 12112 20502 12164
rect 18506 12084 18512 12096
rect 17803 12056 18512 12084
rect 17803 12053 17815 12056
rect 17757 12047 17815 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19334 12044 19340 12096
rect 19392 12044 19398 12096
rect 19886 12044 19892 12096
rect 19944 12044 19950 12096
rect 20640 12084 20668 12183
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 20911 12217 20969 12223
rect 20911 12183 20923 12217
rect 20957 12214 20969 12217
rect 21100 12214 21128 12328
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 24854 12356 24860 12368
rect 23799 12328 24860 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 23569 12291 23627 12297
rect 23569 12288 23581 12291
rect 21468 12260 23581 12288
rect 20957 12186 21128 12214
rect 20957 12183 20969 12186
rect 20911 12177 20969 12183
rect 21174 12180 21180 12232
rect 21232 12180 21238 12232
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21468 12229 21496 12260
rect 23569 12257 23581 12260
rect 23615 12257 23627 12291
rect 24872 12288 24900 12316
rect 24872 12260 25544 12288
rect 23569 12251 23627 12257
rect 21453 12223 21511 12229
rect 21453 12220 21465 12223
rect 21324 12192 21465 12220
rect 21324 12180 21330 12192
rect 21453 12189 21465 12192
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 22922 12180 22928 12232
rect 22980 12180 22986 12232
rect 25314 12220 25320 12232
rect 23492 12192 25320 12220
rect 21192 12152 21220 12180
rect 22940 12152 22968 12180
rect 21192 12124 22968 12152
rect 21361 12087 21419 12093
rect 21361 12084 21373 12087
rect 20640 12056 21373 12084
rect 21361 12053 21373 12056
rect 21407 12084 21419 12087
rect 23492 12084 23520 12192
rect 25314 12180 25320 12192
rect 25372 12220 25378 12232
rect 25516 12229 25544 12260
rect 25409 12223 25467 12229
rect 25409 12220 25421 12223
rect 25372 12192 25421 12220
rect 25372 12180 25378 12192
rect 25409 12189 25421 12192
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 25501 12223 25559 12229
rect 25501 12189 25513 12223
rect 25547 12189 25559 12223
rect 25501 12183 25559 12189
rect 24026 12112 24032 12164
rect 24084 12112 24090 12164
rect 24946 12112 24952 12164
rect 25004 12112 25010 12164
rect 25165 12155 25223 12161
rect 25165 12121 25177 12155
rect 25211 12152 25223 12155
rect 25211 12124 25452 12152
rect 25211 12121 25223 12124
rect 25165 12115 25223 12121
rect 21407 12056 23520 12084
rect 21407 12053 21419 12056
rect 21361 12047 21419 12053
rect 25314 12044 25320 12096
rect 25372 12044 25378 12096
rect 25424 12093 25452 12124
rect 25682 12112 25688 12164
rect 25740 12112 25746 12164
rect 25409 12087 25467 12093
rect 25409 12053 25421 12087
rect 25455 12053 25467 12087
rect 25409 12047 25467 12053
rect 1104 11994 30820 12016
rect 1104 11942 5324 11994
rect 5376 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 12752 11994
rect 12804 11942 12816 11994
rect 12868 11942 12880 11994
rect 12932 11942 12944 11994
rect 12996 11942 13008 11994
rect 13060 11942 20180 11994
rect 20232 11942 20244 11994
rect 20296 11942 20308 11994
rect 20360 11942 20372 11994
rect 20424 11942 20436 11994
rect 20488 11942 27608 11994
rect 27660 11942 27672 11994
rect 27724 11942 27736 11994
rect 27788 11942 27800 11994
rect 27852 11942 27864 11994
rect 27916 11942 30820 11994
rect 1104 11920 30820 11942
rect 4982 11880 4988 11892
rect 2976 11852 4988 11880
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 2976 11753 3004 11852
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5261 11883 5319 11889
rect 5261 11849 5273 11883
rect 5307 11880 5319 11883
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5307 11852 6377 11880
rect 5307 11849 5319 11852
rect 5261 11843 5319 11849
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 7462 11883 7520 11889
rect 7462 11849 7474 11883
rect 7508 11880 7520 11883
rect 7558 11880 7564 11892
rect 7508 11852 7564 11880
rect 7508 11849 7520 11852
rect 7462 11843 7520 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7653 11883 7711 11889
rect 7653 11849 7665 11883
rect 7699 11880 7711 11883
rect 8386 11880 8392 11892
rect 7699 11852 8392 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 9858 11840 9864 11892
rect 9916 11840 9922 11892
rect 11606 11840 11612 11892
rect 11664 11840 11670 11892
rect 13078 11840 13084 11892
rect 13136 11880 13142 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13136 11852 13461 11880
rect 13136 11840 13142 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 13538 11840 13544 11892
rect 13596 11840 13602 11892
rect 17221 11883 17279 11889
rect 17221 11849 17233 11883
rect 17267 11880 17279 11883
rect 17678 11880 17684 11892
rect 17267 11852 17684 11880
rect 17267 11849 17279 11852
rect 17221 11843 17279 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 17862 11840 17868 11892
rect 17920 11840 17926 11892
rect 18340 11852 19196 11880
rect 4246 11772 4252 11824
rect 4304 11772 4310 11824
rect 7377 11815 7435 11821
rect 7377 11812 7389 11815
rect 6104 11784 7389 11812
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4580 11716 5181 11744
rect 4580 11704 4586 11716
rect 5169 11713 5181 11716
rect 5215 11744 5227 11747
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5215 11716 5641 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 4488 11648 5365 11676
rect 4488 11636 4494 11648
rect 5353 11645 5365 11648
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4396 11580 4813 11608
rect 4396 11568 4402 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 4801 11571 4859 11577
rect 6104 11552 6132 11784
rect 7377 11781 7389 11784
rect 7423 11812 7435 11815
rect 8570 11812 8576 11824
rect 7423 11784 8064 11812
rect 7423 11781 7435 11784
rect 7377 11775 7435 11781
rect 6822 11704 6828 11756
rect 6880 11704 6886 11756
rect 7285 11747 7343 11753
rect 7285 11713 7297 11747
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7561 11747 7619 11753
rect 7561 11713 7573 11747
rect 7607 11744 7619 11747
rect 7742 11744 7748 11756
rect 7607 11716 7748 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 6549 11679 6607 11685
rect 6549 11676 6561 11679
rect 6288 11648 6561 11676
rect 6288 11552 6316 11648
rect 6549 11645 6561 11648
rect 6595 11645 6607 11679
rect 6549 11639 6607 11645
rect 6641 11679 6699 11685
rect 6641 11645 6653 11679
rect 6687 11645 6699 11679
rect 6641 11639 6699 11645
rect 6656 11608 6684 11639
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 7300 11676 7328 11707
rect 7742 11704 7748 11716
rect 7800 11744 7806 11756
rect 8036 11753 8064 11784
rect 8496 11784 8576 11812
rect 8021 11747 8079 11753
rect 7800 11716 7972 11744
rect 7800 11704 7806 11716
rect 7944 11685 7972 11716
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8297 11747 8355 11753
rect 8067 11716 8248 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 7300 11648 7849 11676
rect 7300 11620 7328 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 7975 11648 8064 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 7282 11608 7288 11620
rect 6656 11580 7288 11608
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 3970 11540 3976 11552
rect 1627 11512 3976 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4580 11512 4721 11540
rect 4580 11500 4586 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 4709 11503 4767 11509
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5718 11540 5724 11552
rect 5316 11512 5724 11540
rect 5316 11500 5322 11512
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 6086 11500 6092 11552
rect 6144 11500 6150 11552
rect 6270 11500 6276 11552
rect 6328 11500 6334 11552
rect 8036 11540 8064 11648
rect 8110 11636 8116 11688
rect 8168 11636 8174 11688
rect 8220 11608 8248 11716
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8386 11744 8392 11756
rect 8343 11716 8392 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 8496 11753 8524 11784
rect 8570 11772 8576 11784
rect 8628 11812 8634 11824
rect 9582 11812 9588 11824
rect 8628 11784 9588 11812
rect 8628 11772 8634 11784
rect 9582 11772 9588 11784
rect 9640 11772 9646 11824
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 8849 11747 8907 11753
rect 8849 11713 8861 11747
rect 8895 11713 8907 11747
rect 8849 11707 8907 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10778 11744 10784 11756
rect 10275 11716 10784 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 8754 11676 8760 11688
rect 8619 11648 8760 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 8864 11608 8892 11707
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 11624 11744 11652 11840
rect 11563 11716 11652 11744
rect 11701 11747 11759 11753
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 13449 11747 13507 11753
rect 11747 11716 12020 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11992 11688 12020 11716
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13556 11744 13584 11840
rect 18340 11824 18368 11852
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 18322 11812 18328 11824
rect 14056 11784 18328 11812
rect 14056 11772 14062 11784
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 18506 11772 18512 11824
rect 18564 11812 18570 11824
rect 19168 11812 19196 11852
rect 19242 11840 19248 11892
rect 19300 11840 19306 11892
rect 22646 11880 22652 11892
rect 19720 11852 22652 11880
rect 19720 11812 19748 11852
rect 22646 11840 22652 11852
rect 22704 11880 22710 11892
rect 22704 11852 22876 11880
rect 22704 11840 22710 11852
rect 18564 11784 19104 11812
rect 19168 11784 19748 11812
rect 18564 11772 18570 11784
rect 13633 11747 13691 11753
rect 13633 11744 13645 11747
rect 13556 11716 13645 11744
rect 13449 11707 13507 11713
rect 13633 11713 13645 11716
rect 13679 11713 13691 11747
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 13633 11707 13691 11713
rect 16408 11716 16773 11744
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10686 11676 10692 11688
rect 10183 11648 10692 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 10744 11648 11621 11676
rect 10744 11636 10750 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11974 11636 11980 11688
rect 12032 11636 12038 11688
rect 13464 11676 13492 11707
rect 13464 11648 13584 11676
rect 8220 11580 8892 11608
rect 9214 11568 9220 11620
rect 9272 11568 9278 11620
rect 9232 11540 9260 11568
rect 13556 11552 13584 11648
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 16408 11676 16436 11716
rect 16761 11713 16773 11716
rect 16807 11744 16819 11747
rect 17034 11744 17040 11756
rect 16807 11716 17040 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11744 17371 11747
rect 17359 11716 17448 11744
rect 17359 11713 17371 11716
rect 17313 11707 17371 11713
rect 17420 11676 17448 11716
rect 17678 11704 17684 11756
rect 17736 11744 17742 11756
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17736 11716 17877 11744
rect 17736 11704 17742 11716
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 18414 11744 18420 11756
rect 18187 11716 18420 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 15436 11648 16436 11676
rect 15436 11636 15442 11648
rect 16408 11620 16436 11648
rect 17052 11648 17448 11676
rect 16390 11568 16396 11620
rect 16448 11568 16454 11620
rect 8036 11512 9260 11540
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10045 11543 10103 11549
rect 10045 11540 10057 11543
rect 10008 11512 10057 11540
rect 10008 11500 10014 11512
rect 10045 11509 10057 11512
rect 10091 11509 10103 11543
rect 10045 11503 10103 11509
rect 13538 11500 13544 11552
rect 13596 11500 13602 11552
rect 15933 11543 15991 11549
rect 15933 11509 15945 11543
rect 15979 11540 15991 11543
rect 16482 11540 16488 11552
rect 15979 11512 16488 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 17052 11549 17080 11648
rect 17420 11608 17448 11648
rect 17773 11679 17831 11685
rect 17773 11645 17785 11679
rect 17819 11676 17831 11679
rect 18064 11676 18092 11707
rect 18414 11704 18420 11716
rect 18472 11744 18478 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18472 11716 18613 11744
rect 18472 11704 18478 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18874 11704 18880 11756
rect 18932 11744 18938 11756
rect 19076 11744 19104 11784
rect 19518 11744 19524 11756
rect 18932 11716 19012 11744
rect 19076 11716 19524 11744
rect 18932 11704 18938 11716
rect 17819 11648 18092 11676
rect 18233 11679 18291 11685
rect 17819 11645 17831 11648
rect 17773 11639 17831 11645
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18782 11676 18788 11688
rect 18279 11648 18788 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18248 11608 18276 11639
rect 18782 11636 18788 11648
rect 18840 11636 18846 11688
rect 18984 11685 19012 11716
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 19720 11744 19748 11784
rect 19886 11772 19892 11824
rect 19944 11812 19950 11824
rect 20073 11815 20131 11821
rect 20073 11812 20085 11815
rect 19944 11784 20085 11812
rect 19944 11772 19950 11784
rect 20073 11781 20085 11784
rect 20119 11781 20131 11815
rect 20073 11775 20131 11781
rect 20257 11815 20315 11821
rect 20257 11781 20269 11815
rect 20303 11812 20315 11815
rect 20990 11812 20996 11824
rect 20303 11784 20996 11812
rect 20303 11781 20315 11784
rect 20257 11775 20315 11781
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 19720 11716 19809 11744
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 22848 11753 22876 11852
rect 22922 11840 22928 11892
rect 22980 11880 22986 11892
rect 23575 11883 23633 11889
rect 23575 11880 23587 11883
rect 22980 11852 23587 11880
rect 22980 11840 22986 11852
rect 23575 11849 23587 11852
rect 23621 11849 23633 11883
rect 23575 11843 23633 11849
rect 23845 11883 23903 11889
rect 23845 11849 23857 11883
rect 23891 11880 23903 11883
rect 24026 11880 24032 11892
rect 23891 11852 24032 11880
rect 23891 11849 23903 11852
rect 23845 11843 23903 11849
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 25314 11840 25320 11892
rect 25372 11840 25378 11892
rect 24857 11815 24915 11821
rect 24857 11812 24869 11815
rect 23768 11784 24869 11812
rect 23768 11753 23796 11784
rect 24857 11781 24869 11784
rect 24903 11781 24915 11815
rect 24857 11775 24915 11781
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21692 11716 21833 11744
rect 21692 11704 21698 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 21821 11707 21879 11713
rect 21928 11716 22753 11744
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19613 11679 19671 11685
rect 19613 11676 19625 11679
rect 19116 11648 19625 11676
rect 19116 11636 19122 11648
rect 19613 11645 19625 11648
rect 19659 11645 19671 11679
rect 19613 11639 19671 11645
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11645 19763 11679
rect 19705 11639 19763 11645
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 20070 11676 20076 11688
rect 19935 11648 20076 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 17420 11580 18276 11608
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 19334 11608 19340 11620
rect 18555 11580 19340 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 19334 11568 19340 11580
rect 19392 11608 19398 11620
rect 19720 11608 19748 11639
rect 20070 11636 20076 11648
rect 20128 11676 20134 11688
rect 21928 11676 21956 11716
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 22741 11707 22799 11713
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 23477 11747 23535 11753
rect 23477 11713 23489 11747
rect 23523 11713 23535 11747
rect 23477 11707 23535 11713
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 23753 11747 23811 11753
rect 23753 11713 23765 11747
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 20128 11648 21956 11676
rect 22189 11679 22247 11685
rect 20128 11636 20134 11648
rect 22189 11645 22201 11679
rect 22235 11676 22247 11679
rect 22554 11676 22560 11688
rect 22235 11648 22560 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 22554 11636 22560 11648
rect 22612 11636 22618 11688
rect 22922 11636 22928 11688
rect 22980 11636 22986 11688
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11676 23075 11679
rect 23063 11648 23152 11676
rect 23063 11645 23075 11648
rect 23017 11639 23075 11645
rect 19392 11580 19748 11608
rect 20441 11611 20499 11617
rect 19392 11568 19398 11580
rect 20441 11577 20453 11611
rect 20487 11577 20499 11611
rect 20441 11571 20499 11577
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11509 17095 11543
rect 17037 11503 17095 11509
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 18782 11549 18788 11552
rect 17405 11543 17463 11549
rect 17405 11540 17417 11543
rect 17276 11512 17417 11540
rect 17276 11500 17282 11512
rect 17405 11509 17417 11512
rect 17451 11509 17463 11543
rect 17405 11503 17463 11509
rect 18325 11543 18383 11549
rect 18325 11509 18337 11543
rect 18371 11540 18383 11543
rect 18766 11543 18788 11549
rect 18766 11540 18778 11543
rect 18371 11512 18778 11540
rect 18371 11509 18383 11512
rect 18325 11503 18383 11509
rect 18766 11509 18778 11512
rect 18766 11503 18788 11509
rect 18782 11500 18788 11503
rect 18840 11500 18846 11552
rect 18874 11500 18880 11552
rect 18932 11500 18938 11552
rect 19426 11500 19432 11552
rect 19484 11500 19490 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 20456 11540 20484 11571
rect 20714 11568 20720 11620
rect 20772 11608 20778 11620
rect 22281 11611 22339 11617
rect 22281 11608 22293 11611
rect 20772 11580 22293 11608
rect 20772 11568 20778 11580
rect 22281 11577 22293 11580
rect 22327 11577 22339 11611
rect 22281 11571 22339 11577
rect 23124 11552 23152 11648
rect 23201 11611 23259 11617
rect 23201 11577 23213 11611
rect 23247 11577 23259 11611
rect 23492 11608 23520 11707
rect 23676 11676 23704 11707
rect 23934 11704 23940 11756
rect 23992 11744 23998 11756
rect 24121 11747 24179 11753
rect 24121 11744 24133 11747
rect 23992 11716 24133 11744
rect 23992 11704 23998 11716
rect 24121 11713 24133 11716
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24394 11744 24400 11756
rect 24351 11716 24400 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 24486 11704 24492 11756
rect 24544 11704 24550 11756
rect 24673 11747 24731 11753
rect 24673 11713 24685 11747
rect 24719 11744 24731 11747
rect 24762 11744 24768 11756
rect 24719 11716 24768 11744
rect 24719 11713 24731 11716
rect 24673 11707 24731 11713
rect 24026 11676 24032 11688
rect 23676 11648 24032 11676
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 24213 11679 24271 11685
rect 24213 11645 24225 11679
rect 24259 11676 24271 11679
rect 24688 11676 24716 11707
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 24872 11744 24900 11775
rect 24949 11747 25007 11753
rect 24949 11744 24961 11747
rect 24872 11716 24961 11744
rect 24949 11713 24961 11716
rect 24995 11713 25007 11747
rect 24949 11707 25007 11713
rect 25133 11747 25191 11753
rect 25133 11713 25145 11747
rect 25179 11744 25191 11747
rect 25222 11744 25228 11756
rect 25179 11716 25228 11744
rect 25179 11713 25191 11716
rect 25133 11707 25191 11713
rect 25222 11704 25228 11716
rect 25280 11704 25286 11756
rect 25332 11744 25360 11840
rect 25501 11747 25559 11753
rect 25501 11744 25513 11747
rect 25332 11716 25513 11744
rect 25501 11713 25513 11716
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25593 11747 25651 11753
rect 25593 11713 25605 11747
rect 25639 11744 25651 11747
rect 25869 11747 25927 11753
rect 25639 11716 25820 11744
rect 25639 11713 25651 11716
rect 25593 11707 25651 11713
rect 24259 11648 24716 11676
rect 25041 11679 25099 11685
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 25041 11645 25053 11679
rect 25087 11676 25099 11679
rect 25682 11676 25688 11688
rect 25087 11648 25688 11676
rect 25087 11645 25099 11648
rect 25041 11639 25099 11645
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 23750 11608 23756 11620
rect 23492 11580 23756 11608
rect 23201 11571 23259 11577
rect 22002 11549 22008 11552
rect 19576 11512 20484 11540
rect 21986 11543 22008 11549
rect 19576 11500 19582 11512
rect 21986 11509 21998 11543
rect 21986 11503 22008 11509
rect 22002 11500 22008 11503
rect 22060 11500 22066 11552
rect 22097 11543 22155 11549
rect 22097 11509 22109 11543
rect 22143 11540 22155 11543
rect 22186 11540 22192 11552
rect 22143 11512 22192 11540
rect 22143 11509 22155 11512
rect 22097 11503 22155 11509
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 23106 11500 23112 11552
rect 23164 11500 23170 11552
rect 23216 11540 23244 11571
rect 23750 11568 23756 11580
rect 23808 11568 23814 11620
rect 25792 11608 25820 11716
rect 25869 11713 25881 11747
rect 25915 11744 25927 11747
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 25915 11716 26985 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 30193 11747 30251 11753
rect 30193 11744 30205 11747
rect 27672 11716 30205 11744
rect 27672 11704 27678 11716
rect 30193 11713 30205 11716
rect 30239 11713 30251 11747
rect 30193 11707 30251 11713
rect 26142 11636 26148 11688
rect 26200 11636 26206 11688
rect 24228 11580 24716 11608
rect 24228 11540 24256 11580
rect 23216 11512 24256 11540
rect 24688 11540 24716 11580
rect 25240 11580 25820 11608
rect 25240 11540 25268 11580
rect 24688 11512 25268 11540
rect 25317 11543 25375 11549
rect 25317 11509 25329 11543
rect 25363 11540 25375 11543
rect 25682 11540 25688 11552
rect 25363 11512 25688 11540
rect 25363 11509 25375 11512
rect 25317 11503 25375 11509
rect 25682 11500 25688 11512
rect 25740 11500 25746 11552
rect 25777 11543 25835 11549
rect 25777 11509 25789 11543
rect 25823 11540 25835 11543
rect 26160 11540 26188 11636
rect 30374 11568 30380 11620
rect 30432 11568 30438 11620
rect 25823 11512 26188 11540
rect 25823 11509 25835 11512
rect 25777 11503 25835 11509
rect 1104 11450 30820 11472
rect 1104 11398 4664 11450
rect 4716 11398 4728 11450
rect 4780 11398 4792 11450
rect 4844 11398 4856 11450
rect 4908 11398 4920 11450
rect 4972 11398 12092 11450
rect 12144 11398 12156 11450
rect 12208 11398 12220 11450
rect 12272 11398 12284 11450
rect 12336 11398 12348 11450
rect 12400 11398 19520 11450
rect 19572 11398 19584 11450
rect 19636 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 26948 11450
rect 27000 11398 27012 11450
rect 27064 11398 27076 11450
rect 27128 11398 27140 11450
rect 27192 11398 27204 11450
rect 27256 11398 30820 11450
rect 1104 11376 30820 11398
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3292 11308 3433 11336
rect 3292 11296 3298 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 4246 11336 4252 11348
rect 4203 11308 4252 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4338 11296 4344 11348
rect 4396 11296 4402 11348
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4580 11308 4997 11336
rect 4580 11296 4586 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 6270 11296 6276 11348
rect 6328 11296 6334 11348
rect 7282 11296 7288 11348
rect 7340 11296 7346 11348
rect 8294 11296 8300 11348
rect 8352 11296 8358 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8665 11339 8723 11345
rect 8665 11336 8677 11339
rect 8444 11308 8677 11336
rect 8444 11296 8450 11308
rect 8665 11305 8677 11308
rect 8711 11305 8723 11339
rect 8665 11299 8723 11305
rect 9306 11296 9312 11348
rect 9364 11296 9370 11348
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 13538 11336 13544 11348
rect 13495 11308 13544 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 14277 11339 14335 11345
rect 14277 11305 14289 11339
rect 14323 11336 14335 11339
rect 15378 11336 15384 11348
rect 14323 11308 15384 11336
rect 14323 11305 14335 11308
rect 14277 11299 14335 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 15948 11308 16589 11336
rect 4356 11200 4384 11296
rect 3620 11172 4384 11200
rect 4816 11240 9260 11268
rect 3620 11141 3648 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 1688 11064 1716 11095
rect 4246 11092 4252 11144
rect 4304 11092 4310 11144
rect 4816 11132 4844 11240
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5629 11203 5687 11209
rect 5399 11172 5580 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 4356 11104 4844 11132
rect 4893 11135 4951 11141
rect 4356 11064 4384 11104
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 5258 11132 5264 11144
rect 4939 11104 5264 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 1688 11036 4384 11064
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 4908 11064 4936 11095
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 5552 11141 5580 11172
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 8205 11203 8263 11209
rect 5675 11172 8064 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6086 11132 6092 11144
rect 5767 11104 6092 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6196 11141 6224 11172
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6362 11092 6368 11144
rect 6420 11092 6426 11144
rect 6840 11141 6868 11172
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 6825 11135 6883 11141
rect 6825 11101 6837 11135
rect 6871 11101 6883 11135
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6825 11095 6883 11101
rect 6932 11104 7021 11132
rect 4488 11036 4936 11064
rect 4488 11024 4494 11036
rect 6748 11008 6776 11095
rect 6932 11076 6960 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7098 11092 7104 11144
rect 7156 11092 7162 11144
rect 7742 11092 7748 11144
rect 7800 11132 7806 11144
rect 8036 11141 8064 11172
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 8386 11200 8392 11212
rect 8251 11172 8392 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7800 11104 7849 11132
rect 7800 11092 7806 11104
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11101 8355 11135
rect 9232 11132 9260 11240
rect 9324 11200 9352 11296
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 13814 11268 13820 11280
rect 11388 11240 13820 11268
rect 11388 11228 11394 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 15948 11200 15976 11308
rect 16577 11305 16589 11308
rect 16623 11336 16635 11339
rect 17586 11336 17592 11348
rect 16623 11308 17592 11336
rect 16623 11305 16635 11308
rect 16577 11299 16635 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 18509 11339 18567 11345
rect 18509 11305 18521 11339
rect 18555 11336 18567 11339
rect 19058 11336 19064 11348
rect 18555 11308 19064 11336
rect 18555 11305 18567 11308
rect 18509 11299 18567 11305
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 21634 11296 21640 11348
rect 21692 11296 21698 11348
rect 22557 11339 22615 11345
rect 22557 11305 22569 11339
rect 22603 11336 22615 11339
rect 22922 11336 22928 11348
rect 22603 11308 22928 11336
rect 22603 11305 22615 11308
rect 22557 11299 22615 11305
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 23106 11296 23112 11348
rect 23164 11336 23170 11348
rect 23201 11339 23259 11345
rect 23201 11336 23213 11339
rect 23164 11308 23213 11336
rect 23164 11296 23170 11308
rect 23201 11305 23213 11308
rect 23247 11305 23259 11339
rect 23201 11299 23259 11305
rect 23569 11339 23627 11345
rect 23569 11305 23581 11339
rect 23615 11336 23627 11339
rect 23934 11336 23940 11348
rect 23615 11308 23940 11336
rect 23615 11305 23627 11308
rect 23569 11299 23627 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 24762 11296 24768 11348
rect 24820 11336 24826 11348
rect 27157 11339 27215 11345
rect 27157 11336 27169 11339
rect 24820 11308 27169 11336
rect 24820 11296 24826 11308
rect 27157 11305 27169 11308
rect 27203 11336 27215 11339
rect 27614 11336 27620 11348
rect 27203 11308 27620 11336
rect 27203 11305 27215 11308
rect 27157 11299 27215 11305
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 24581 11271 24639 11277
rect 16040 11240 21864 11268
rect 16040 11209 16068 11240
rect 21836 11212 21864 11240
rect 24581 11237 24593 11271
rect 24627 11268 24639 11271
rect 25222 11268 25228 11280
rect 24627 11240 25228 11268
rect 24627 11237 24639 11240
rect 24581 11231 24639 11237
rect 25222 11228 25228 11240
rect 25280 11268 25286 11280
rect 25406 11268 25412 11280
rect 25280 11240 25412 11268
rect 25280 11228 25286 11240
rect 25406 11228 25412 11240
rect 25464 11228 25470 11280
rect 9324 11172 15976 11200
rect 16025 11203 16083 11209
rect 16025 11169 16037 11203
rect 16071 11169 16083 11203
rect 16025 11163 16083 11169
rect 16482 11160 16488 11212
rect 16540 11160 16546 11212
rect 18601 11203 18659 11209
rect 18340 11172 18552 11200
rect 11146 11132 11152 11144
rect 9232 11104 11152 11132
rect 8297 11095 8355 11101
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 8312 11064 8340 11095
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11440 11104 11529 11132
rect 11440 11076 11468 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 11664 11104 11805 11132
rect 11664 11092 11670 11104
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 13173 11135 13231 11141
rect 13173 11101 13185 11135
rect 13219 11132 13231 11135
rect 13219 11104 13308 11132
rect 13219 11101 13231 11104
rect 13173 11095 13231 11101
rect 9858 11064 9864 11076
rect 6972 11036 8340 11064
rect 8404 11036 9864 11064
rect 6972 11024 6978 11036
rect 1486 10956 1492 11008
rect 1544 10956 1550 11008
rect 6730 10956 6736 11008
rect 6788 10956 6794 11008
rect 8202 10956 8208 11008
rect 8260 10996 8266 11008
rect 8404 10996 8432 11036
rect 9858 11024 9864 11036
rect 9916 11024 9922 11076
rect 11422 11024 11428 11076
rect 11480 11024 11486 11076
rect 12066 11064 12072 11076
rect 11624 11036 12072 11064
rect 8260 10968 8432 10996
rect 8260 10956 8266 10968
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 11624 11005 11652 11036
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 13280 11008 13308 11104
rect 16298 11092 16304 11144
rect 16356 11092 16362 11144
rect 16393 11135 16451 11141
rect 16393 11101 16405 11135
rect 16439 11101 16451 11135
rect 16500 11132 16528 11160
rect 18340 11141 18368 11172
rect 16669 11135 16727 11141
rect 16669 11132 16681 11135
rect 16500 11104 16681 11132
rect 16393 11095 16451 11101
rect 16669 11101 16681 11104
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 15102 11024 15108 11076
rect 15160 11024 15166 11076
rect 15749 11067 15807 11073
rect 15749 11033 15761 11067
rect 15795 11064 15807 11067
rect 16117 11067 16175 11073
rect 16117 11064 16129 11067
rect 15795 11036 16129 11064
rect 15795 11033 15807 11036
rect 15749 11027 15807 11033
rect 16117 11033 16129 11036
rect 16163 11033 16175 11067
rect 16408 11064 16436 11095
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18524 11132 18552 11172
rect 18601 11169 18613 11203
rect 18647 11200 18659 11203
rect 18647 11172 18920 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 18892 11144 18920 11172
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 21818 11160 21824 11212
rect 21876 11200 21882 11212
rect 21876 11172 25268 11200
rect 21876 11160 21882 11172
rect 18782 11132 18788 11144
rect 18524 11104 18788 11132
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18874 11092 18880 11144
rect 18932 11092 18938 11144
rect 19444 11064 19472 11160
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11132 22799 11135
rect 22787 11104 23060 11132
rect 22787 11101 22799 11104
rect 22741 11095 22799 11101
rect 16408 11036 19472 11064
rect 16117 11027 16175 11033
rect 21266 11024 21272 11076
rect 21324 11024 21330 11076
rect 21453 11067 21511 11073
rect 21453 11033 21465 11067
rect 21499 11064 21511 11067
rect 21910 11064 21916 11076
rect 21499 11036 21916 11064
rect 21499 11033 21511 11036
rect 21453 11027 21511 11033
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 22925 11067 22983 11073
rect 22925 11033 22937 11067
rect 22971 11033 22983 11067
rect 23032 11064 23060 11104
rect 23106 11092 23112 11144
rect 23164 11092 23170 11144
rect 23293 11135 23351 11141
rect 23293 11101 23305 11135
rect 23339 11132 23351 11135
rect 23477 11135 23535 11141
rect 23477 11132 23489 11135
rect 23339 11104 23489 11132
rect 23339 11101 23351 11104
rect 23293 11095 23351 11101
rect 23477 11101 23489 11104
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 23492 11064 23520 11095
rect 23934 11092 23940 11144
rect 23992 11132 23998 11144
rect 24486 11132 24492 11144
rect 23992 11104 24492 11132
rect 23992 11092 23998 11104
rect 24486 11092 24492 11104
rect 24544 11092 24550 11144
rect 24673 11135 24731 11141
rect 24673 11101 24685 11135
rect 24719 11132 24731 11135
rect 24762 11132 24768 11144
rect 24719 11104 24768 11132
rect 24719 11101 24731 11104
rect 24673 11095 24731 11101
rect 24762 11092 24768 11104
rect 24820 11092 24826 11144
rect 25240 11132 25268 11172
rect 25682 11160 25688 11212
rect 25740 11160 25746 11212
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 25240 11104 25421 11132
rect 25409 11101 25421 11104
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 30282 11092 30288 11144
rect 30340 11132 30346 11144
rect 30469 11135 30527 11141
rect 30469 11132 30481 11135
rect 30340 11104 30481 11132
rect 30340 11092 30346 11104
rect 30469 11101 30481 11104
rect 30515 11101 30527 11135
rect 30469 11095 30527 11101
rect 23658 11064 23664 11076
rect 23032 11036 23664 11064
rect 22925 11027 22983 11033
rect 11609 10999 11667 11005
rect 11609 10996 11621 10999
rect 11112 10968 11621 10996
rect 11112 10956 11118 10968
rect 11609 10965 11621 10968
rect 11655 10965 11667 10999
rect 11609 10959 11667 10965
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11756 10968 11989 10996
rect 11756 10956 11762 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 13262 10956 13268 11008
rect 13320 10956 13326 11008
rect 13630 10956 13636 11008
rect 13688 10956 13694 11008
rect 22940 10996 22968 11027
rect 23658 11024 23664 11036
rect 23716 11064 23722 11076
rect 23716 11036 26096 11064
rect 23716 11024 23722 11036
rect 23014 10996 23020 11008
rect 22940 10968 23020 10996
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 26068 10996 26096 11036
rect 26234 11024 26240 11076
rect 26292 11024 26298 11076
rect 26988 11036 30328 11064
rect 26988 10996 27016 11036
rect 30300 11005 30328 11036
rect 26068 10968 27016 10996
rect 30285 10999 30343 11005
rect 30285 10965 30297 10999
rect 30331 10965 30343 10999
rect 30285 10959 30343 10965
rect 1104 10906 30820 10928
rect 1104 10854 5324 10906
rect 5376 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 12752 10906
rect 12804 10854 12816 10906
rect 12868 10854 12880 10906
rect 12932 10854 12944 10906
rect 12996 10854 13008 10906
rect 13060 10854 20180 10906
rect 20232 10854 20244 10906
rect 20296 10854 20308 10906
rect 20360 10854 20372 10906
rect 20424 10854 20436 10906
rect 20488 10854 27608 10906
rect 27660 10854 27672 10906
rect 27724 10854 27736 10906
rect 27788 10854 27800 10906
rect 27852 10854 27864 10906
rect 27916 10854 30820 10906
rect 1104 10832 30820 10854
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 6420 10764 6469 10792
rect 6420 10752 6426 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 6914 10792 6920 10804
rect 6871 10764 6920 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 8294 10752 8300 10804
rect 8352 10752 8358 10804
rect 8570 10752 8576 10804
rect 8628 10752 8634 10804
rect 11146 10792 11152 10804
rect 10244 10764 11152 10792
rect 6730 10724 6736 10736
rect 6656 10696 6736 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 4522 10656 4528 10668
rect 1719 10628 4528 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 6656 10665 6684 10696
rect 6730 10684 6736 10696
rect 6788 10724 6794 10736
rect 8312 10724 8340 10752
rect 9401 10727 9459 10733
rect 9401 10724 9413 10727
rect 6788 10696 8340 10724
rect 9048 10696 9413 10724
rect 6788 10684 6794 10696
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6917 10659 6975 10665
rect 6917 10625 6929 10659
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 6932 10588 6960 10619
rect 8202 10616 8208 10668
rect 8260 10616 8266 10668
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 9048 10665 9076 10696
rect 9401 10693 9413 10696
rect 9447 10693 9459 10727
rect 10244 10724 10272 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 15160 10764 15209 10792
rect 15160 10752 15166 10764
rect 15197 10761 15209 10764
rect 15243 10761 15255 10795
rect 15197 10755 15255 10761
rect 18141 10795 18199 10801
rect 18141 10761 18153 10795
rect 18187 10792 18199 10795
rect 18414 10792 18420 10804
rect 18187 10764 18420 10792
rect 18187 10761 18199 10764
rect 18141 10755 18199 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 20057 10795 20115 10801
rect 20057 10761 20069 10795
rect 20103 10792 20115 10795
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20103 10764 20637 10792
rect 20103 10761 20115 10764
rect 20057 10755 20115 10761
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 21177 10795 21235 10801
rect 21177 10761 21189 10795
rect 21223 10792 21235 10795
rect 21469 10795 21527 10801
rect 21469 10792 21481 10795
rect 21223 10764 21481 10792
rect 21223 10761 21235 10764
rect 21177 10755 21235 10761
rect 21469 10761 21481 10764
rect 21515 10761 21527 10795
rect 21469 10755 21527 10761
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22922 10792 22928 10804
rect 22060 10752 22094 10792
rect 9401 10687 9459 10693
rect 9692 10696 10272 10724
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8496 10628 9045 10656
rect 7098 10588 7104 10600
rect 6932 10560 7104 10588
rect 7098 10548 7104 10560
rect 7156 10588 7162 10600
rect 8110 10588 8116 10600
rect 7156 10560 8116 10588
rect 7156 10548 7162 10560
rect 8110 10548 8116 10560
rect 8168 10588 8174 10600
rect 8496 10588 8524 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9692 10665 9720 10696
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9677 10659 9735 10665
rect 9677 10625 9689 10659
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 8168 10560 8524 10588
rect 8168 10548 8174 10560
rect 8938 10548 8944 10600
rect 8996 10548 9002 10600
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9600 10588 9628 10619
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9824 10628 9873 10656
rect 9824 10616 9830 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10656 10011 10659
rect 10134 10656 10140 10668
rect 9999 10628 10140 10656
rect 9999 10625 10011 10628
rect 9953 10619 10011 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10244 10665 10272 10696
rect 10410 10684 10416 10736
rect 10468 10724 10474 10736
rect 10965 10727 11023 10733
rect 10468 10696 10916 10724
rect 10468 10684 10474 10696
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10318 10616 10324 10668
rect 10376 10616 10382 10668
rect 10594 10616 10600 10668
rect 10652 10616 10658 10668
rect 10888 10665 10916 10696
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11422 10724 11428 10736
rect 11011 10696 11428 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11422 10684 11428 10696
rect 11480 10724 11486 10736
rect 13630 10724 13636 10736
rect 11480 10696 13636 10724
rect 11480 10684 11486 10696
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11054 10616 11060 10668
rect 11112 10616 11118 10668
rect 11238 10616 11244 10668
rect 11296 10616 11302 10668
rect 11333 10659 11391 10665
rect 11333 10625 11345 10659
rect 11379 10656 11391 10659
rect 11606 10656 11612 10668
rect 11379 10628 11612 10656
rect 11379 10625 11391 10628
rect 11333 10619 11391 10625
rect 11606 10616 11612 10628
rect 11664 10656 11670 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11664 10628 11713 10656
rect 11664 10616 11670 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 12452 10665 12480 10696
rect 13630 10684 13636 10696
rect 13688 10724 13694 10736
rect 20257 10727 20315 10733
rect 13688 10696 13768 10724
rect 13688 10684 13694 10696
rect 12437 10659 12495 10665
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12483 10628 12517 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13262 10656 13268 10668
rect 13219 10628 13268 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13740 10665 13768 10696
rect 18432 10696 18736 10724
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15746 10656 15752 10668
rect 15344 10628 15752 10656
rect 15344 10616 15350 10628
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 17460 10628 17785 10656
rect 17460 10616 17466 10628
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 17773 10619 17831 10625
rect 17954 10616 17960 10668
rect 18012 10656 18018 10668
rect 18432 10665 18460 10696
rect 18708 10665 18736 10696
rect 20257 10693 20269 10727
rect 20303 10724 20315 10727
rect 20916 10724 20944 10752
rect 21269 10727 21327 10733
rect 21269 10724 21281 10727
rect 20303 10696 21281 10724
rect 20303 10693 20315 10696
rect 20257 10687 20315 10693
rect 21269 10693 21281 10696
rect 21315 10693 21327 10727
rect 21269 10687 21327 10693
rect 21358 10684 21364 10736
rect 21416 10724 21422 10736
rect 22066 10724 22094 10752
rect 22388 10764 22928 10792
rect 21416 10696 22232 10724
rect 21416 10684 21422 10696
rect 18417 10659 18475 10665
rect 18417 10656 18429 10659
rect 18012 10628 18429 10656
rect 18012 10616 18018 10628
rect 18417 10625 18429 10628
rect 18463 10625 18475 10659
rect 18417 10619 18475 10625
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 18693 10619 18751 10625
rect 18877 10659 18935 10665
rect 18877 10625 18889 10659
rect 18923 10656 18935 10659
rect 20625 10659 20683 10665
rect 18923 10628 20116 10656
rect 18923 10625 18935 10628
rect 18877 10619 18935 10625
rect 9600 10560 10732 10588
rect 9217 10551 9275 10557
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 9232 10520 9260 10551
rect 10704 10529 10732 10560
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 18616 10588 18644 10619
rect 18782 10588 18788 10600
rect 13280 10560 14228 10588
rect 18616 10560 18788 10588
rect 6236 10492 9260 10520
rect 10045 10523 10103 10529
rect 6236 10480 6242 10492
rect 10045 10489 10057 10523
rect 10091 10489 10103 10523
rect 10045 10483 10103 10489
rect 10689 10523 10747 10529
rect 10689 10489 10701 10523
rect 10735 10489 10747 10523
rect 11698 10520 11704 10532
rect 10689 10483 10747 10489
rect 11440 10492 11704 10520
rect 934 10412 940 10464
rect 992 10452 998 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 992 10424 1501 10452
rect 992 10412 998 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 1489 10415 1547 10421
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9582 10452 9588 10464
rect 8904 10424 9588 10452
rect 8904 10412 8910 10424
rect 9582 10412 9588 10424
rect 9640 10452 9646 10464
rect 10060 10452 10088 10483
rect 9640 10424 10088 10452
rect 10505 10455 10563 10461
rect 9640 10412 9646 10424
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11440 10452 11468 10492
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 13280 10520 13308 10560
rect 12032 10492 13308 10520
rect 12032 10480 12038 10492
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 13998 10520 14004 10532
rect 13596 10492 14004 10520
rect 13596 10480 13602 10492
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 14200 10529 14228 10560
rect 18782 10548 18788 10560
rect 18840 10588 18846 10600
rect 18892 10588 18920 10619
rect 18840 10560 18920 10588
rect 18840 10548 18846 10560
rect 14185 10523 14243 10529
rect 14185 10489 14197 10523
rect 14231 10489 14243 10523
rect 14185 10483 14243 10489
rect 10551 10424 11468 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 13633 10455 13691 10461
rect 13633 10452 13645 10455
rect 11664 10424 13645 10452
rect 11664 10412 11670 10424
rect 13633 10421 13645 10424
rect 13679 10452 13691 10455
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13679 10424 13829 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 18230 10412 18236 10464
rect 18288 10412 18294 10464
rect 18782 10412 18788 10464
rect 18840 10412 18846 10464
rect 19889 10455 19947 10461
rect 19889 10421 19901 10455
rect 19935 10452 19947 10455
rect 19978 10452 19984 10464
rect 19935 10424 19984 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 20088 10461 20116 10628
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20640 10588 20668 10619
rect 20806 10616 20812 10668
rect 20864 10616 20870 10668
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10656 20959 10659
rect 21726 10656 21732 10668
rect 20947 10628 21732 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 21726 10616 21732 10628
rect 21784 10616 21790 10668
rect 22204 10665 22232 10696
rect 22388 10665 22416 10764
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 26234 10752 26240 10804
rect 26292 10752 26298 10804
rect 30285 10795 30343 10801
rect 30285 10761 30297 10795
rect 30331 10761 30343 10795
rect 30285 10755 30343 10761
rect 22465 10727 22523 10733
rect 22465 10693 22477 10727
rect 22511 10724 22523 10727
rect 23569 10727 23627 10733
rect 22511 10696 22876 10724
rect 22511 10693 22523 10696
rect 22465 10687 22523 10693
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21836 10628 22017 10656
rect 21082 10588 21088 10600
rect 20640 10560 21088 10588
rect 21082 10548 21088 10560
rect 21140 10548 21146 10600
rect 21177 10591 21235 10597
rect 21177 10557 21189 10591
rect 21223 10588 21235 10591
rect 21836 10588 21864 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 21223 10560 21864 10588
rect 22020 10588 22048 10619
rect 22204 10588 22232 10619
rect 22554 10616 22560 10668
rect 22612 10616 22618 10668
rect 22646 10616 22652 10668
rect 22704 10616 22710 10668
rect 22848 10665 22876 10696
rect 23569 10693 23581 10727
rect 23615 10724 23627 10727
rect 23658 10724 23664 10736
rect 23615 10696 23664 10724
rect 23615 10693 23627 10696
rect 23569 10687 23627 10693
rect 23658 10684 23664 10696
rect 23716 10684 23722 10736
rect 23753 10727 23811 10733
rect 23753 10693 23765 10727
rect 23799 10724 23811 10727
rect 24118 10724 24124 10736
rect 23799 10696 24124 10724
rect 23799 10693 23811 10696
rect 23753 10687 23811 10693
rect 24118 10684 24124 10696
rect 24176 10724 24182 10736
rect 30300 10724 30328 10755
rect 24176 10696 30328 10724
rect 24176 10684 24182 10696
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 22925 10659 22983 10665
rect 22925 10625 22937 10659
rect 22971 10625 22983 10659
rect 22925 10619 22983 10625
rect 22940 10588 22968 10619
rect 23014 10616 23020 10668
rect 23072 10616 23078 10668
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 22020 10560 22094 10588
rect 22204 10560 23397 10588
rect 21223 10557 21235 10560
rect 21177 10551 21235 10557
rect 20806 10480 20812 10532
rect 20864 10520 20870 10532
rect 21821 10523 21879 10529
rect 21821 10520 21833 10523
rect 20864 10492 21833 10520
rect 20864 10480 20870 10492
rect 20073 10455 20131 10461
rect 20073 10421 20085 10455
rect 20119 10452 20131 10455
rect 20714 10452 20720 10464
rect 20119 10424 20720 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21358 10452 21364 10464
rect 21039 10424 21364 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21358 10412 21364 10424
rect 21416 10412 21422 10464
rect 21468 10461 21496 10492
rect 21821 10489 21833 10492
rect 21867 10489 21879 10523
rect 21821 10483 21879 10489
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 22066 10520 22094 10560
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 24026 10588 24032 10600
rect 23385 10551 23443 10557
rect 23584 10560 24032 10588
rect 23584 10532 23612 10560
rect 24026 10548 24032 10560
rect 24084 10588 24090 10600
rect 24596 10588 24624 10619
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 26145 10659 26203 10665
rect 26145 10656 26157 10659
rect 24912 10628 26157 10656
rect 24912 10616 24918 10628
rect 26145 10625 26157 10628
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 30469 10659 30527 10665
rect 30469 10625 30481 10659
rect 30515 10656 30527 10659
rect 30926 10656 30932 10668
rect 30515 10628 30932 10656
rect 30515 10625 30527 10628
rect 30469 10619 30527 10625
rect 30926 10616 30932 10628
rect 30984 10616 30990 10668
rect 24084 10560 24624 10588
rect 24084 10548 24090 10560
rect 23293 10523 23351 10529
rect 21968 10492 23152 10520
rect 21968 10480 21974 10492
rect 21453 10455 21511 10461
rect 21453 10421 21465 10455
rect 21499 10421 21511 10455
rect 21453 10415 21511 10421
rect 21634 10412 21640 10464
rect 21692 10412 21698 10464
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21784 10424 22017 10452
rect 21784 10412 21790 10424
rect 22005 10421 22017 10424
rect 22051 10452 22063 10455
rect 23014 10452 23020 10464
rect 22051 10424 23020 10452
rect 22051 10421 22063 10424
rect 22005 10415 22063 10421
rect 23014 10412 23020 10424
rect 23072 10412 23078 10464
rect 23124 10452 23152 10492
rect 23293 10489 23305 10523
rect 23339 10520 23351 10523
rect 23474 10520 23480 10532
rect 23339 10492 23480 10520
rect 23339 10489 23351 10492
rect 23293 10483 23351 10489
rect 23474 10480 23480 10492
rect 23532 10480 23538 10532
rect 23566 10480 23572 10532
rect 23624 10480 23630 10532
rect 23750 10480 23756 10532
rect 23808 10520 23814 10532
rect 24394 10520 24400 10532
rect 23808 10492 24400 10520
rect 23808 10480 23814 10492
rect 24394 10480 24400 10492
rect 24452 10520 24458 10532
rect 24452 10492 24716 10520
rect 24452 10480 24458 10492
rect 23934 10452 23940 10464
rect 23124 10424 23940 10452
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24688 10461 24716 10492
rect 24673 10455 24731 10461
rect 24673 10421 24685 10455
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 25041 10455 25099 10461
rect 25041 10421 25053 10455
rect 25087 10452 25099 10455
rect 25130 10452 25136 10464
rect 25087 10424 25136 10452
rect 25087 10421 25099 10424
rect 25041 10415 25099 10421
rect 25130 10412 25136 10424
rect 25188 10412 25194 10464
rect 1104 10362 30820 10384
rect 1104 10310 4664 10362
rect 4716 10310 4728 10362
rect 4780 10310 4792 10362
rect 4844 10310 4856 10362
rect 4908 10310 4920 10362
rect 4972 10310 12092 10362
rect 12144 10310 12156 10362
rect 12208 10310 12220 10362
rect 12272 10310 12284 10362
rect 12336 10310 12348 10362
rect 12400 10310 19520 10362
rect 19572 10310 19584 10362
rect 19636 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 26948 10362
rect 27000 10310 27012 10362
rect 27064 10310 27076 10362
rect 27128 10310 27140 10362
rect 27192 10310 27204 10362
rect 27256 10310 30820 10362
rect 1104 10288 30820 10310
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 8938 10208 8944 10260
rect 8996 10248 9002 10260
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8996 10220 9413 10248
rect 8996 10208 9002 10220
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 9769 10251 9827 10257
rect 9769 10217 9781 10251
rect 9815 10248 9827 10251
rect 10594 10248 10600 10260
rect 9815 10220 10600 10248
rect 9815 10217 9827 10220
rect 9769 10211 9827 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11572 10220 14136 10248
rect 11572 10208 11578 10220
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 12618 10180 12624 10192
rect 12406 10152 12624 10180
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 5902 10072 5908 10124
rect 5960 10072 5966 10124
rect 5997 10115 6055 10121
rect 5997 10081 6009 10115
rect 6043 10112 6055 10115
rect 6178 10112 6184 10124
rect 6043 10084 6184 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 7834 10112 7840 10124
rect 7791 10084 7840 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 7834 10072 7840 10084
rect 7892 10112 7898 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7892 10084 8125 10112
rect 7892 10072 7898 10084
rect 8113 10081 8125 10084
rect 8159 10112 8171 10115
rect 8220 10112 8248 10140
rect 8159 10084 8248 10112
rect 8389 10115 8447 10121
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 12406 10112 12434 10152
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 14108 10121 14136 10220
rect 18230 10208 18236 10260
rect 18288 10208 18294 10260
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 21542 10248 21548 10260
rect 19392 10220 21548 10248
rect 19392 10208 19398 10220
rect 21542 10208 21548 10220
rect 21600 10248 21606 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21600 10220 21925 10248
rect 21600 10208 21606 10220
rect 21913 10217 21925 10220
rect 21959 10248 21971 10251
rect 23198 10248 23204 10260
rect 21959 10220 23204 10248
rect 21959 10217 21971 10220
rect 21913 10211 21971 10217
rect 23198 10208 23204 10220
rect 23256 10208 23262 10260
rect 23385 10251 23443 10257
rect 23385 10217 23397 10251
rect 23431 10217 23443 10251
rect 23385 10211 23443 10217
rect 17405 10183 17463 10189
rect 17405 10180 17417 10183
rect 17144 10152 17417 10180
rect 8389 10075 8447 10081
rect 9692 10084 12434 10112
rect 14093 10115 14151 10121
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 4893 10047 4951 10053
rect 4893 10044 4905 10047
rect 1719 10016 4905 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 4893 10013 4905 10016
rect 4939 10044 4951 10047
rect 4982 10044 4988 10056
rect 4939 10016 4988 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5828 10044 5856 10072
rect 6638 10044 6644 10056
rect 5828 10016 6644 10044
rect 5721 10007 5779 10013
rect 5736 9976 5764 10007
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 6730 10004 6736 10056
rect 6788 10004 6794 10056
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7147 10016 7880 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 5902 9976 5908 9988
rect 5736 9948 5908 9976
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 6748 9976 6776 10004
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 6748 9948 7389 9976
rect 7377 9945 7389 9948
rect 7423 9945 7435 9979
rect 7377 9939 7435 9945
rect 7558 9936 7564 9988
rect 7616 9936 7622 9988
rect 7852 9976 7880 10016
rect 7926 10004 7932 10056
rect 7984 10004 7990 10056
rect 8018 10004 8024 10056
rect 8076 10004 8082 10056
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 8128 10016 8217 10044
rect 8036 9976 8064 10004
rect 8128 9988 8156 10016
rect 8205 10013 8217 10016
rect 8251 10013 8263 10047
rect 8404 10044 8432 10075
rect 8481 10047 8539 10053
rect 8481 10044 8493 10047
rect 8404 10016 8493 10044
rect 8205 10007 8263 10013
rect 8481 10013 8493 10016
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8662 10004 8668 10056
rect 8720 10004 8726 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9490 10044 9496 10056
rect 9447 10016 9496 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 7852 9948 8064 9976
rect 8110 9936 8116 9988
rect 8168 9936 8174 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9416 9976 9444 10007
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9582 10004 9588 10056
rect 9640 10004 9646 10056
rect 9692 10053 9720 10084
rect 10428 10056 10456 10084
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 9950 10004 9956 10056
rect 10008 10004 10014 10056
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11606 10044 11612 10056
rect 11296 10016 11612 10044
rect 11296 10004 11302 10016
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11900 10053 11928 10084
rect 14093 10081 14105 10115
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11756 10016 11805 10044
rect 11756 10004 11762 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 11974 10004 11980 10056
rect 12032 10004 12038 10056
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 12084 10016 12357 10044
rect 8444 9948 9444 9976
rect 9968 9976 9996 10004
rect 11992 9976 12020 10004
rect 9968 9948 12020 9976
rect 8444 9936 8450 9948
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5224 9880 5457 9908
rect 5224 9868 5230 9880
rect 5445 9877 5457 9880
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 5537 9911 5595 9917
rect 5537 9877 5549 9911
rect 5583 9908 5595 9911
rect 5718 9908 5724 9920
rect 5583 9880 5724 9908
rect 5583 9877 5595 9880
rect 5537 9871 5595 9877
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 7524 9880 8585 9908
rect 7524 9868 7530 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 12084 9908 12112 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 12253 9979 12311 9985
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 12544 9976 12572 10007
rect 15470 10004 15476 10056
rect 15528 10004 15534 10056
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 16298 10004 16304 10056
rect 16356 10004 16362 10056
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 12299 9948 12572 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 14366 9936 14372 9988
rect 14424 9936 14430 9988
rect 16408 9976 16436 10007
rect 16574 10004 16580 10056
rect 16632 10004 16638 10056
rect 17144 10053 17172 10152
rect 17405 10149 17417 10152
rect 17451 10180 17463 10183
rect 18248 10180 18276 10208
rect 17451 10152 18276 10180
rect 17451 10149 17463 10152
rect 17405 10143 17463 10149
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 17267 10084 17632 10112
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10013 17555 10047
rect 17497 10007 17555 10013
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16408 9948 16681 9976
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16868 9976 16896 10007
rect 17221 9979 17279 9985
rect 17221 9976 17233 9979
rect 16868 9948 17233 9976
rect 16669 9939 16727 9945
rect 17221 9945 17233 9948
rect 17267 9945 17279 9979
rect 17221 9939 17279 9945
rect 11848 9880 12112 9908
rect 12437 9911 12495 9917
rect 11848 9868 11854 9880
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12618 9908 12624 9920
rect 12483 9880 12624 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 15838 9868 15844 9920
rect 15896 9868 15902 9920
rect 15930 9868 15936 9920
rect 15988 9868 15994 9920
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9908 17095 9911
rect 17126 9908 17132 9920
rect 17083 9880 17132 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 17126 9868 17132 9880
rect 17184 9908 17190 9920
rect 17402 9908 17408 9920
rect 17184 9880 17408 9908
rect 17184 9868 17190 9880
rect 17402 9868 17408 9880
rect 17460 9908 17466 9920
rect 17512 9908 17540 10007
rect 17604 9976 17632 10084
rect 17972 10044 18000 10152
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 18800 10112 18828 10208
rect 20070 10180 20076 10192
rect 18095 10084 18828 10112
rect 19306 10152 20076 10180
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17972 10016 18153 10044
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10044 18383 10047
rect 19306 10044 19334 10152
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 20162 10140 20168 10192
rect 20220 10140 20226 10192
rect 20622 10140 20628 10192
rect 20680 10180 20686 10192
rect 21450 10180 21456 10192
rect 20680 10152 21456 10180
rect 20680 10140 20686 10152
rect 21450 10140 21456 10152
rect 21508 10180 21514 10192
rect 23400 10180 23428 10211
rect 23566 10208 23572 10260
rect 23624 10208 23630 10260
rect 23661 10251 23719 10257
rect 23661 10217 23673 10251
rect 23707 10248 23719 10251
rect 23750 10248 23756 10260
rect 23707 10220 23756 10248
rect 23707 10217 23719 10220
rect 23661 10211 23719 10217
rect 23750 10208 23756 10220
rect 23808 10208 23814 10260
rect 23934 10208 23940 10260
rect 23992 10248 23998 10260
rect 30285 10251 30343 10257
rect 30285 10248 30297 10251
rect 23992 10220 30297 10248
rect 23992 10208 23998 10220
rect 30285 10217 30297 10220
rect 30331 10217 30343 10251
rect 30285 10211 30343 10217
rect 23845 10183 23903 10189
rect 23845 10180 23857 10183
rect 21508 10152 22029 10180
rect 23400 10152 23857 10180
rect 21508 10140 21514 10152
rect 19794 10072 19800 10124
rect 19852 10072 19858 10124
rect 18371 10016 19334 10044
rect 18371 10013 18383 10016
rect 18325 10007 18383 10013
rect 19702 10004 19708 10056
rect 19760 10004 19766 10056
rect 20088 10053 20116 10140
rect 20180 10112 20208 10140
rect 20349 10115 20407 10121
rect 20349 10112 20361 10115
rect 20180 10084 20361 10112
rect 20349 10081 20361 10084
rect 20395 10081 20407 10115
rect 20349 10075 20407 10081
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 22001 10112 22029 10152
rect 23845 10149 23857 10152
rect 23891 10180 23903 10183
rect 24946 10180 24952 10192
rect 23891 10152 24952 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 25501 10183 25559 10189
rect 25501 10180 25513 10183
rect 25056 10152 25513 10180
rect 24489 10115 24547 10121
rect 24489 10112 24501 10115
rect 20579 10084 21588 10112
rect 22001 10084 24501 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 17604 9948 18184 9976
rect 18156 9920 18184 9948
rect 17460 9880 17540 9908
rect 17460 9868 17466 9880
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17736 9880 17877 9908
rect 17736 9868 17742 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 18138 9868 18144 9920
rect 18196 9868 18202 9920
rect 19904 9908 19932 10007
rect 20180 9976 20208 10007
rect 20254 10004 20260 10056
rect 20312 10044 20318 10056
rect 20625 10047 20683 10053
rect 20625 10044 20637 10047
rect 20312 10016 20637 10044
rect 20312 10004 20318 10016
rect 20625 10013 20637 10016
rect 20671 10013 20683 10047
rect 20625 10007 20683 10013
rect 20809 10047 20867 10053
rect 20809 10013 20821 10047
rect 20855 10044 20867 10047
rect 20898 10044 20904 10056
rect 20855 10016 20904 10044
rect 20855 10013 20867 10016
rect 20809 10007 20867 10013
rect 20438 9976 20444 9988
rect 20180 9948 20444 9976
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 20530 9936 20536 9988
rect 20588 9976 20594 9988
rect 20824 9976 20852 10007
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 20588 9948 20852 9976
rect 20588 9936 20594 9948
rect 20548 9908 20576 9936
rect 21008 9920 21036 10007
rect 21560 9976 21588 10084
rect 24489 10081 24501 10084
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 24673 10115 24731 10121
rect 24673 10081 24685 10115
rect 24719 10112 24731 10115
rect 24857 10115 24915 10121
rect 24857 10112 24869 10115
rect 24719 10084 24869 10112
rect 24719 10081 24731 10084
rect 24673 10075 24731 10081
rect 24857 10081 24869 10084
rect 24903 10081 24915 10115
rect 25056 10112 25084 10152
rect 25501 10149 25513 10152
rect 25547 10149 25559 10183
rect 25501 10143 25559 10149
rect 24857 10075 24915 10081
rect 24964 10084 25084 10112
rect 21634 10004 21640 10056
rect 21692 10004 21698 10056
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 22005 10047 22063 10053
rect 22005 10013 22017 10047
rect 22051 10044 22063 10047
rect 22370 10044 22376 10056
rect 22051 10016 22376 10044
rect 22051 10013 22063 10016
rect 22005 10007 22063 10013
rect 21744 9976 21772 10007
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 23109 10047 23167 10053
rect 23109 10044 23121 10047
rect 22612 10016 23121 10044
rect 22612 10004 22618 10016
rect 23109 10013 23121 10016
rect 23155 10044 23167 10047
rect 24118 10044 24124 10056
rect 23155 10016 24124 10044
rect 23155 10013 23167 10016
rect 23109 10007 23167 10013
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10044 24823 10047
rect 24964 10044 24992 10084
rect 25314 10072 25320 10124
rect 25372 10072 25378 10124
rect 24811 10016 24992 10044
rect 24811 10013 24823 10016
rect 24765 10007 24823 10013
rect 25038 10004 25044 10056
rect 25096 10004 25102 10056
rect 25130 10004 25136 10056
rect 25188 10004 25194 10056
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10044 25283 10047
rect 25406 10044 25412 10056
rect 25271 10016 25412 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 25406 10004 25412 10016
rect 25464 10044 25470 10056
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 25464 10016 25697 10044
rect 25464 10004 25470 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10013 25835 10047
rect 25777 10007 25835 10013
rect 21560 9948 21772 9976
rect 23198 9936 23204 9988
rect 23256 9976 23262 9988
rect 23750 9976 23756 9988
rect 23256 9948 23756 9976
rect 23256 9936 23262 9948
rect 23750 9936 23756 9948
rect 23808 9936 23814 9988
rect 19904 9880 20576 9908
rect 20990 9868 20996 9920
rect 21048 9868 21054 9920
rect 21453 9911 21511 9917
rect 21453 9877 21465 9911
rect 21499 9908 21511 9911
rect 22094 9908 22100 9920
rect 21499 9880 22100 9908
rect 21499 9877 21511 9880
rect 21453 9871 21511 9877
rect 22094 9868 22100 9880
rect 22152 9868 22158 9920
rect 24486 9868 24492 9920
rect 24544 9868 24550 9920
rect 25056 9908 25084 10004
rect 25148 9976 25176 10004
rect 25501 9979 25559 9985
rect 25501 9976 25513 9979
rect 25148 9948 25513 9976
rect 25501 9945 25513 9948
rect 25547 9945 25559 9979
rect 25792 9976 25820 10007
rect 30282 10004 30288 10056
rect 30340 10044 30346 10056
rect 30469 10047 30527 10053
rect 30469 10044 30481 10047
rect 30340 10016 30481 10044
rect 30340 10004 30346 10016
rect 30469 10013 30481 10016
rect 30515 10013 30527 10047
rect 30469 10007 30527 10013
rect 25501 9939 25559 9945
rect 25608 9948 25820 9976
rect 25608 9908 25636 9948
rect 25056 9880 25636 9908
rect 1104 9818 30820 9840
rect 1104 9766 5324 9818
rect 5376 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 12752 9818
rect 12804 9766 12816 9818
rect 12868 9766 12880 9818
rect 12932 9766 12944 9818
rect 12996 9766 13008 9818
rect 13060 9766 20180 9818
rect 20232 9766 20244 9818
rect 20296 9766 20308 9818
rect 20360 9766 20372 9818
rect 20424 9766 20436 9818
rect 20488 9766 27608 9818
rect 27660 9766 27672 9818
rect 27724 9766 27736 9818
rect 27788 9766 27800 9818
rect 27852 9766 27864 9818
rect 27916 9766 30820 9818
rect 1104 9744 30820 9766
rect 5166 9664 5172 9716
rect 5224 9664 5230 9716
rect 6730 9664 6736 9716
rect 6788 9664 6794 9716
rect 7193 9707 7251 9713
rect 7193 9673 7205 9707
rect 7239 9704 7251 9707
rect 7558 9704 7564 9716
rect 7239 9676 7564 9704
rect 7239 9673 7251 9676
rect 7193 9667 7251 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 8110 9704 8116 9716
rect 7668 9676 8116 9704
rect 4522 9596 4528 9648
rect 4580 9596 4586 9648
rect 5184 9636 5212 9664
rect 7668 9636 7696 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 10594 9664 10600 9716
rect 10652 9664 10658 9716
rect 11146 9664 11152 9716
rect 11204 9664 11210 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 15028 9676 15301 9704
rect 5184 9608 5488 9636
rect 5460 9577 5488 9608
rect 5828 9608 7512 9636
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 5828 9577 5856 9608
rect 7484 9580 7512 9608
rect 7576 9608 7696 9636
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9537 5871 9571
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 5813 9531 5871 9537
rect 6104 9540 6561 9568
rect 6104 9512 6132 9540
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 6914 9568 6920 9580
rect 6595 9540 6920 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4982 9500 4988 9512
rect 3651 9472 4988 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5123 9472 5304 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5276 9432 5304 9472
rect 5350 9460 5356 9512
rect 5408 9460 5414 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5552 9472 6009 9500
rect 5552 9432 5580 9472
rect 5997 9469 6009 9472
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6086 9460 6092 9512
rect 6144 9460 6150 9512
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 6454 9460 6460 9512
rect 6512 9460 6518 9512
rect 5276 9404 5580 9432
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 6472 9432 6500 9460
rect 5684 9404 6500 9432
rect 6748 9432 6776 9540
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7107 9574 7165 9577
rect 7024 9571 7165 9574
rect 7024 9546 7119 9571
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7024 9500 7052 9546
rect 7107 9537 7119 9546
rect 7153 9537 7165 9571
rect 7107 9531 7165 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 6880 9472 7052 9500
rect 6880 9460 6886 9472
rect 7300 9432 7328 9531
rect 7466 9528 7472 9580
rect 7524 9528 7530 9580
rect 7576 9577 7604 9608
rect 7834 9596 7840 9648
rect 7892 9596 7898 9648
rect 11606 9636 11612 9648
rect 10980 9608 11612 9636
rect 7561 9571 7619 9577
rect 7561 9537 7573 9571
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 8018 9568 8024 9580
rect 7699 9540 8024 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 8018 9528 8024 9540
rect 8076 9568 8082 9580
rect 8294 9568 8300 9580
rect 8076 9540 8300 9568
rect 8076 9528 8082 9540
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 10980 9577 11008 9608
rect 11606 9596 11612 9608
rect 11664 9636 11670 9648
rect 11882 9636 11888 9648
rect 11664 9608 11888 9636
rect 11664 9596 11670 9608
rect 11882 9596 11888 9608
rect 11940 9636 11946 9648
rect 12621 9639 12679 9645
rect 12621 9636 12633 9639
rect 11940 9608 12633 9636
rect 11940 9596 11946 9608
rect 12621 9605 12633 9608
rect 12667 9605 12679 9639
rect 12621 9599 12679 9605
rect 12894 9596 12900 9648
rect 12952 9636 12958 9648
rect 13354 9636 13360 9648
rect 12952 9608 13360 9636
rect 12952 9596 12958 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 14921 9639 14979 9645
rect 14921 9605 14933 9639
rect 14967 9636 14979 9639
rect 15028 9636 15056 9676
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 15335 9676 16068 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 14967 9608 15056 9636
rect 15105 9639 15163 9645
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 15930 9636 15936 9648
rect 15151 9608 15936 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 15930 9596 15936 9608
rect 15988 9596 15994 9648
rect 16040 9636 16068 9676
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 18046 9704 18052 9716
rect 16264 9676 18052 9704
rect 16264 9664 16270 9676
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 19886 9664 19892 9716
rect 19944 9664 19950 9716
rect 20990 9704 20996 9716
rect 20364 9676 20996 9704
rect 17310 9636 17316 9648
rect 16040 9608 17316 9636
rect 17310 9596 17316 9608
rect 17368 9636 17374 9648
rect 17368 9608 17632 9636
rect 17368 9596 17374 9608
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11422 9568 11428 9580
rect 11287 9540 11428 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 8662 9460 8668 9512
rect 8720 9460 8726 9512
rect 10686 9460 10692 9512
rect 10744 9500 10750 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10744 9472 10885 9500
rect 10744 9460 10750 9472
rect 10873 9469 10885 9472
rect 10919 9500 10931 9503
rect 11072 9500 11100 9531
rect 11422 9528 11428 9540
rect 11480 9568 11486 9580
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 11480 9540 12817 9568
rect 11480 9528 11486 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 12805 9531 12863 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9568 13047 9571
rect 13078 9568 13084 9580
rect 13035 9540 13084 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 10919 9472 11100 9500
rect 12820 9500 12848 9531
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 14148 9540 14841 9568
rect 14148 9528 14154 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15528 9540 15577 9568
rect 15528 9528 15534 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 15657 9571 15715 9577
rect 15657 9537 15669 9571
rect 15703 9568 15715 9571
rect 15746 9568 15752 9580
rect 15703 9540 15752 9568
rect 15703 9537 15715 9540
rect 15657 9531 15715 9537
rect 15746 9528 15752 9540
rect 15804 9568 15810 9580
rect 16942 9568 16948 9580
rect 15804 9540 16948 9568
rect 15804 9528 15810 9540
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17604 9577 17632 9608
rect 17770 9596 17776 9648
rect 17828 9596 17834 9648
rect 18064 9636 18092 9664
rect 20254 9636 20260 9648
rect 18064 9608 20260 9636
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 17221 9571 17279 9577
rect 17221 9537 17233 9571
rect 17267 9568 17279 9571
rect 17589 9571 17647 9577
rect 17267 9540 17540 9568
rect 17267 9537 17279 9540
rect 17221 9531 17279 9537
rect 13170 9500 13176 9512
rect 12820 9472 13176 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 17313 9503 17371 9509
rect 14424 9472 15148 9500
rect 14424 9460 14430 9472
rect 6748 9404 7328 9432
rect 7837 9435 7895 9441
rect 5684 9392 5690 9404
rect 7837 9401 7849 9435
rect 7883 9432 7895 9435
rect 8680 9432 8708 9460
rect 7883 9404 8708 9432
rect 7883 9401 7895 9404
rect 7837 9395 7895 9401
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 13446 9432 13452 9444
rect 9824 9404 13452 9432
rect 9824 9392 9830 9404
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 15120 9441 15148 9472
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 15105 9435 15163 9441
rect 15105 9401 15117 9435
rect 15151 9401 15163 9435
rect 17328 9432 17356 9463
rect 17402 9460 17408 9512
rect 17460 9460 17466 9512
rect 17512 9500 17540 9540
rect 17589 9537 17601 9571
rect 17635 9537 17647 9571
rect 17589 9531 17647 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9568 19579 9571
rect 19702 9568 19708 9580
rect 19567 9540 19708 9568
rect 19567 9537 19579 9540
rect 19521 9531 19579 9537
rect 19702 9528 19708 9540
rect 19760 9568 19766 9580
rect 20364 9577 20392 9676
rect 20990 9664 20996 9676
rect 21048 9704 21054 9716
rect 22278 9704 22284 9716
rect 21048 9676 22284 9704
rect 21048 9664 21054 9676
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 22370 9664 22376 9716
rect 22428 9664 22434 9716
rect 24394 9596 24400 9648
rect 24452 9596 24458 9648
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 19760 9540 20361 9568
rect 19760 9528 19766 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 20530 9528 20536 9580
rect 20588 9528 20594 9580
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9568 21879 9571
rect 21867 9540 21956 9568
rect 21867 9537 21879 9540
rect 21821 9531 21879 9537
rect 18322 9500 18328 9512
rect 17512 9472 18328 9500
rect 18322 9460 18328 9472
rect 18380 9500 18386 9512
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 18380 9472 19625 9500
rect 18380 9460 18386 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 20257 9503 20315 9509
rect 20257 9469 20269 9503
rect 20303 9500 20315 9503
rect 20548 9500 20576 9528
rect 21928 9512 21956 9540
rect 22066 9540 23152 9568
rect 20303 9472 20576 9500
rect 20303 9469 20315 9472
rect 20257 9463 20315 9469
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 18966 9432 18972 9444
rect 17328 9404 18972 9432
rect 15105 9395 15163 9401
rect 18966 9392 18972 9404
rect 19024 9392 19030 9444
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 19981 9435 20039 9441
rect 19981 9432 19993 9435
rect 19484 9404 19993 9432
rect 19484 9392 19490 9404
rect 19981 9401 19993 9404
rect 20027 9401 20039 9435
rect 19981 9395 20039 9401
rect 21818 9392 21824 9444
rect 21876 9432 21882 9444
rect 22066 9432 22094 9540
rect 23124 9509 23152 9540
rect 23017 9503 23075 9509
rect 23017 9469 23029 9503
rect 23063 9469 23075 9503
rect 23017 9463 23075 9469
rect 23109 9503 23167 9509
rect 23109 9469 23121 9503
rect 23155 9469 23167 9503
rect 23109 9463 23167 9469
rect 23032 9432 23060 9463
rect 23382 9460 23388 9512
rect 23440 9460 23446 9512
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9500 24915 9503
rect 24946 9500 24952 9512
rect 24903 9472 24952 9500
rect 24903 9469 24915 9472
rect 24857 9463 24915 9469
rect 24946 9460 24952 9472
rect 25004 9500 25010 9512
rect 25590 9500 25596 9512
rect 25004 9472 25596 9500
rect 25004 9460 25010 9472
rect 25590 9460 25596 9472
rect 25648 9460 25654 9512
rect 21876 9404 22094 9432
rect 22204 9404 23060 9432
rect 21876 9392 21882 9404
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 6270 9364 6276 9376
rect 5583 9336 6276 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10781 9367 10839 9373
rect 10781 9364 10793 9367
rect 10376 9336 10793 9364
rect 10376 9324 10382 9336
rect 10781 9333 10793 9336
rect 10827 9333 10839 9367
rect 10781 9327 10839 9333
rect 19705 9367 19763 9373
rect 19705 9333 19717 9367
rect 19751 9364 19763 9367
rect 20162 9364 20168 9376
rect 19751 9336 20168 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 20162 9324 20168 9336
rect 20220 9364 20226 9376
rect 20349 9367 20407 9373
rect 20349 9364 20361 9367
rect 20220 9336 20361 9364
rect 20220 9324 20226 9336
rect 20349 9333 20361 9336
rect 20395 9364 20407 9367
rect 21450 9364 21456 9376
rect 20395 9336 21456 9364
rect 20395 9333 20407 9336
rect 20349 9327 20407 9333
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 22097 9367 22155 9373
rect 22097 9333 22109 9367
rect 22143 9364 22155 9367
rect 22204 9364 22232 9404
rect 22143 9336 22232 9364
rect 22143 9333 22155 9336
rect 22097 9327 22155 9333
rect 22278 9324 22284 9376
rect 22336 9324 22342 9376
rect 23032 9364 23060 9404
rect 23566 9364 23572 9376
rect 23032 9336 23572 9364
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 24946 9324 24952 9376
rect 25004 9324 25010 9376
rect 1104 9274 30820 9296
rect 1104 9222 4664 9274
rect 4716 9222 4728 9274
rect 4780 9222 4792 9274
rect 4844 9222 4856 9274
rect 4908 9222 4920 9274
rect 4972 9222 12092 9274
rect 12144 9222 12156 9274
rect 12208 9222 12220 9274
rect 12272 9222 12284 9274
rect 12336 9222 12348 9274
rect 12400 9222 19520 9274
rect 19572 9222 19584 9274
rect 19636 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 26948 9274
rect 27000 9222 27012 9274
rect 27064 9222 27076 9274
rect 27128 9222 27140 9274
rect 27192 9222 27204 9274
rect 27256 9222 30820 9274
rect 1104 9200 30820 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 4430 9160 4436 9172
rect 1627 9132 4436 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4580 9132 4629 9160
rect 4580 9120 4586 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 4617 9123 4675 9129
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5960 9132 6101 9160
rect 5960 9120 5966 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 7374 9160 7380 9172
rect 6328 9132 7380 9160
rect 6328 9120 6334 9132
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 8754 9160 8760 9172
rect 7524 9132 8760 9160
rect 7524 9120 7530 9132
rect 8754 9120 8760 9132
rect 8812 9120 8818 9172
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 11422 9120 11428 9172
rect 11480 9120 11486 9172
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9160 17003 9163
rect 17034 9160 17040 9172
rect 16991 9132 17040 9160
rect 16991 9129 17003 9132
rect 16945 9123 17003 9129
rect 17034 9120 17040 9132
rect 17092 9120 17098 9172
rect 18322 9120 18328 9172
rect 18380 9120 18386 9172
rect 18966 9120 18972 9172
rect 19024 9160 19030 9172
rect 19429 9163 19487 9169
rect 19429 9160 19441 9163
rect 19024 9132 19441 9160
rect 19024 9120 19030 9132
rect 19429 9129 19441 9132
rect 19475 9160 19487 9163
rect 20806 9160 20812 9172
rect 19475 9132 20812 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 21910 9120 21916 9172
rect 21968 9120 21974 9172
rect 22278 9120 22284 9172
rect 22336 9120 22342 9172
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 22465 9163 22523 9169
rect 22465 9160 22477 9163
rect 22428 9132 22477 9160
rect 22428 9120 22434 9132
rect 22465 9129 22477 9132
rect 22511 9129 22523 9163
rect 22465 9123 22523 9129
rect 23293 9163 23351 9169
rect 23293 9129 23305 9163
rect 23339 9160 23351 9163
rect 23382 9160 23388 9172
rect 23339 9132 23388 9160
rect 23339 9129 23351 9132
rect 23293 9123 23351 9129
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 23750 9120 23756 9172
rect 23808 9120 23814 9172
rect 24486 9120 24492 9172
rect 24544 9120 24550 9172
rect 24946 9120 24952 9172
rect 25004 9120 25010 9172
rect 30374 9120 30380 9172
rect 30432 9120 30438 9172
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9092 5871 9095
rect 6362 9092 6368 9104
rect 5859 9064 6368 9092
rect 5859 9061 5871 9064
rect 5813 9055 5871 9061
rect 6362 9052 6368 9064
rect 6420 9092 6426 9104
rect 6822 9092 6828 9104
rect 6420 9064 6828 9092
rect 6420 9052 6426 9064
rect 6822 9052 6828 9064
rect 6880 9052 6886 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 9030 9092 9036 9104
rect 8527 9064 9036 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 9030 9052 9036 9064
rect 9088 9052 9094 9104
rect 9600 9064 9720 9092
rect 6086 9024 6092 9036
rect 6012 8996 6092 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 4246 8916 4252 8968
rect 4304 8956 4310 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 4304 8928 4721 8956
rect 4304 8916 4310 8928
rect 4709 8925 4721 8928
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 4724 8888 4752 8919
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 6012 8965 6040 8996
rect 6086 8984 6092 8996
rect 6144 9024 6150 9036
rect 6144 8996 6316 9024
rect 6144 8984 6150 8996
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5040 8928 5733 8956
rect 5040 8916 5046 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5721 8919 5779 8925
rect 5920 8928 6009 8956
rect 5920 8900 5948 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5997 8919 6055 8925
rect 6104 8928 6193 8956
rect 5166 8888 5172 8900
rect 4724 8860 5172 8888
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 5902 8848 5908 8900
rect 5960 8848 5966 8900
rect 6104 8832 6132 8928
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 6288 8956 6316 8996
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 6696 8996 8033 9024
rect 6696 8984 6702 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 9024 8447 9027
rect 9600 9024 9628 9064
rect 8435 8996 8524 9024
rect 8435 8993 8447 8996
rect 8389 8987 8447 8993
rect 8496 8968 8524 8996
rect 9324 8996 9628 9024
rect 9692 9024 9720 9064
rect 9950 9052 9956 9104
rect 10008 9092 10014 9104
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 10008 9064 10149 9092
rect 10008 9052 10014 9064
rect 10137 9061 10149 9064
rect 10183 9061 10195 9095
rect 10336 9092 10364 9120
rect 10336 9064 10916 9092
rect 10137 9055 10195 9061
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 9692 8996 10517 9024
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6288 8928 7573 8956
rect 6181 8919 6239 8925
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 8478 8916 8484 8968
rect 8536 8916 8542 8968
rect 8610 8959 8668 8965
rect 8610 8925 8622 8959
rect 8656 8956 8668 8959
rect 9214 8956 9220 8968
rect 8656 8928 9220 8956
rect 8656 8925 8668 8928
rect 8610 8919 8668 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9324 8965 9352 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 9950 8916 9956 8968
rect 10008 8956 10014 8968
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10008 8928 10425 8956
rect 10008 8916 10014 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 7929 8891 7987 8897
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 7975 8860 8769 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 8757 8857 8769 8860
rect 8803 8857 8815 8891
rect 8757 8851 8815 8857
rect 6086 8780 6092 8832
rect 6144 8780 6150 8832
rect 7760 8820 7788 8851
rect 9398 8848 9404 8900
rect 9456 8848 9462 8900
rect 9490 8848 9496 8900
rect 9548 8848 9554 8900
rect 9674 8897 9680 8900
rect 9631 8891 9680 8897
rect 9631 8888 9643 8891
rect 9587 8860 9643 8888
rect 9631 8857 9643 8860
rect 9677 8857 9680 8891
rect 9631 8851 9680 8857
rect 9674 8848 9680 8851
rect 9732 8848 9738 8900
rect 9861 8891 9919 8897
rect 9861 8857 9873 8891
rect 9907 8888 9919 8891
rect 10612 8888 10640 8919
rect 10686 8916 10692 8968
rect 10744 8916 10750 8968
rect 10888 8965 10916 9064
rect 11440 8965 11468 9120
rect 13265 9095 13323 9101
rect 13265 9092 13277 9095
rect 12406 9064 13277 9092
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 11790 8956 11796 8968
rect 11655 8928 11796 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 12406 8888 12434 9064
rect 13265 9061 13277 9064
rect 13311 9061 13323 9095
rect 17126 9092 17132 9104
rect 13265 9055 13323 9061
rect 15304 9064 17132 9092
rect 15304 9033 15332 9064
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 17218 9052 17224 9104
rect 17276 9092 17282 9104
rect 18141 9095 18199 9101
rect 18141 9092 18153 9095
rect 17276 9064 18153 9092
rect 17276 9052 17282 9064
rect 18141 9061 18153 9064
rect 18187 9092 18199 9095
rect 18785 9095 18843 9101
rect 18785 9092 18797 9095
rect 18187 9064 18797 9092
rect 18187 9061 18199 9064
rect 18141 9055 18199 9061
rect 18785 9061 18797 9064
rect 18831 9061 18843 9095
rect 18785 9055 18843 9061
rect 19245 9095 19303 9101
rect 19245 9061 19257 9095
rect 19291 9061 19303 9095
rect 19245 9055 19303 9061
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 12728 8996 13829 9024
rect 12728 8965 12756 8996
rect 13817 8993 13829 8996
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 15289 9027 15347 9033
rect 15289 8993 15301 9027
rect 15335 8993 15347 9027
rect 15289 8987 15347 8993
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 9024 15623 9027
rect 15654 9024 15660 9036
rect 15611 8996 15660 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 15654 8984 15660 8996
rect 15712 9024 15718 9036
rect 17957 9027 18015 9033
rect 15712 8996 17632 9024
rect 15712 8984 15718 8996
rect 12713 8959 12771 8965
rect 12713 8925 12725 8959
rect 12759 8925 12771 8959
rect 12713 8919 12771 8925
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8956 13231 8959
rect 13354 8956 13360 8968
rect 13219 8928 13360 8956
rect 13219 8925 13231 8928
rect 13173 8919 13231 8925
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 13495 8928 13737 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 9907 8860 10456 8888
rect 10612 8860 12817 8888
rect 9907 8857 9919 8860
rect 9861 8851 9919 8857
rect 10428 8832 10456 8860
rect 12805 8857 12817 8860
rect 12851 8857 12863 8891
rect 13015 8891 13073 8897
rect 13015 8888 13027 8891
rect 12805 8851 12863 8857
rect 12912 8860 13027 8888
rect 7834 8820 7840 8832
rect 7760 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 9122 8780 9128 8832
rect 9180 8780 9186 8832
rect 10410 8780 10416 8832
rect 10468 8780 10474 8832
rect 10781 8823 10839 8829
rect 10781 8789 10793 8823
rect 10827 8820 10839 8823
rect 10962 8820 10968 8832
rect 10827 8792 10968 8820
rect 10827 8789 10839 8792
rect 10781 8783 10839 8789
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 11296 8792 11529 8820
rect 11296 8780 11302 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 12526 8780 12532 8832
rect 12584 8780 12590 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 12912 8820 12940 8860
rect 13015 8857 13027 8860
rect 13061 8857 13073 8891
rect 13015 8851 13073 8857
rect 13464 8832 13492 8919
rect 13906 8916 13912 8968
rect 13964 8916 13970 8968
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15838 8956 15844 8968
rect 15252 8928 15844 8956
rect 15252 8916 15258 8928
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 17221 8959 17279 8965
rect 17132 8937 17190 8943
rect 13633 8891 13691 8897
rect 13633 8857 13645 8891
rect 13679 8888 13691 8891
rect 13924 8888 13952 8916
rect 17132 8903 17144 8937
rect 17178 8903 17190 8937
rect 17221 8925 17233 8959
rect 17267 8956 17279 8959
rect 17310 8956 17316 8968
rect 17267 8928 17316 8956
rect 17267 8925 17279 8928
rect 17221 8919 17279 8925
rect 17310 8916 17316 8928
rect 17368 8916 17374 8968
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17604 8956 17632 8996
rect 17957 8993 17969 9027
rect 18003 9024 18015 9027
rect 18046 9024 18052 9036
rect 18003 8996 18052 9024
rect 18003 8993 18015 8996
rect 17957 8987 18015 8993
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 19260 9024 19288 9055
rect 20530 9052 20536 9104
rect 20588 9052 20594 9104
rect 22296 9092 22324 9120
rect 22296 9064 22600 9092
rect 18248 8996 19288 9024
rect 18248 8965 18276 8996
rect 20070 8984 20076 9036
rect 20128 8984 20134 9036
rect 20165 9027 20223 9033
rect 20165 8993 20177 9027
rect 20211 9024 20223 9027
rect 20211 8996 21036 9024
rect 20211 8993 20223 8996
rect 20165 8987 20223 8993
rect 18233 8959 18291 8965
rect 17604 8928 18092 8956
rect 17132 8900 17190 8903
rect 13679 8860 13952 8888
rect 13679 8857 13691 8860
rect 13633 8851 13691 8857
rect 17126 8848 17132 8900
rect 17184 8848 17190 8900
rect 18064 8888 18092 8928
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18966 8916 18972 8968
rect 19024 8916 19030 8968
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8956 19119 8959
rect 19426 8956 19432 8968
rect 19107 8928 19432 8956
rect 19107 8925 19119 8928
rect 19061 8919 19119 8925
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 18509 8891 18567 8897
rect 18509 8888 18521 8891
rect 18064 8860 18521 8888
rect 18509 8857 18521 8860
rect 18555 8857 18567 8891
rect 18509 8851 18567 8857
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 18693 8891 18751 8897
rect 18693 8888 18705 8891
rect 18656 8860 18705 8888
rect 18656 8848 18662 8860
rect 18693 8857 18705 8860
rect 18739 8888 18751 8891
rect 18785 8891 18843 8897
rect 18785 8888 18797 8891
rect 18739 8860 18797 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 18785 8857 18797 8860
rect 18831 8888 18843 8891
rect 19613 8891 19671 8897
rect 19613 8888 19625 8891
rect 18831 8860 19625 8888
rect 18831 8857 18843 8860
rect 18785 8851 18843 8857
rect 19613 8857 19625 8860
rect 19659 8857 19671 8891
rect 19613 8851 19671 8857
rect 12676 8792 12940 8820
rect 12676 8780 12682 8792
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 18230 8780 18236 8832
rect 18288 8780 18294 8832
rect 19426 8829 19432 8832
rect 19413 8823 19432 8829
rect 19413 8789 19425 8823
rect 19413 8783 19432 8789
rect 19426 8780 19432 8783
rect 19484 8780 19490 8832
rect 19886 8780 19892 8832
rect 19944 8780 19950 8832
rect 20088 8820 20116 8984
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20180 8928 20269 8956
rect 20180 8900 20208 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20438 8956 20444 8968
rect 20395 8928 20444 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 20438 8916 20444 8928
rect 20496 8916 20502 8968
rect 20732 8965 20760 8996
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8925 20775 8959
rect 20717 8919 20775 8925
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 21008 8956 21036 8996
rect 21634 8984 21640 9036
rect 21692 9024 21698 9036
rect 21692 8996 22416 9024
rect 21692 8984 21698 8996
rect 21652 8956 21680 8984
rect 22388 8965 22416 8996
rect 22572 8965 22600 9064
rect 23566 9052 23572 9104
rect 23624 9052 23630 9104
rect 24504 9092 24532 9120
rect 23676 9064 24532 9092
rect 23584 9024 23612 9052
rect 23400 8996 23612 9024
rect 21008 8928 21680 8956
rect 22097 8959 22155 8965
rect 20809 8919 20867 8925
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22373 8959 22431 8965
rect 22373 8925 22385 8959
rect 22419 8925 22431 8959
rect 22373 8919 22431 8925
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 20162 8848 20168 8900
rect 20220 8888 20226 8900
rect 20533 8891 20591 8897
rect 20533 8888 20545 8891
rect 20220 8860 20545 8888
rect 20220 8848 20226 8860
rect 20533 8857 20545 8860
rect 20579 8857 20591 8891
rect 20533 8851 20591 8857
rect 20824 8820 20852 8919
rect 22112 8888 22140 8919
rect 23400 8888 23428 8996
rect 23474 8916 23480 8968
rect 23532 8916 23538 8968
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8956 23627 8959
rect 23676 8956 23704 9064
rect 23615 8928 23704 8956
rect 23845 8959 23903 8965
rect 23615 8925 23627 8928
rect 23569 8919 23627 8925
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24964 8956 24992 9120
rect 23891 8928 24992 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 25590 8916 25596 8968
rect 25648 8956 25654 8968
rect 30193 8959 30251 8965
rect 30193 8956 30205 8959
rect 25648 8928 30205 8956
rect 25648 8916 25654 8928
rect 30193 8925 30205 8928
rect 30239 8925 30251 8959
rect 30193 8919 30251 8925
rect 22112 8860 23428 8888
rect 20088 8792 20852 8820
rect 1104 8730 30820 8752
rect 1104 8678 5324 8730
rect 5376 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 12752 8730
rect 12804 8678 12816 8730
rect 12868 8678 12880 8730
rect 12932 8678 12944 8730
rect 12996 8678 13008 8730
rect 13060 8678 20180 8730
rect 20232 8678 20244 8730
rect 20296 8678 20308 8730
rect 20360 8678 20372 8730
rect 20424 8678 20436 8730
rect 20488 8678 27608 8730
rect 27660 8678 27672 8730
rect 27724 8678 27736 8730
rect 27788 8678 27800 8730
rect 27852 8678 27864 8730
rect 27916 8678 30820 8730
rect 1104 8656 30820 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 5902 8616 5908 8628
rect 1627 8588 5908 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 7009 8619 7067 8625
rect 7009 8585 7021 8619
rect 7055 8616 7067 8619
rect 7650 8616 7656 8628
rect 7055 8588 7656 8616
rect 7055 8585 7067 8588
rect 7009 8579 7067 8585
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8128 8588 9045 8616
rect 5813 8551 5871 8557
rect 5813 8517 5825 8551
rect 5859 8517 5871 8551
rect 5813 8511 5871 8517
rect 6029 8551 6087 8557
rect 6029 8517 6041 8551
rect 6075 8548 6087 8551
rect 6546 8548 6552 8560
rect 6075 8520 6552 8548
rect 6075 8517 6087 8520
rect 6029 8511 6087 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 5828 8480 5856 8511
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 8128 8557 8156 8588
rect 9033 8585 9045 8588
rect 9079 8616 9091 8619
rect 9398 8616 9404 8628
rect 9079 8588 9404 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10413 8619 10471 8625
rect 9548 8588 10364 8616
rect 9548 8576 9554 8588
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 7760 8520 8125 8548
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 5828 8452 6040 8480
rect 6012 8424 6040 8452
rect 6196 8452 7297 8480
rect 5994 8372 6000 8424
rect 6052 8372 6058 8424
rect 6196 8353 6224 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7466 8480 7472 8492
rect 7423 8452 7472 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7650 8489 7656 8492
rect 7635 8483 7656 8489
rect 7635 8449 7647 8483
rect 7635 8443 7656 8449
rect 7650 8440 7656 8443
rect 7708 8440 7714 8492
rect 6362 8372 6368 8424
rect 6420 8372 6426 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7760 8412 7788 8520
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 9214 8508 9220 8560
rect 9272 8508 9278 8560
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 8076 8452 8217 8480
rect 8076 8440 8082 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 8352 8452 8401 8480
rect 8352 8440 8358 8452
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 9232 8480 9260 8508
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 9232 8452 9413 8480
rect 8389 8443 8447 8449
rect 9401 8449 9413 8452
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10336 8480 10364 8588
rect 10413 8585 10425 8619
rect 10459 8616 10471 8619
rect 10686 8616 10692 8628
rect 10459 8588 10692 8616
rect 10459 8585 10471 8588
rect 10413 8579 10471 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 12713 8619 12771 8625
rect 10796 8588 12434 8616
rect 10796 8480 10824 8588
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 12406 8548 12434 8588
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 13078 8616 13084 8628
rect 12759 8588 13084 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 15654 8576 15660 8628
rect 15712 8576 15718 8628
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16298 8616 16304 8628
rect 16071 8588 16304 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 17494 8576 17500 8628
rect 17552 8576 17558 8628
rect 19886 8576 19892 8628
rect 19944 8576 19950 8628
rect 20530 8576 20536 8628
rect 20588 8576 20594 8628
rect 20806 8576 20812 8628
rect 20864 8576 20870 8628
rect 21634 8576 21640 8628
rect 21692 8576 21698 8628
rect 24305 8619 24363 8625
rect 24305 8585 24317 8619
rect 24351 8616 24363 8619
rect 24394 8616 24400 8628
rect 24351 8588 24400 8616
rect 24351 8585 24363 8588
rect 24305 8579 24363 8585
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 13906 8548 13912 8560
rect 11020 8520 11192 8548
rect 12406 8520 13912 8548
rect 11020 8508 11026 8520
rect 11164 8489 11192 8520
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 9732 8452 10272 8480
rect 10336 8452 10824 8480
rect 11149 8483 11207 8489
rect 9732 8440 9738 8452
rect 6788 8384 7788 8412
rect 6788 8372 6794 8384
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8536 8384 9321 8412
rect 8536 8372 8542 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8313 6239 8347
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 6181 8307 6239 8313
rect 6656 8316 7757 8344
rect 5997 8279 6055 8285
rect 5997 8245 6009 8279
rect 6043 8276 6055 8279
rect 6086 8276 6092 8288
rect 6043 8248 6092 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6086 8236 6092 8248
rect 6144 8276 6150 8288
rect 6656 8276 6684 8316
rect 7745 8313 7757 8316
rect 7791 8313 7803 8347
rect 7745 8307 7803 8313
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 8386 8344 8392 8356
rect 8343 8316 8392 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 9324 8288 9352 8375
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 9950 8412 9956 8424
rect 9640 8384 9956 8412
rect 9640 8372 9646 8384
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10244 8412 10272 8452
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11238 8440 11244 8492
rect 11296 8440 11302 8492
rect 13446 8480 13452 8492
rect 12544 8452 13452 8480
rect 11057 8415 11115 8421
rect 10244 8384 10824 8412
rect 10321 8347 10379 8353
rect 9646 8316 10272 8344
rect 6144 8248 6684 8276
rect 6144 8236 6150 8248
rect 7098 8236 7104 8288
rect 7156 8236 7162 8288
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7561 8279 7619 8285
rect 7561 8276 7573 8279
rect 7432 8248 7573 8276
rect 7432 8236 7438 8248
rect 7561 8245 7573 8248
rect 7607 8245 7619 8279
rect 7561 8239 7619 8245
rect 9030 8236 9036 8288
rect 9088 8276 9094 8288
rect 9214 8276 9220 8288
rect 9088 8248 9220 8276
rect 9088 8236 9094 8248
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9646 8276 9674 8316
rect 9364 8248 9674 8276
rect 10244 8276 10272 8316
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 10410 8344 10416 8356
rect 10367 8316 10416 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10796 8353 10824 8384
rect 11057 8381 11069 8415
rect 11103 8412 11115 8415
rect 11256 8412 11284 8440
rect 11103 8384 11284 8412
rect 11103 8381 11115 8384
rect 11057 8375 11115 8381
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8313 10839 8347
rect 12544 8344 12572 8452
rect 13446 8440 13452 8452
rect 13504 8480 13510 8492
rect 15672 8489 15700 8576
rect 17512 8548 17540 8576
rect 17681 8551 17739 8557
rect 17681 8548 17693 8551
rect 17512 8520 17693 8548
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13504 8452 13737 8480
rect 13504 8440 13510 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17218 8480 17224 8492
rect 17083 8452 17224 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 17512 8489 17540 8520
rect 17681 8517 17693 8520
rect 17727 8517 17739 8551
rect 17681 8511 17739 8517
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8480 17831 8483
rect 17862 8480 17868 8492
rect 17819 8452 17868 8480
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 12676 8384 13185 8412
rect 12676 8372 12682 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 15795 8384 16865 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 17328 8412 17356 8443
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 17954 8440 17960 8492
rect 18012 8440 18018 8492
rect 19904 8480 19932 8576
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19904 8452 19993 8480
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8480 20131 8483
rect 20548 8480 20576 8576
rect 20119 8452 20576 8480
rect 20993 8483 21051 8489
rect 20119 8449 20131 8452
rect 20073 8443 20131 8449
rect 20993 8449 21005 8483
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 17402 8412 17408 8424
rect 17328 8384 17408 8412
rect 16853 8375 16911 8381
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 10781 8307 10839 8313
rect 10888 8316 12817 8344
rect 10888 8276 10916 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 13188 8344 13216 8375
rect 17402 8372 17408 8384
rect 17460 8412 17466 8424
rect 17972 8412 18000 8440
rect 17460 8384 18000 8412
rect 19797 8415 19855 8421
rect 17460 8372 17466 8384
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 20622 8412 20628 8424
rect 19843 8384 20628 8412
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 13357 8347 13415 8353
rect 13357 8344 13369 8347
rect 13188 8316 13369 8344
rect 12805 8307 12863 8313
rect 13357 8313 13369 8316
rect 13403 8313 13415 8347
rect 21008 8344 21036 8443
rect 21174 8440 21180 8492
rect 21232 8440 21238 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21652 8480 21680 8576
rect 22094 8508 22100 8560
rect 22152 8508 22158 8560
rect 23106 8508 23112 8560
rect 23164 8508 23170 8560
rect 21315 8452 21680 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 24397 8483 24455 8489
rect 24397 8480 24409 8483
rect 23716 8452 24409 8480
rect 23716 8440 23722 8452
rect 24397 8449 24409 8452
rect 24443 8480 24455 8483
rect 24854 8480 24860 8492
rect 24443 8452 24860 8480
rect 24443 8449 24455 8452
rect 24397 8443 24455 8449
rect 24854 8440 24860 8452
rect 24912 8440 24918 8492
rect 30193 8483 30251 8489
rect 30193 8449 30205 8483
rect 30239 8449 30251 8483
rect 30193 8443 30251 8449
rect 21082 8372 21088 8424
rect 21140 8412 21146 8424
rect 21818 8412 21824 8424
rect 21140 8384 21824 8412
rect 21140 8372 21146 8384
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 22186 8412 22192 8424
rect 21928 8384 22192 8412
rect 21928 8344 21956 8384
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 30208 8412 30236 8443
rect 23624 8384 30236 8412
rect 23624 8372 23630 8384
rect 21008 8316 21956 8344
rect 13357 8307 13415 8313
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 30377 8347 30435 8353
rect 30377 8344 30389 8347
rect 30340 8316 30389 8344
rect 30340 8304 30346 8316
rect 30377 8313 30389 8316
rect 30423 8313 30435 8347
rect 30377 8307 30435 8313
rect 10244 8248 10916 8276
rect 19889 8279 19947 8285
rect 9364 8236 9370 8248
rect 19889 8245 19901 8279
rect 19935 8276 19947 8279
rect 19978 8276 19984 8288
rect 19935 8248 19984 8276
rect 19935 8245 19947 8248
rect 19889 8239 19947 8245
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 1104 8186 30820 8208
rect 1104 8134 4664 8186
rect 4716 8134 4728 8186
rect 4780 8134 4792 8186
rect 4844 8134 4856 8186
rect 4908 8134 4920 8186
rect 4972 8134 12092 8186
rect 12144 8134 12156 8186
rect 12208 8134 12220 8186
rect 12272 8134 12284 8186
rect 12336 8134 12348 8186
rect 12400 8134 19520 8186
rect 19572 8134 19584 8186
rect 19636 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 26948 8186
rect 27000 8134 27012 8186
rect 27064 8134 27076 8186
rect 27128 8134 27140 8186
rect 27192 8134 27204 8186
rect 27256 8134 30820 8186
rect 1104 8112 30820 8134
rect 6362 8072 6368 8084
rect 4724 8044 6368 8072
rect 4724 7945 4752 8044
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6604 8044 6653 8072
rect 6604 8032 6610 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 7377 8075 7435 8081
rect 7377 8041 7389 8075
rect 7423 8041 7435 8075
rect 7377 8035 7435 8041
rect 6380 8004 6408 8032
rect 7392 8004 7420 8035
rect 7926 8032 7932 8084
rect 7984 8032 7990 8084
rect 8294 8032 8300 8084
rect 8352 8032 8358 8084
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17644 8044 17785 8072
rect 17644 8032 17650 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 18509 8075 18567 8081
rect 18509 8041 18521 8075
rect 18555 8072 18567 8075
rect 18598 8072 18604 8084
rect 18555 8044 18604 8072
rect 18555 8041 18567 8044
rect 18509 8035 18567 8041
rect 6380 7976 7420 8004
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 1688 7908 4721 7936
rect 1688 7877 1716 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 6181 7939 6239 7945
rect 6181 7905 6193 7939
rect 6227 7936 6239 7939
rect 7098 7936 7104 7948
rect 6227 7908 7104 7936
rect 6227 7905 6239 7908
rect 6181 7899 6239 7905
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 5718 7760 5724 7812
rect 5776 7760 5782 7812
rect 6564 7800 6592 7831
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7392 7868 7420 7976
rect 7745 8007 7803 8013
rect 7745 7973 7757 8007
rect 7791 8004 7803 8007
rect 7834 8004 7840 8016
rect 7791 7976 7840 8004
rect 7791 7973 7803 7976
rect 7745 7967 7803 7973
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7392 7840 7849 7868
rect 7285 7831 7343 7837
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7300 7800 7328 7831
rect 7944 7800 7972 8032
rect 17788 8004 17816 8035
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8041 20223 8075
rect 20165 8035 20223 8041
rect 19334 8004 19340 8016
rect 17788 7976 19340 8004
rect 19334 7964 19340 7976
rect 19392 8004 19398 8016
rect 20180 8004 20208 8035
rect 21174 8032 21180 8084
rect 21232 8032 21238 8084
rect 21358 8032 21364 8084
rect 21416 8032 21422 8084
rect 21450 8032 21456 8084
rect 21508 8072 21514 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 21508 8044 21833 8072
rect 21508 8032 21514 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22373 8075 22431 8081
rect 22373 8072 22385 8075
rect 22244 8044 22385 8072
rect 22244 8032 22250 8044
rect 22373 8041 22385 8044
rect 22419 8041 22431 8075
rect 22373 8035 22431 8041
rect 23017 8075 23075 8081
rect 23017 8041 23029 8075
rect 23063 8072 23075 8075
rect 23106 8072 23112 8084
rect 23063 8044 23112 8072
rect 23063 8041 23075 8044
rect 23017 8035 23075 8041
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 19392 7976 20208 8004
rect 21192 8004 21220 8032
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 21192 7976 21741 8004
rect 19392 7964 19398 7976
rect 21729 7973 21741 7976
rect 21775 8004 21787 8007
rect 21775 7976 21864 8004
rect 21775 7973 21787 7976
rect 21729 7967 21787 7973
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12584 7908 12633 7936
rect 12584 7896 12590 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12805 7939 12863 7945
rect 12805 7905 12817 7939
rect 12851 7936 12863 7939
rect 13078 7936 13084 7948
rect 12851 7908 13084 7936
rect 12851 7905 12863 7908
rect 12805 7899 12863 7905
rect 13078 7896 13084 7908
rect 13136 7936 13142 7948
rect 16574 7936 16580 7948
rect 13136 7908 16580 7936
rect 13136 7896 13142 7908
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 17954 7896 17960 7948
rect 18012 7936 18018 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 18012 7908 18061 7936
rect 18012 7896 18018 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17678 7868 17684 7880
rect 17635 7840 17684 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 6380 7772 7972 7800
rect 17512 7800 17540 7831
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18141 7871 18199 7877
rect 18141 7868 18153 7871
rect 17920 7840 18153 7868
rect 17920 7828 17926 7840
rect 18141 7837 18153 7840
rect 18187 7868 18199 7871
rect 18414 7868 18420 7880
rect 18187 7840 18420 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 19886 7828 19892 7880
rect 19944 7828 19950 7880
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20533 7871 20591 7877
rect 20533 7868 20545 7871
rect 20303 7840 20545 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 20533 7837 20545 7840
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20990 7828 20996 7880
rect 21048 7868 21054 7880
rect 21085 7871 21143 7877
rect 21085 7868 21097 7871
rect 21048 7840 21097 7868
rect 21048 7828 21054 7840
rect 21085 7837 21097 7840
rect 21131 7868 21143 7871
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 21131 7840 21281 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 21269 7837 21281 7840
rect 21315 7837 21327 7871
rect 21836 7868 21864 7976
rect 21910 7964 21916 8016
rect 21968 8004 21974 8016
rect 22465 8007 22523 8013
rect 22465 8004 22477 8007
rect 21968 7976 22477 8004
rect 21968 7964 21974 7976
rect 22465 7973 22477 7976
rect 22511 7973 22523 8007
rect 22465 7967 22523 7973
rect 22281 7871 22339 7877
rect 22281 7868 22293 7871
rect 21836 7840 22293 7868
rect 21269 7831 21327 7837
rect 22281 7837 22293 7840
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23658 7868 23664 7880
rect 23155 7840 23664 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 18230 7800 18236 7812
rect 17512 7772 18236 7800
rect 6380 7744 6408 7772
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 21284 7800 21312 7831
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 21284 7772 22845 7800
rect 22833 7769 22845 7772
rect 22879 7769 22891 7803
rect 22833 7763 22891 7769
rect 934 7692 940 7744
rect 992 7732 998 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 992 7704 1501 7732
rect 992 7692 998 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 6362 7692 6368 7744
rect 6420 7692 6426 7744
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 12161 7735 12219 7741
rect 12161 7732 12173 7735
rect 12032 7704 12173 7732
rect 12032 7692 12038 7704
rect 12161 7701 12173 7704
rect 12207 7701 12219 7735
rect 12161 7695 12219 7701
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12618 7732 12624 7744
rect 12575 7704 12624 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17092 7704 17325 7732
rect 17092 7692 17098 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 19426 7692 19432 7744
rect 19484 7732 19490 7744
rect 19705 7735 19763 7741
rect 19705 7732 19717 7735
rect 19484 7704 19717 7732
rect 19484 7692 19490 7704
rect 19705 7701 19717 7704
rect 19751 7701 19763 7735
rect 19705 7695 19763 7701
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21910 7732 21916 7744
rect 21416 7704 21916 7732
rect 21416 7692 21422 7704
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 23124 7732 23152 7831
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 22336 7704 23152 7732
rect 22336 7692 22342 7704
rect 1104 7642 30820 7664
rect 1104 7590 5324 7642
rect 5376 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 12752 7642
rect 12804 7590 12816 7642
rect 12868 7590 12880 7642
rect 12932 7590 12944 7642
rect 12996 7590 13008 7642
rect 13060 7590 20180 7642
rect 20232 7590 20244 7642
rect 20296 7590 20308 7642
rect 20360 7590 20372 7642
rect 20424 7590 20436 7642
rect 20488 7590 27608 7642
rect 27660 7590 27672 7642
rect 27724 7590 27736 7642
rect 27788 7590 27800 7642
rect 27852 7590 27864 7642
rect 27916 7590 30820 7642
rect 1104 7568 30820 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7497 1639 7531
rect 1581 7491 1639 7497
rect 1596 7460 1624 7491
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 11514 7528 11520 7540
rect 6512 7500 11520 7528
rect 6512 7488 6518 7500
rect 6362 7460 6368 7472
rect 1596 7432 6368 7460
rect 6362 7420 6368 7432
rect 6420 7420 6426 7472
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5224 7364 5641 7392
rect 5224 7352 5230 7364
rect 5629 7361 5641 7364
rect 5675 7392 5687 7395
rect 5675 7364 6960 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 6932 7188 6960 7364
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8588 7401 8616 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 12434 7528 12440 7540
rect 11624 7500 12440 7528
rect 10505 7463 10563 7469
rect 10505 7460 10517 7463
rect 10074 7432 10517 7460
rect 10505 7429 10517 7432
rect 10551 7429 10563 7463
rect 11624 7460 11652 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12676 7500 13277 7528
rect 12676 7488 12682 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 13449 7463 13507 7469
rect 13449 7460 13461 7463
rect 10505 7423 10563 7429
rect 10612 7432 11652 7460
rect 13018 7432 13461 7460
rect 10612 7401 10640 7432
rect 13449 7429 13461 7432
rect 13495 7429 13507 7463
rect 13449 7423 13507 7429
rect 16945 7463 17003 7469
rect 16945 7429 16957 7463
rect 16991 7460 17003 7463
rect 17034 7460 17040 7472
rect 16991 7432 17040 7460
rect 16991 7429 17003 7432
rect 16945 7423 17003 7429
rect 17034 7420 17040 7432
rect 17092 7420 17098 7472
rect 19337 7463 19395 7469
rect 19337 7429 19349 7463
rect 19383 7460 19395 7463
rect 19426 7460 19432 7472
rect 19383 7432 19432 7460
rect 19383 7429 19395 7432
rect 19337 7423 19395 7429
rect 19426 7420 19432 7432
rect 19484 7420 19490 7472
rect 20070 7420 20076 7472
rect 20128 7420 20134 7472
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8496 7296 8861 7324
rect 8496 7265 8524 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 8481 7259 8539 7265
rect 8481 7225 8493 7259
rect 8527 7225 8539 7259
rect 10612 7256 10640 7355
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 11790 7284 11796 7336
rect 11848 7284 11854 7336
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 13372 7324 13400 7355
rect 12492 7296 13400 7324
rect 16684 7324 16712 7355
rect 18046 7352 18052 7404
rect 18104 7352 18110 7404
rect 19061 7395 19119 7401
rect 19061 7361 19073 7395
rect 19107 7361 19119 7395
rect 19061 7355 19119 7361
rect 19076 7324 19104 7355
rect 21082 7324 21088 7336
rect 16684 7296 21088 7324
rect 12492 7284 12498 7296
rect 21082 7284 21088 7296
rect 21140 7284 21146 7336
rect 8481 7219 8539 7225
rect 9876 7228 10640 7256
rect 9876 7188 9904 7228
rect 6932 7160 9904 7188
rect 10321 7191 10379 7197
rect 10321 7157 10333 7191
rect 10367 7188 10379 7191
rect 10410 7188 10416 7200
rect 10367 7160 10416 7188
rect 10367 7157 10379 7160
rect 10321 7151 10379 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 18414 7148 18420 7200
rect 18472 7148 18478 7200
rect 20809 7191 20867 7197
rect 20809 7157 20821 7191
rect 20855 7188 20867 7191
rect 20990 7188 20996 7200
rect 20855 7160 20996 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 1104 7098 30820 7120
rect 1104 7046 4664 7098
rect 4716 7046 4728 7098
rect 4780 7046 4792 7098
rect 4844 7046 4856 7098
rect 4908 7046 4920 7098
rect 4972 7046 12092 7098
rect 12144 7046 12156 7098
rect 12208 7046 12220 7098
rect 12272 7046 12284 7098
rect 12336 7046 12348 7098
rect 12400 7046 19520 7098
rect 19572 7046 19584 7098
rect 19636 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 26948 7098
rect 27000 7046 27012 7098
rect 27064 7046 27076 7098
rect 27128 7046 27140 7098
rect 27192 7046 27204 7098
rect 27256 7046 30820 7098
rect 1104 7024 30820 7046
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8352 6956 8953 6984
rect 8352 6944 8358 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 11885 6987 11943 6993
rect 11885 6984 11897 6987
rect 11848 6956 11897 6984
rect 11848 6944 11854 6956
rect 11885 6953 11897 6956
rect 11931 6953 11943 6987
rect 11885 6947 11943 6953
rect 20070 6944 20076 6996
rect 20128 6944 20134 6996
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 9180 6820 9413 6848
rect 9180 6808 9186 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 13078 6848 13084 6860
rect 9631 6820 13084 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 10410 6780 10416 6792
rect 9355 6752 10416 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12069 6783 12127 6789
rect 12069 6780 12081 6783
rect 12032 6752 12081 6780
rect 12032 6740 12038 6752
rect 12069 6749 12081 6752
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 17000 6752 17141 6780
rect 17000 6740 17006 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 18064 6780 18092 6808
rect 17267 6752 18092 6780
rect 19981 6783 20039 6789
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 22278 6780 22284 6792
rect 20027 6752 22284 6780
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 17144 6712 17172 6743
rect 19996 6712 20024 6743
rect 22278 6740 22284 6752
rect 22336 6740 22342 6792
rect 17144 6684 20024 6712
rect 1104 6554 30820 6576
rect 1104 6502 5324 6554
rect 5376 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 12752 6554
rect 12804 6502 12816 6554
rect 12868 6502 12880 6554
rect 12932 6502 12944 6554
rect 12996 6502 13008 6554
rect 13060 6502 20180 6554
rect 20232 6502 20244 6554
rect 20296 6502 20308 6554
rect 20360 6502 20372 6554
rect 20424 6502 20436 6554
rect 20488 6502 27608 6554
rect 27660 6502 27672 6554
rect 27724 6502 27736 6554
rect 27788 6502 27800 6554
rect 27852 6502 27864 6554
rect 27916 6502 30820 6554
rect 1104 6480 30820 6502
rect 1104 6010 30820 6032
rect 1104 5958 4664 6010
rect 4716 5958 4728 6010
rect 4780 5958 4792 6010
rect 4844 5958 4856 6010
rect 4908 5958 4920 6010
rect 4972 5958 12092 6010
rect 12144 5958 12156 6010
rect 12208 5958 12220 6010
rect 12272 5958 12284 6010
rect 12336 5958 12348 6010
rect 12400 5958 19520 6010
rect 19572 5958 19584 6010
rect 19636 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 26948 6010
rect 27000 5958 27012 6010
rect 27064 5958 27076 6010
rect 27128 5958 27140 6010
rect 27192 5958 27204 6010
rect 27256 5958 30820 6010
rect 1104 5936 30820 5958
rect 1104 5466 30820 5488
rect 1104 5414 5324 5466
rect 5376 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 12752 5466
rect 12804 5414 12816 5466
rect 12868 5414 12880 5466
rect 12932 5414 12944 5466
rect 12996 5414 13008 5466
rect 13060 5414 20180 5466
rect 20232 5414 20244 5466
rect 20296 5414 20308 5466
rect 20360 5414 20372 5466
rect 20424 5414 20436 5466
rect 20488 5414 27608 5466
rect 27660 5414 27672 5466
rect 27724 5414 27736 5466
rect 27788 5414 27800 5466
rect 27852 5414 27864 5466
rect 27916 5414 30820 5466
rect 1104 5392 30820 5414
rect 1104 4922 30820 4944
rect 1104 4870 4664 4922
rect 4716 4870 4728 4922
rect 4780 4870 4792 4922
rect 4844 4870 4856 4922
rect 4908 4870 4920 4922
rect 4972 4870 12092 4922
rect 12144 4870 12156 4922
rect 12208 4870 12220 4922
rect 12272 4870 12284 4922
rect 12336 4870 12348 4922
rect 12400 4870 19520 4922
rect 19572 4870 19584 4922
rect 19636 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 26948 4922
rect 27000 4870 27012 4922
rect 27064 4870 27076 4922
rect 27128 4870 27140 4922
rect 27192 4870 27204 4922
rect 27256 4870 30820 4922
rect 1104 4848 30820 4870
rect 1104 4378 30820 4400
rect 1104 4326 5324 4378
rect 5376 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 12752 4378
rect 12804 4326 12816 4378
rect 12868 4326 12880 4378
rect 12932 4326 12944 4378
rect 12996 4326 13008 4378
rect 13060 4326 20180 4378
rect 20232 4326 20244 4378
rect 20296 4326 20308 4378
rect 20360 4326 20372 4378
rect 20424 4326 20436 4378
rect 20488 4326 27608 4378
rect 27660 4326 27672 4378
rect 27724 4326 27736 4378
rect 27788 4326 27800 4378
rect 27852 4326 27864 4378
rect 27916 4326 30820 4378
rect 1104 4304 30820 4326
rect 1104 3834 30820 3856
rect 1104 3782 4664 3834
rect 4716 3782 4728 3834
rect 4780 3782 4792 3834
rect 4844 3782 4856 3834
rect 4908 3782 4920 3834
rect 4972 3782 12092 3834
rect 12144 3782 12156 3834
rect 12208 3782 12220 3834
rect 12272 3782 12284 3834
rect 12336 3782 12348 3834
rect 12400 3782 19520 3834
rect 19572 3782 19584 3834
rect 19636 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 26948 3834
rect 27000 3782 27012 3834
rect 27064 3782 27076 3834
rect 27128 3782 27140 3834
rect 27192 3782 27204 3834
rect 27256 3782 30820 3834
rect 1104 3760 30820 3782
rect 1104 3290 30820 3312
rect 1104 3238 5324 3290
rect 5376 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 12752 3290
rect 12804 3238 12816 3290
rect 12868 3238 12880 3290
rect 12932 3238 12944 3290
rect 12996 3238 13008 3290
rect 13060 3238 20180 3290
rect 20232 3238 20244 3290
rect 20296 3238 20308 3290
rect 20360 3238 20372 3290
rect 20424 3238 20436 3290
rect 20488 3238 27608 3290
rect 27660 3238 27672 3290
rect 27724 3238 27736 3290
rect 27788 3238 27800 3290
rect 27852 3238 27864 3290
rect 27916 3238 30820 3290
rect 1104 3216 30820 3238
rect 1104 2746 30820 2768
rect 1104 2694 4664 2746
rect 4716 2694 4728 2746
rect 4780 2694 4792 2746
rect 4844 2694 4856 2746
rect 4908 2694 4920 2746
rect 4972 2694 12092 2746
rect 12144 2694 12156 2746
rect 12208 2694 12220 2746
rect 12272 2694 12284 2746
rect 12336 2694 12348 2746
rect 12400 2694 19520 2746
rect 19572 2694 19584 2746
rect 19636 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 26948 2746
rect 27000 2694 27012 2746
rect 27064 2694 27076 2746
rect 27128 2694 27140 2746
rect 27192 2694 27204 2746
rect 27256 2694 30820 2746
rect 1104 2672 30820 2694
rect 9306 2592 9312 2644
rect 9364 2592 9370 2644
rect 9950 2592 9956 2644
rect 10008 2592 10014 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11112 2604 11897 2632
rect 11112 2592 11118 2604
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 13817 2635 13875 2641
rect 13817 2601 13829 2635
rect 13863 2632 13875 2635
rect 13998 2632 14004 2644
rect 13863 2604 14004 2632
rect 13863 2601 13875 2604
rect 13817 2595 13875 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16114 2592 16120 2644
rect 16172 2592 16178 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17126 2632 17132 2644
rect 17083 2604 17132 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 17862 2632 17868 2644
rect 17727 2604 17868 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18966 2592 18972 2644
rect 19024 2592 19030 2644
rect 21450 2592 21456 2644
rect 21508 2632 21514 2644
rect 21545 2635 21603 2641
rect 21545 2632 21557 2635
rect 21508 2604 21557 2632
rect 21508 2592 21514 2604
rect 21545 2601 21557 2604
rect 21591 2601 21603 2635
rect 21545 2595 21603 2601
rect 15197 2567 15255 2573
rect 15197 2533 15209 2567
rect 15243 2564 15255 2567
rect 16132 2564 16160 2592
rect 15243 2536 16160 2564
rect 15243 2533 15255 2536
rect 15197 2527 15255 2533
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 15838 2388 15844 2440
rect 15896 2388 15902 2440
rect 16482 2388 16488 2440
rect 16540 2388 16546 2440
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 20990 2388 20996 2440
rect 21048 2388 21054 2440
rect 21358 2388 21364 2440
rect 21416 2388 21422 2440
rect 15010 2320 15016 2372
rect 15068 2320 15074 2372
rect 16942 2320 16948 2372
rect 17000 2320 17006 2372
rect 17586 2320 17592 2372
rect 17644 2320 17650 2372
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12308 2264 12449 2292
rect 12308 2252 12314 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 15654 2252 15660 2304
rect 15712 2252 15718 2304
rect 16298 2252 16304 2304
rect 16356 2252 16362 2304
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20680 2264 20821 2292
rect 20680 2252 20686 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 1104 2202 30820 2224
rect 1104 2150 5324 2202
rect 5376 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 12752 2202
rect 12804 2150 12816 2202
rect 12868 2150 12880 2202
rect 12932 2150 12944 2202
rect 12996 2150 13008 2202
rect 13060 2150 20180 2202
rect 20232 2150 20244 2202
rect 20296 2150 20308 2202
rect 20360 2150 20372 2202
rect 20424 2150 20436 2202
rect 20488 2150 27608 2202
rect 27660 2150 27672 2202
rect 27724 2150 27736 2202
rect 27788 2150 27800 2202
rect 27852 2150 27864 2202
rect 27916 2150 30820 2202
rect 1104 2128 30820 2150
<< via1 >>
rect 5324 29350 5376 29402
rect 5388 29350 5440 29402
rect 5452 29350 5504 29402
rect 5516 29350 5568 29402
rect 5580 29350 5632 29402
rect 12752 29350 12804 29402
rect 12816 29350 12868 29402
rect 12880 29350 12932 29402
rect 12944 29350 12996 29402
rect 13008 29350 13060 29402
rect 20180 29350 20232 29402
rect 20244 29350 20296 29402
rect 20308 29350 20360 29402
rect 20372 29350 20424 29402
rect 20436 29350 20488 29402
rect 27608 29350 27660 29402
rect 27672 29350 27724 29402
rect 27736 29350 27788 29402
rect 27800 29350 27852 29402
rect 27864 29350 27916 29402
rect 12348 29248 12400 29300
rect 13084 29248 13136 29300
rect 14280 29248 14332 29300
rect 15752 29291 15804 29300
rect 15752 29257 15761 29291
rect 15761 29257 15795 29291
rect 15795 29257 15804 29291
rect 15752 29248 15804 29257
rect 18696 29248 18748 29300
rect 19616 29248 19668 29300
rect 20628 29248 20680 29300
rect 21916 29248 21968 29300
rect 14832 29180 14884 29232
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 15660 29155 15712 29164
rect 15660 29121 15669 29155
rect 15669 29121 15703 29155
rect 15703 29121 15712 29155
rect 15660 29112 15712 29121
rect 19340 29155 19392 29164
rect 19340 29121 19349 29155
rect 19349 29121 19383 29155
rect 19383 29121 19392 29155
rect 19340 29112 19392 29121
rect 19892 29155 19944 29164
rect 19892 29121 19901 29155
rect 19901 29121 19935 29155
rect 19935 29121 19944 29155
rect 19892 29112 19944 29121
rect 20812 29155 20864 29164
rect 20812 29121 20821 29155
rect 20821 29121 20855 29155
rect 20855 29121 20864 29155
rect 20812 29112 20864 29121
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 22100 29112 22152 29121
rect 13268 29044 13320 29096
rect 12532 28976 12584 29028
rect 15200 29019 15252 29028
rect 15200 28985 15209 29019
rect 15209 28985 15243 29019
rect 15243 28985 15252 29019
rect 15200 28976 15252 28985
rect 4664 28806 4716 28858
rect 4728 28806 4780 28858
rect 4792 28806 4844 28858
rect 4856 28806 4908 28858
rect 4920 28806 4972 28858
rect 12092 28806 12144 28858
rect 12156 28806 12208 28858
rect 12220 28806 12272 28858
rect 12284 28806 12336 28858
rect 12348 28806 12400 28858
rect 19520 28806 19572 28858
rect 19584 28806 19636 28858
rect 19648 28806 19700 28858
rect 19712 28806 19764 28858
rect 19776 28806 19828 28858
rect 26948 28806 27000 28858
rect 27012 28806 27064 28858
rect 27076 28806 27128 28858
rect 27140 28806 27192 28858
rect 27204 28806 27256 28858
rect 5324 28262 5376 28314
rect 5388 28262 5440 28314
rect 5452 28262 5504 28314
rect 5516 28262 5568 28314
rect 5580 28262 5632 28314
rect 12752 28262 12804 28314
rect 12816 28262 12868 28314
rect 12880 28262 12932 28314
rect 12944 28262 12996 28314
rect 13008 28262 13060 28314
rect 20180 28262 20232 28314
rect 20244 28262 20296 28314
rect 20308 28262 20360 28314
rect 20372 28262 20424 28314
rect 20436 28262 20488 28314
rect 27608 28262 27660 28314
rect 27672 28262 27724 28314
rect 27736 28262 27788 28314
rect 27800 28262 27852 28314
rect 27864 28262 27916 28314
rect 4664 27718 4716 27770
rect 4728 27718 4780 27770
rect 4792 27718 4844 27770
rect 4856 27718 4908 27770
rect 4920 27718 4972 27770
rect 12092 27718 12144 27770
rect 12156 27718 12208 27770
rect 12220 27718 12272 27770
rect 12284 27718 12336 27770
rect 12348 27718 12400 27770
rect 19520 27718 19572 27770
rect 19584 27718 19636 27770
rect 19648 27718 19700 27770
rect 19712 27718 19764 27770
rect 19776 27718 19828 27770
rect 26948 27718 27000 27770
rect 27012 27718 27064 27770
rect 27076 27718 27128 27770
rect 27140 27718 27192 27770
rect 27204 27718 27256 27770
rect 5324 27174 5376 27226
rect 5388 27174 5440 27226
rect 5452 27174 5504 27226
rect 5516 27174 5568 27226
rect 5580 27174 5632 27226
rect 12752 27174 12804 27226
rect 12816 27174 12868 27226
rect 12880 27174 12932 27226
rect 12944 27174 12996 27226
rect 13008 27174 13060 27226
rect 20180 27174 20232 27226
rect 20244 27174 20296 27226
rect 20308 27174 20360 27226
rect 20372 27174 20424 27226
rect 20436 27174 20488 27226
rect 27608 27174 27660 27226
rect 27672 27174 27724 27226
rect 27736 27174 27788 27226
rect 27800 27174 27852 27226
rect 27864 27174 27916 27226
rect 4664 26630 4716 26682
rect 4728 26630 4780 26682
rect 4792 26630 4844 26682
rect 4856 26630 4908 26682
rect 4920 26630 4972 26682
rect 12092 26630 12144 26682
rect 12156 26630 12208 26682
rect 12220 26630 12272 26682
rect 12284 26630 12336 26682
rect 12348 26630 12400 26682
rect 19520 26630 19572 26682
rect 19584 26630 19636 26682
rect 19648 26630 19700 26682
rect 19712 26630 19764 26682
rect 19776 26630 19828 26682
rect 26948 26630 27000 26682
rect 27012 26630 27064 26682
rect 27076 26630 27128 26682
rect 27140 26630 27192 26682
rect 27204 26630 27256 26682
rect 5324 26086 5376 26138
rect 5388 26086 5440 26138
rect 5452 26086 5504 26138
rect 5516 26086 5568 26138
rect 5580 26086 5632 26138
rect 12752 26086 12804 26138
rect 12816 26086 12868 26138
rect 12880 26086 12932 26138
rect 12944 26086 12996 26138
rect 13008 26086 13060 26138
rect 20180 26086 20232 26138
rect 20244 26086 20296 26138
rect 20308 26086 20360 26138
rect 20372 26086 20424 26138
rect 20436 26086 20488 26138
rect 27608 26086 27660 26138
rect 27672 26086 27724 26138
rect 27736 26086 27788 26138
rect 27800 26086 27852 26138
rect 27864 26086 27916 26138
rect 20076 25848 20128 25900
rect 22744 25848 22796 25900
rect 21180 25644 21232 25696
rect 4664 25542 4716 25594
rect 4728 25542 4780 25594
rect 4792 25542 4844 25594
rect 4856 25542 4908 25594
rect 4920 25542 4972 25594
rect 12092 25542 12144 25594
rect 12156 25542 12208 25594
rect 12220 25542 12272 25594
rect 12284 25542 12336 25594
rect 12348 25542 12400 25594
rect 19520 25542 19572 25594
rect 19584 25542 19636 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 26948 25542 27000 25594
rect 27012 25542 27064 25594
rect 27076 25542 27128 25594
rect 27140 25542 27192 25594
rect 27204 25542 27256 25594
rect 18972 25440 19024 25492
rect 14740 25304 14792 25356
rect 18420 25304 18472 25356
rect 14924 25236 14976 25288
rect 14832 25168 14884 25220
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 16212 25211 16264 25220
rect 16212 25177 16221 25211
rect 16221 25177 16255 25211
rect 16255 25177 16264 25211
rect 16212 25168 16264 25177
rect 17224 25168 17276 25220
rect 17868 25168 17920 25220
rect 20076 25236 20128 25288
rect 24216 25304 24268 25356
rect 20536 25168 20588 25220
rect 21180 25168 21232 25220
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 16028 25100 16080 25152
rect 18144 25100 18196 25152
rect 18788 25100 18840 25152
rect 19432 25143 19484 25152
rect 19432 25109 19441 25143
rect 19441 25109 19475 25143
rect 19475 25109 19484 25143
rect 19432 25100 19484 25109
rect 21364 25100 21416 25152
rect 22836 25168 22888 25220
rect 22284 25100 22336 25152
rect 22560 25100 22612 25152
rect 24676 25211 24728 25220
rect 24676 25177 24685 25211
rect 24685 25177 24719 25211
rect 24719 25177 24728 25211
rect 24676 25168 24728 25177
rect 25228 25168 25280 25220
rect 24860 25100 24912 25152
rect 5324 24998 5376 25050
rect 5388 24998 5440 25050
rect 5452 24998 5504 25050
rect 5516 24998 5568 25050
rect 5580 24998 5632 25050
rect 12752 24998 12804 25050
rect 12816 24998 12868 25050
rect 12880 24998 12932 25050
rect 12944 24998 12996 25050
rect 13008 24998 13060 25050
rect 20180 24998 20232 25050
rect 20244 24998 20296 25050
rect 20308 24998 20360 25050
rect 20372 24998 20424 25050
rect 20436 24998 20488 25050
rect 27608 24998 27660 25050
rect 27672 24998 27724 25050
rect 27736 24998 27788 25050
rect 27800 24998 27852 25050
rect 27864 24998 27916 25050
rect 17224 24939 17276 24948
rect 17224 24905 17233 24939
rect 17233 24905 17267 24939
rect 17267 24905 17276 24939
rect 17224 24896 17276 24905
rect 20536 24896 20588 24948
rect 22560 24896 22612 24948
rect 22836 24896 22888 24948
rect 24676 24896 24728 24948
rect 25228 24939 25280 24948
rect 25228 24905 25237 24939
rect 25237 24905 25271 24939
rect 25271 24905 25280 24939
rect 25228 24896 25280 24905
rect 14740 24871 14792 24880
rect 14740 24837 14749 24871
rect 14749 24837 14783 24871
rect 14783 24837 14792 24871
rect 14740 24828 14792 24837
rect 15752 24828 15804 24880
rect 19432 24828 19484 24880
rect 14188 24760 14240 24812
rect 16028 24760 16080 24812
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 18328 24803 18380 24812
rect 18328 24769 18337 24803
rect 18337 24769 18371 24803
rect 18371 24769 18380 24803
rect 18328 24760 18380 24769
rect 12624 24735 12676 24744
rect 12624 24701 12633 24735
rect 12633 24701 12667 24735
rect 12667 24701 12676 24735
rect 12624 24692 12676 24701
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 14464 24735 14516 24744
rect 14464 24701 14473 24735
rect 14473 24701 14507 24735
rect 14507 24701 14516 24735
rect 14464 24692 14516 24701
rect 15936 24692 15988 24744
rect 14556 24556 14608 24608
rect 16120 24692 16172 24744
rect 17960 24599 18012 24608
rect 17960 24565 17969 24599
rect 17969 24565 18003 24599
rect 18003 24565 18012 24599
rect 17960 24556 18012 24565
rect 18420 24735 18472 24744
rect 18420 24701 18429 24735
rect 18429 24701 18463 24735
rect 18463 24701 18472 24735
rect 18420 24692 18472 24701
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 20628 24803 20680 24812
rect 20628 24769 20637 24803
rect 20637 24769 20671 24803
rect 20671 24769 20680 24803
rect 20628 24760 20680 24769
rect 20720 24692 20772 24744
rect 21364 24760 21416 24812
rect 21824 24760 21876 24812
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22836 24803 22888 24812
rect 22836 24769 22845 24803
rect 22845 24769 22879 24803
rect 22879 24769 22888 24803
rect 22836 24760 22888 24769
rect 23204 24692 23256 24744
rect 23756 24692 23808 24744
rect 24124 24803 24176 24812
rect 24124 24769 24133 24803
rect 24133 24769 24167 24803
rect 24167 24769 24176 24803
rect 24124 24760 24176 24769
rect 19984 24556 20036 24608
rect 20444 24556 20496 24608
rect 21916 24556 21968 24608
rect 22284 24556 22336 24608
rect 23204 24556 23256 24608
rect 23296 24556 23348 24608
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 25964 24760 26016 24812
rect 25596 24556 25648 24608
rect 4664 24454 4716 24506
rect 4728 24454 4780 24506
rect 4792 24454 4844 24506
rect 4856 24454 4908 24506
rect 4920 24454 4972 24506
rect 12092 24454 12144 24506
rect 12156 24454 12208 24506
rect 12220 24454 12272 24506
rect 12284 24454 12336 24506
rect 12348 24454 12400 24506
rect 19520 24454 19572 24506
rect 19584 24454 19636 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 26948 24454 27000 24506
rect 27012 24454 27064 24506
rect 27076 24454 27128 24506
rect 27140 24454 27192 24506
rect 27204 24454 27256 24506
rect 12624 24352 12676 24404
rect 14188 24395 14240 24404
rect 14188 24361 14197 24395
rect 14197 24361 14231 24395
rect 14231 24361 14240 24395
rect 14188 24352 14240 24361
rect 14464 24352 14516 24404
rect 16212 24352 16264 24404
rect 13084 24148 13136 24200
rect 17960 24352 18012 24404
rect 18696 24352 18748 24404
rect 20076 24352 20128 24404
rect 20628 24352 20680 24404
rect 14372 24148 14424 24200
rect 14832 24191 14884 24200
rect 14832 24157 14841 24191
rect 14841 24157 14875 24191
rect 14875 24157 14884 24191
rect 14832 24148 14884 24157
rect 14924 24191 14976 24200
rect 14924 24157 14933 24191
rect 14933 24157 14967 24191
rect 14967 24157 14976 24191
rect 14924 24148 14976 24157
rect 14556 24080 14608 24132
rect 14280 24012 14332 24064
rect 15384 24080 15436 24132
rect 17224 24148 17276 24200
rect 17500 24216 17552 24268
rect 17868 24216 17920 24268
rect 18604 24284 18656 24336
rect 20444 24284 20496 24336
rect 16120 24080 16172 24132
rect 16948 24012 17000 24064
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 18144 24080 18196 24132
rect 18788 24123 18840 24132
rect 18788 24089 18797 24123
rect 18797 24089 18831 24123
rect 18831 24089 18840 24123
rect 20628 24216 20680 24268
rect 21824 24395 21876 24404
rect 21824 24361 21833 24395
rect 21833 24361 21867 24395
rect 21867 24361 21876 24395
rect 21824 24352 21876 24361
rect 21916 24352 21968 24404
rect 22376 24352 22428 24404
rect 22836 24352 22888 24404
rect 19984 24148 20036 24200
rect 20904 24259 20956 24268
rect 20904 24225 20914 24259
rect 20914 24225 20948 24259
rect 20948 24225 20956 24259
rect 20904 24216 20956 24225
rect 21088 24216 21140 24268
rect 18788 24080 18840 24089
rect 20720 24080 20772 24132
rect 21732 24191 21784 24200
rect 21732 24157 21741 24191
rect 21741 24157 21775 24191
rect 21775 24157 21784 24191
rect 21732 24148 21784 24157
rect 22284 24148 22336 24200
rect 23664 24284 23716 24336
rect 25136 24284 25188 24336
rect 25504 24216 25556 24268
rect 21272 24080 21324 24132
rect 21364 24123 21416 24132
rect 21364 24089 21373 24123
rect 21373 24089 21407 24123
rect 21407 24089 21416 24123
rect 21364 24080 21416 24089
rect 21456 24080 21508 24132
rect 23296 24080 23348 24132
rect 24952 24148 25004 24200
rect 17500 24055 17552 24064
rect 17500 24021 17509 24055
rect 17509 24021 17543 24055
rect 17543 24021 17552 24055
rect 17500 24012 17552 24021
rect 20996 24012 21048 24064
rect 23020 24055 23072 24064
rect 23020 24021 23029 24055
rect 23029 24021 23063 24055
rect 23063 24021 23072 24055
rect 23020 24012 23072 24021
rect 23388 24012 23440 24064
rect 23480 24012 23532 24064
rect 24124 24012 24176 24064
rect 24492 24055 24544 24064
rect 24492 24021 24501 24055
rect 24501 24021 24535 24055
rect 24535 24021 24544 24055
rect 24492 24012 24544 24021
rect 24860 24012 24912 24064
rect 26056 24080 26108 24132
rect 25504 24012 25556 24064
rect 5324 23910 5376 23962
rect 5388 23910 5440 23962
rect 5452 23910 5504 23962
rect 5516 23910 5568 23962
rect 5580 23910 5632 23962
rect 12752 23910 12804 23962
rect 12816 23910 12868 23962
rect 12880 23910 12932 23962
rect 12944 23910 12996 23962
rect 13008 23910 13060 23962
rect 20180 23910 20232 23962
rect 20244 23910 20296 23962
rect 20308 23910 20360 23962
rect 20372 23910 20424 23962
rect 20436 23910 20488 23962
rect 27608 23910 27660 23962
rect 27672 23910 27724 23962
rect 27736 23910 27788 23962
rect 27800 23910 27852 23962
rect 27864 23910 27916 23962
rect 13084 23808 13136 23860
rect 15016 23808 15068 23860
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 17224 23808 17276 23860
rect 17500 23808 17552 23860
rect 18144 23851 18196 23860
rect 18144 23817 18153 23851
rect 18153 23817 18187 23851
rect 18187 23817 18196 23851
rect 18144 23808 18196 23817
rect 18604 23808 18656 23860
rect 18880 23808 18932 23860
rect 1492 23715 1544 23724
rect 1492 23681 1501 23715
rect 1501 23681 1535 23715
rect 1535 23681 1544 23715
rect 1492 23672 1544 23681
rect 11980 23740 12032 23792
rect 13912 23740 13964 23792
rect 14648 23740 14700 23792
rect 11796 23715 11848 23724
rect 11796 23681 11830 23715
rect 11830 23681 11848 23715
rect 11796 23672 11848 23681
rect 14372 23672 14424 23724
rect 14832 23715 14884 23724
rect 14832 23681 14841 23715
rect 14841 23681 14875 23715
rect 14875 23681 14884 23715
rect 14832 23672 14884 23681
rect 17960 23715 18012 23724
rect 17960 23681 17969 23715
rect 17969 23681 18003 23715
rect 18003 23681 18012 23715
rect 17960 23672 18012 23681
rect 18512 23715 18564 23724
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 20628 23808 20680 23860
rect 20720 23808 20772 23860
rect 20904 23851 20956 23860
rect 20904 23817 20913 23851
rect 20913 23817 20947 23851
rect 20947 23817 20956 23851
rect 20904 23808 20956 23817
rect 19984 23740 20036 23792
rect 24124 23808 24176 23860
rect 22284 23740 22336 23792
rect 19432 23672 19484 23724
rect 6920 23536 6972 23588
rect 13268 23536 13320 23588
rect 14924 23468 14976 23520
rect 16120 23536 16172 23588
rect 16948 23468 17000 23520
rect 17132 23468 17184 23520
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 18880 23604 18932 23656
rect 20904 23672 20956 23724
rect 20076 23604 20128 23656
rect 21456 23672 21508 23724
rect 23388 23740 23440 23792
rect 23480 23715 23532 23724
rect 23480 23681 23489 23715
rect 23489 23681 23523 23715
rect 23523 23681 23532 23715
rect 23480 23672 23532 23681
rect 23664 23672 23716 23724
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 21180 23536 21232 23588
rect 22192 23579 22244 23588
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 22192 23536 22244 23545
rect 23020 23536 23072 23588
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24032 23647 24084 23656
rect 24032 23613 24041 23647
rect 24041 23613 24075 23647
rect 24075 23613 24084 23647
rect 24032 23604 24084 23613
rect 24124 23647 24176 23656
rect 24124 23613 24133 23647
rect 24133 23613 24167 23647
rect 24167 23613 24176 23647
rect 24124 23604 24176 23613
rect 25504 23808 25556 23860
rect 26056 23851 26108 23860
rect 26056 23817 26065 23851
rect 26065 23817 26099 23851
rect 26099 23817 26108 23851
rect 26056 23808 26108 23817
rect 25964 23715 26016 23724
rect 25964 23681 25973 23715
rect 25973 23681 26007 23715
rect 26007 23681 26016 23715
rect 25964 23672 26016 23681
rect 30288 23672 30340 23724
rect 25412 23647 25464 23656
rect 25412 23613 25421 23647
rect 25421 23613 25455 23647
rect 25455 23613 25464 23647
rect 25412 23604 25464 23613
rect 25596 23647 25648 23656
rect 25596 23613 25605 23647
rect 25605 23613 25639 23647
rect 25639 23613 25648 23647
rect 25596 23604 25648 23613
rect 26056 23536 26108 23588
rect 18604 23468 18656 23520
rect 20352 23468 20404 23520
rect 20904 23468 20956 23520
rect 21364 23468 21416 23520
rect 21548 23468 21600 23520
rect 23480 23468 23532 23520
rect 24124 23468 24176 23520
rect 4664 23366 4716 23418
rect 4728 23366 4780 23418
rect 4792 23366 4844 23418
rect 4856 23366 4908 23418
rect 4920 23366 4972 23418
rect 12092 23366 12144 23418
rect 12156 23366 12208 23418
rect 12220 23366 12272 23418
rect 12284 23366 12336 23418
rect 12348 23366 12400 23418
rect 19520 23366 19572 23418
rect 19584 23366 19636 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 26948 23366 27000 23418
rect 27012 23366 27064 23418
rect 27076 23366 27128 23418
rect 27140 23366 27192 23418
rect 27204 23366 27256 23418
rect 11796 23264 11848 23316
rect 12256 23307 12308 23316
rect 12256 23273 12265 23307
rect 12265 23273 12299 23307
rect 12299 23273 12308 23307
rect 12256 23264 12308 23273
rect 14924 23264 14976 23316
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 14832 23171 14884 23180
rect 14832 23137 14841 23171
rect 14841 23137 14875 23171
rect 14875 23137 14884 23171
rect 14832 23128 14884 23137
rect 16212 23264 16264 23316
rect 16304 23264 16356 23316
rect 17960 23264 18012 23316
rect 22192 23264 22244 23316
rect 23664 23264 23716 23316
rect 23940 23264 23992 23316
rect 25412 23264 25464 23316
rect 16120 23239 16172 23248
rect 16120 23205 16129 23239
rect 16129 23205 16163 23239
rect 16163 23205 16172 23239
rect 16120 23196 16172 23205
rect 11980 23060 12032 23112
rect 17224 23196 17276 23248
rect 19432 23128 19484 23180
rect 20720 23128 20772 23180
rect 22008 23171 22060 23180
rect 22008 23137 22017 23171
rect 22017 23137 22051 23171
rect 22051 23137 22060 23171
rect 22008 23128 22060 23137
rect 9864 22992 9916 23044
rect 12624 22924 12676 22976
rect 15108 22992 15160 23044
rect 15476 22967 15528 22976
rect 15476 22933 15485 22967
rect 15485 22933 15519 22967
rect 15519 22933 15528 22967
rect 15476 22924 15528 22933
rect 15568 22967 15620 22976
rect 15568 22933 15577 22967
rect 15577 22933 15611 22967
rect 15611 22933 15620 22967
rect 15568 22924 15620 22933
rect 17040 23103 17092 23112
rect 17040 23069 17049 23103
rect 17049 23069 17083 23103
rect 17083 23069 17092 23103
rect 17040 23060 17092 23069
rect 20352 23060 20404 23112
rect 20444 23103 20496 23112
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 21180 23060 21232 23112
rect 23388 23196 23440 23248
rect 23480 23060 23532 23112
rect 16304 22924 16356 22976
rect 16488 22924 16540 22976
rect 18972 22992 19024 23044
rect 23848 23103 23900 23112
rect 23848 23069 23857 23103
rect 23857 23069 23891 23103
rect 23891 23069 23900 23103
rect 23848 23060 23900 23069
rect 24492 23060 24544 23112
rect 18696 22924 18748 22976
rect 20536 22924 20588 22976
rect 21088 22924 21140 22976
rect 22284 22924 22336 22976
rect 25872 23060 25924 23112
rect 24860 23035 24912 23044
rect 24860 23001 24869 23035
rect 24869 23001 24903 23035
rect 24903 23001 24912 23035
rect 24860 22992 24912 23001
rect 24952 23035 25004 23044
rect 24952 23001 24961 23035
rect 24961 23001 24995 23035
rect 24995 23001 25004 23035
rect 24952 22992 25004 23001
rect 25596 22924 25648 22976
rect 5324 22822 5376 22874
rect 5388 22822 5440 22874
rect 5452 22822 5504 22874
rect 5516 22822 5568 22874
rect 5580 22822 5632 22874
rect 12752 22822 12804 22874
rect 12816 22822 12868 22874
rect 12880 22822 12932 22874
rect 12944 22822 12996 22874
rect 13008 22822 13060 22874
rect 20180 22822 20232 22874
rect 20244 22822 20296 22874
rect 20308 22822 20360 22874
rect 20372 22822 20424 22874
rect 20436 22822 20488 22874
rect 27608 22822 27660 22874
rect 27672 22822 27724 22874
rect 27736 22822 27788 22874
rect 27800 22822 27852 22874
rect 27864 22822 27916 22874
rect 12624 22720 12676 22772
rect 14832 22720 14884 22772
rect 18328 22720 18380 22772
rect 12256 22695 12308 22704
rect 12256 22661 12265 22695
rect 12265 22661 12299 22695
rect 12299 22661 12308 22695
rect 12256 22652 12308 22661
rect 4436 22584 4488 22636
rect 940 22448 992 22500
rect 6092 22584 6144 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 7656 22584 7708 22636
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 8300 22559 8352 22568
rect 8300 22525 8309 22559
rect 8309 22525 8343 22559
rect 8343 22525 8352 22559
rect 8300 22516 8352 22525
rect 9956 22559 10008 22568
rect 9956 22525 9965 22559
rect 9965 22525 9999 22559
rect 9999 22525 10008 22559
rect 9956 22516 10008 22525
rect 11612 22559 11664 22568
rect 11612 22525 11621 22559
rect 11621 22525 11655 22559
rect 11655 22525 11664 22559
rect 11612 22516 11664 22525
rect 13820 22559 13872 22568
rect 13820 22525 13829 22559
rect 13829 22525 13863 22559
rect 13863 22525 13872 22559
rect 13820 22516 13872 22525
rect 14924 22516 14976 22568
rect 5080 22380 5132 22432
rect 5356 22380 5408 22432
rect 7012 22423 7064 22432
rect 7012 22389 7021 22423
rect 7021 22389 7055 22423
rect 7055 22389 7064 22423
rect 7012 22380 7064 22389
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 9864 22380 9916 22432
rect 18788 22720 18840 22772
rect 20536 22720 20588 22772
rect 18972 22652 19024 22704
rect 21272 22720 21324 22772
rect 21732 22720 21784 22772
rect 22560 22720 22612 22772
rect 18604 22516 18656 22568
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 21088 22652 21140 22704
rect 23204 22652 23256 22704
rect 24032 22652 24084 22704
rect 25872 22763 25924 22772
rect 25872 22729 25881 22763
rect 25881 22729 25915 22763
rect 25915 22729 25924 22763
rect 25872 22720 25924 22729
rect 20996 22627 21048 22636
rect 20996 22593 21010 22627
rect 21010 22593 21044 22627
rect 21044 22593 21048 22627
rect 20996 22584 21048 22593
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 20904 22516 20956 22568
rect 12808 22380 12860 22432
rect 14556 22380 14608 22432
rect 15016 22423 15068 22432
rect 15016 22389 15025 22423
rect 15025 22389 15059 22423
rect 15059 22389 15068 22423
rect 15016 22380 15068 22389
rect 15568 22380 15620 22432
rect 16120 22380 16172 22432
rect 17040 22380 17092 22432
rect 17592 22380 17644 22432
rect 19064 22448 19116 22500
rect 22284 22627 22336 22636
rect 22284 22593 22293 22627
rect 22293 22593 22327 22627
rect 22327 22593 22336 22627
rect 22284 22584 22336 22593
rect 21456 22559 21508 22568
rect 21456 22525 21465 22559
rect 21465 22525 21499 22559
rect 21499 22525 21508 22559
rect 21456 22516 21508 22525
rect 22008 22516 22060 22568
rect 22192 22448 22244 22500
rect 20076 22380 20128 22432
rect 20904 22380 20956 22432
rect 22560 22627 22612 22636
rect 22560 22593 22595 22627
rect 22595 22593 22612 22627
rect 22560 22584 22612 22593
rect 22744 22559 22796 22568
rect 22744 22525 22753 22559
rect 22753 22525 22787 22559
rect 22787 22525 22796 22559
rect 22744 22516 22796 22525
rect 23388 22584 23440 22636
rect 25596 22584 25648 22636
rect 26056 22584 26108 22636
rect 26240 22627 26292 22636
rect 26240 22593 26249 22627
rect 26249 22593 26283 22627
rect 26283 22593 26292 22627
rect 26240 22584 26292 22593
rect 30932 22584 30984 22636
rect 24860 22516 24912 22568
rect 25504 22559 25556 22568
rect 25504 22525 25513 22559
rect 25513 22525 25547 22559
rect 25547 22525 25556 22559
rect 25504 22516 25556 22525
rect 23204 22448 23256 22500
rect 24032 22380 24084 22432
rect 24952 22380 25004 22432
rect 4664 22278 4716 22330
rect 4728 22278 4780 22330
rect 4792 22278 4844 22330
rect 4856 22278 4908 22330
rect 4920 22278 4972 22330
rect 12092 22278 12144 22330
rect 12156 22278 12208 22330
rect 12220 22278 12272 22330
rect 12284 22278 12336 22330
rect 12348 22278 12400 22330
rect 19520 22278 19572 22330
rect 19584 22278 19636 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 26948 22278 27000 22330
rect 27012 22278 27064 22330
rect 27076 22278 27128 22330
rect 27140 22278 27192 22330
rect 27204 22278 27256 22330
rect 5172 22219 5224 22228
rect 5172 22185 5181 22219
rect 5181 22185 5215 22219
rect 5215 22185 5224 22219
rect 5172 22176 5224 22185
rect 5724 22176 5776 22228
rect 6736 22176 6788 22228
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 3792 22015 3844 22024
rect 3792 21981 3801 22015
rect 3801 21981 3835 22015
rect 3835 21981 3844 22015
rect 5816 22015 5868 22024
rect 3792 21972 3844 21981
rect 5816 21981 5825 22015
rect 5825 21981 5859 22015
rect 5859 21981 5868 22015
rect 5816 21972 5868 21981
rect 9404 22176 9456 22228
rect 11612 22219 11664 22228
rect 11612 22185 11621 22219
rect 11621 22185 11655 22219
rect 11655 22185 11664 22219
rect 11612 22176 11664 22185
rect 12808 22176 12860 22228
rect 7656 22083 7708 22092
rect 7656 22049 7665 22083
rect 7665 22049 7699 22083
rect 7699 22049 7708 22083
rect 7656 22040 7708 22049
rect 11980 22040 12032 22092
rect 15292 22108 15344 22160
rect 15384 22108 15436 22160
rect 8760 22015 8812 22024
rect 8760 21981 8769 22015
rect 8769 21981 8803 22015
rect 8803 21981 8812 22015
rect 8760 21972 8812 21981
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 9772 21972 9824 22024
rect 9956 21972 10008 22024
rect 10048 21972 10100 22024
rect 14004 21972 14056 22024
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 4620 21904 4672 21956
rect 5356 21904 5408 21956
rect 940 21836 992 21888
rect 5172 21836 5224 21888
rect 6368 21904 6420 21956
rect 10324 21904 10376 21956
rect 7288 21879 7340 21888
rect 7288 21845 7297 21879
rect 7297 21845 7331 21879
rect 7331 21845 7340 21879
rect 7288 21836 7340 21845
rect 8300 21836 8352 21888
rect 8484 21836 8536 21888
rect 9956 21836 10008 21888
rect 13912 21879 13964 21888
rect 13912 21845 13921 21879
rect 13921 21845 13955 21879
rect 13955 21845 13964 21879
rect 13912 21836 13964 21845
rect 14372 21836 14424 21888
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15292 21836 15344 21888
rect 16488 22176 16540 22228
rect 16856 22176 16908 22228
rect 17316 22108 17368 22160
rect 16120 21947 16172 21956
rect 16120 21913 16129 21947
rect 16129 21913 16163 21947
rect 16163 21913 16172 21947
rect 16120 21904 16172 21913
rect 16304 21972 16356 22024
rect 17040 22040 17092 22092
rect 17592 22176 17644 22228
rect 18788 22219 18840 22228
rect 18788 22185 18797 22219
rect 18797 22185 18831 22219
rect 18831 22185 18840 22219
rect 18788 22176 18840 22185
rect 19064 22108 19116 22160
rect 20536 22176 20588 22228
rect 21456 22176 21508 22228
rect 22284 22176 22336 22228
rect 23756 22176 23808 22228
rect 23848 22176 23900 22228
rect 16580 21972 16632 22024
rect 15568 21836 15620 21888
rect 15752 21836 15804 21888
rect 16672 21904 16724 21956
rect 18420 22040 18472 22092
rect 18696 22040 18748 22092
rect 19156 22040 19208 22092
rect 19800 22040 19852 22092
rect 23204 22040 23256 22092
rect 18236 21972 18288 22024
rect 18880 21972 18932 22024
rect 20076 22015 20128 22024
rect 20076 21981 20085 22015
rect 20085 21981 20119 22015
rect 20119 21981 20128 22015
rect 20076 21972 20128 21981
rect 20168 21972 20220 22024
rect 20536 21972 20588 22024
rect 21180 21972 21232 22024
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 16856 21836 16908 21888
rect 18052 21836 18104 21888
rect 18420 21947 18472 21956
rect 18420 21913 18429 21947
rect 18429 21913 18463 21947
rect 18463 21913 18472 21947
rect 18420 21904 18472 21913
rect 20720 21904 20772 21956
rect 20904 21904 20956 21956
rect 22100 21972 22152 22024
rect 23388 21972 23440 22024
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 24032 21972 24084 22024
rect 24124 22015 24176 22024
rect 24124 21981 24133 22015
rect 24133 21981 24167 22015
rect 24167 21981 24176 22015
rect 24124 21972 24176 21981
rect 20996 21836 21048 21888
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 24860 21972 24912 22024
rect 25044 21972 25096 22024
rect 24584 21947 24636 21956
rect 24584 21913 24593 21947
rect 24593 21913 24627 21947
rect 24627 21913 24636 21947
rect 24584 21904 24636 21913
rect 26608 21904 26660 21956
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 5324 21734 5376 21786
rect 5388 21734 5440 21786
rect 5452 21734 5504 21786
rect 5516 21734 5568 21786
rect 5580 21734 5632 21786
rect 12752 21734 12804 21786
rect 12816 21734 12868 21786
rect 12880 21734 12932 21786
rect 12944 21734 12996 21786
rect 13008 21734 13060 21786
rect 20180 21734 20232 21786
rect 20244 21734 20296 21786
rect 20308 21734 20360 21786
rect 20372 21734 20424 21786
rect 20436 21734 20488 21786
rect 27608 21734 27660 21786
rect 27672 21734 27724 21786
rect 27736 21734 27788 21786
rect 27800 21734 27852 21786
rect 27864 21734 27916 21786
rect 4620 21675 4672 21684
rect 4620 21641 4629 21675
rect 4629 21641 4663 21675
rect 4663 21641 4672 21675
rect 4620 21632 4672 21641
rect 6368 21675 6420 21684
rect 6368 21641 6377 21675
rect 6377 21641 6411 21675
rect 6411 21641 6420 21675
rect 6368 21632 6420 21641
rect 5080 21496 5132 21548
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 7288 21632 7340 21684
rect 9772 21632 9824 21684
rect 10324 21632 10376 21684
rect 13820 21632 13872 21684
rect 14832 21632 14884 21684
rect 15200 21675 15252 21684
rect 15200 21641 15227 21675
rect 15227 21641 15252 21675
rect 15200 21632 15252 21641
rect 5816 21428 5868 21480
rect 7012 21539 7064 21548
rect 7012 21505 7046 21539
rect 7046 21505 7064 21539
rect 7012 21496 7064 21505
rect 10048 21564 10100 21616
rect 12440 21564 12492 21616
rect 8300 21496 8352 21548
rect 8484 21539 8536 21548
rect 8484 21505 8518 21539
rect 8518 21505 8536 21539
rect 8484 21496 8536 21505
rect 9864 21539 9916 21548
rect 9864 21505 9873 21539
rect 9873 21505 9907 21539
rect 9907 21505 9916 21539
rect 9864 21496 9916 21505
rect 9956 21496 10008 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 14372 21496 14424 21548
rect 15016 21564 15068 21616
rect 15660 21675 15712 21684
rect 15660 21641 15669 21675
rect 15669 21641 15703 21675
rect 15703 21641 15712 21675
rect 15660 21632 15712 21641
rect 19892 21632 19944 21684
rect 19984 21675 20036 21684
rect 19984 21641 19993 21675
rect 19993 21641 20027 21675
rect 20027 21641 20036 21675
rect 19984 21632 20036 21641
rect 20168 21632 20220 21684
rect 16120 21564 16172 21616
rect 17316 21564 17368 21616
rect 11888 21428 11940 21480
rect 13544 21471 13596 21480
rect 13544 21437 13553 21471
rect 13553 21437 13587 21471
rect 13587 21437 13596 21471
rect 13544 21428 13596 21437
rect 6644 21360 6696 21412
rect 14004 21471 14056 21480
rect 14004 21437 14013 21471
rect 14013 21437 14047 21471
rect 14047 21437 14056 21471
rect 14004 21428 14056 21437
rect 15292 21496 15344 21548
rect 15384 21428 15436 21480
rect 15752 21428 15804 21480
rect 16212 21428 16264 21480
rect 16488 21428 16540 21480
rect 15660 21360 15712 21412
rect 16304 21360 16356 21412
rect 940 21292 992 21344
rect 1676 21292 1728 21344
rect 6920 21292 6972 21344
rect 8944 21292 8996 21344
rect 15568 21292 15620 21344
rect 18788 21607 18840 21616
rect 18788 21573 18797 21607
rect 18797 21573 18831 21607
rect 18831 21573 18840 21607
rect 18788 21564 18840 21573
rect 20996 21675 21048 21684
rect 20996 21641 21005 21675
rect 21005 21641 21039 21675
rect 21039 21641 21048 21675
rect 20996 21632 21048 21641
rect 21088 21632 21140 21684
rect 21272 21632 21324 21684
rect 19156 21496 19208 21548
rect 19892 21496 19944 21548
rect 20352 21496 20404 21548
rect 20536 21496 20588 21548
rect 20996 21496 21048 21548
rect 21548 21564 21600 21616
rect 22376 21607 22428 21616
rect 18696 21292 18748 21344
rect 19984 21428 20036 21480
rect 22376 21573 22385 21607
rect 22385 21573 22419 21607
rect 22419 21573 22428 21607
rect 22376 21564 22428 21573
rect 23388 21632 23440 21684
rect 23480 21564 23532 21616
rect 24584 21632 24636 21684
rect 25044 21675 25096 21684
rect 25044 21641 25053 21675
rect 25053 21641 25087 21675
rect 25087 21641 25096 21675
rect 25044 21632 25096 21641
rect 26240 21632 26292 21684
rect 25320 21564 25372 21616
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 23940 21539 23992 21548
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 24584 21496 24636 21548
rect 24860 21539 24912 21548
rect 24860 21505 24869 21539
rect 24869 21505 24903 21539
rect 24903 21505 24912 21539
rect 24860 21496 24912 21505
rect 19800 21403 19852 21412
rect 19800 21369 19809 21403
rect 19809 21369 19843 21403
rect 19843 21369 19852 21403
rect 19800 21360 19852 21369
rect 19892 21360 19944 21412
rect 21088 21360 21140 21412
rect 26148 21539 26200 21548
rect 26148 21505 26157 21539
rect 26157 21505 26191 21539
rect 26191 21505 26200 21539
rect 26148 21496 26200 21505
rect 30472 21539 30524 21548
rect 30472 21505 30481 21539
rect 30481 21505 30515 21539
rect 30515 21505 30524 21539
rect 30472 21496 30524 21505
rect 26332 21428 26384 21480
rect 26608 21428 26660 21480
rect 22284 21360 22336 21412
rect 26056 21360 26108 21412
rect 20076 21292 20128 21344
rect 22192 21292 22244 21344
rect 24400 21292 24452 21344
rect 26240 21292 26292 21344
rect 4664 21190 4716 21242
rect 4728 21190 4780 21242
rect 4792 21190 4844 21242
rect 4856 21190 4908 21242
rect 4920 21190 4972 21242
rect 12092 21190 12144 21242
rect 12156 21190 12208 21242
rect 12220 21190 12272 21242
rect 12284 21190 12336 21242
rect 12348 21190 12400 21242
rect 19520 21190 19572 21242
rect 19584 21190 19636 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 26948 21190 27000 21242
rect 27012 21190 27064 21242
rect 27076 21190 27128 21242
rect 27140 21190 27192 21242
rect 27204 21190 27256 21242
rect 5172 21088 5224 21140
rect 6092 21131 6144 21140
rect 6092 21097 6101 21131
rect 6101 21097 6135 21131
rect 6135 21097 6144 21131
rect 6092 21088 6144 21097
rect 6644 21088 6696 21140
rect 8944 21088 8996 21140
rect 12440 21088 12492 21140
rect 13544 21088 13596 21140
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 3332 20884 3384 20936
rect 3792 20884 3844 20936
rect 9404 21020 9456 21072
rect 14280 21020 14332 21072
rect 15752 21020 15804 21072
rect 20352 21131 20404 21140
rect 20352 21097 20361 21131
rect 20361 21097 20395 21131
rect 20395 21097 20404 21131
rect 20352 21088 20404 21097
rect 20904 21088 20956 21140
rect 11336 20952 11388 21004
rect 9772 20884 9824 20936
rect 15200 20884 15252 20936
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 18696 20995 18748 21004
rect 18696 20961 18705 20995
rect 18705 20961 18739 20995
rect 18739 20961 18748 20995
rect 22192 21088 22244 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 23848 21088 23900 21140
rect 18696 20952 18748 20961
rect 22376 20995 22428 21004
rect 22376 20961 22385 20995
rect 22385 20961 22419 20995
rect 22419 20961 22428 20995
rect 22376 20952 22428 20961
rect 22744 20952 22796 21004
rect 10232 20816 10284 20868
rect 19432 20884 19484 20936
rect 19892 20884 19944 20936
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 17224 20859 17276 20868
rect 17224 20825 17233 20859
rect 17233 20825 17267 20859
rect 17267 20825 17276 20859
rect 17224 20816 17276 20825
rect 22100 20884 22152 20936
rect 23940 20884 23992 20936
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 24860 21020 24912 21072
rect 22192 20816 22244 20868
rect 22836 20859 22888 20868
rect 22836 20825 22845 20859
rect 22845 20825 22879 20859
rect 22879 20825 22888 20859
rect 22836 20816 22888 20825
rect 22928 20816 22980 20868
rect 23112 20816 23164 20868
rect 24584 20859 24636 20868
rect 24584 20825 24593 20859
rect 24593 20825 24627 20859
rect 24627 20825 24636 20859
rect 24584 20816 24636 20825
rect 24676 20859 24728 20868
rect 24676 20825 24685 20859
rect 24685 20825 24719 20859
rect 24719 20825 24728 20859
rect 24676 20816 24728 20825
rect 24860 20816 24912 20868
rect 8484 20748 8536 20800
rect 8760 20748 8812 20800
rect 9680 20748 9732 20800
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 15476 20748 15528 20800
rect 17040 20748 17092 20800
rect 19248 20791 19300 20800
rect 19248 20757 19257 20791
rect 19257 20757 19291 20791
rect 19291 20757 19300 20791
rect 19248 20748 19300 20757
rect 26056 20952 26108 21004
rect 26332 20816 26384 20868
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 26148 20748 26200 20800
rect 30288 20748 30340 20800
rect 5324 20646 5376 20698
rect 5388 20646 5440 20698
rect 5452 20646 5504 20698
rect 5516 20646 5568 20698
rect 5580 20646 5632 20698
rect 12752 20646 12804 20698
rect 12816 20646 12868 20698
rect 12880 20646 12932 20698
rect 12944 20646 12996 20698
rect 13008 20646 13060 20698
rect 20180 20646 20232 20698
rect 20244 20646 20296 20698
rect 20308 20646 20360 20698
rect 20372 20646 20424 20698
rect 20436 20646 20488 20698
rect 27608 20646 27660 20698
rect 27672 20646 27724 20698
rect 27736 20646 27788 20698
rect 27800 20646 27852 20698
rect 27864 20646 27916 20698
rect 6920 20544 6972 20596
rect 7656 20544 7708 20596
rect 8484 20544 8536 20596
rect 9312 20544 9364 20596
rect 10324 20544 10376 20596
rect 17224 20544 17276 20596
rect 19248 20544 19300 20596
rect 19524 20544 19576 20596
rect 19984 20544 20036 20596
rect 20076 20544 20128 20596
rect 7104 20476 7156 20528
rect 14740 20519 14792 20528
rect 14740 20485 14749 20519
rect 14749 20485 14783 20519
rect 14783 20485 14792 20519
rect 14740 20476 14792 20485
rect 16488 20519 16540 20528
rect 16488 20485 16497 20519
rect 16497 20485 16531 20519
rect 16531 20485 16540 20519
rect 16488 20476 16540 20485
rect 18972 20476 19024 20528
rect 20812 20544 20864 20596
rect 23112 20544 23164 20596
rect 25688 20544 25740 20596
rect 26148 20544 26200 20596
rect 26332 20587 26384 20596
rect 26332 20553 26341 20587
rect 26341 20553 26375 20587
rect 26375 20553 26384 20587
rect 26332 20544 26384 20553
rect 22928 20476 22980 20528
rect 24032 20476 24084 20528
rect 24676 20476 24728 20528
rect 25320 20519 25372 20528
rect 25320 20485 25329 20519
rect 25329 20485 25363 20519
rect 25363 20485 25372 20519
rect 25320 20476 25372 20485
rect 25596 20476 25648 20528
rect 5816 20408 5868 20460
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 9680 20408 9732 20460
rect 11336 20451 11388 20460
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 11336 20417 11345 20451
rect 11345 20417 11379 20451
rect 11379 20417 11388 20451
rect 11336 20408 11388 20417
rect 12624 20408 12676 20460
rect 13544 20408 13596 20460
rect 15844 20408 15896 20460
rect 19432 20451 19484 20460
rect 10048 20340 10100 20392
rect 12532 20340 12584 20392
rect 14280 20340 14332 20392
rect 10324 20315 10376 20324
rect 10324 20281 10333 20315
rect 10333 20281 10367 20315
rect 10367 20281 10376 20315
rect 10324 20272 10376 20281
rect 19432 20417 19433 20451
rect 19433 20417 19467 20451
rect 19467 20417 19484 20451
rect 19432 20408 19484 20417
rect 19984 20451 20036 20460
rect 19984 20417 19993 20451
rect 19993 20417 20027 20451
rect 20027 20417 20036 20451
rect 19984 20408 20036 20417
rect 20076 20408 20128 20460
rect 17960 20340 18012 20392
rect 22376 20451 22428 20460
rect 22376 20417 22385 20451
rect 22385 20417 22419 20451
rect 22419 20417 22428 20451
rect 22376 20408 22428 20417
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 26608 20476 26660 20528
rect 19156 20272 19208 20324
rect 23020 20383 23072 20392
rect 23020 20349 23029 20383
rect 23029 20349 23063 20383
rect 23063 20349 23072 20383
rect 23020 20340 23072 20349
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23296 20340 23348 20349
rect 24492 20340 24544 20392
rect 24860 20340 24912 20392
rect 24952 20272 25004 20324
rect 7380 20204 7432 20256
rect 9772 20204 9824 20256
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 13268 20204 13320 20256
rect 19984 20204 20036 20256
rect 20076 20204 20128 20256
rect 20996 20204 21048 20256
rect 24676 20204 24728 20256
rect 24860 20247 24912 20256
rect 24860 20213 24869 20247
rect 24869 20213 24903 20247
rect 24903 20213 24912 20247
rect 24860 20204 24912 20213
rect 4664 20102 4716 20154
rect 4728 20102 4780 20154
rect 4792 20102 4844 20154
rect 4856 20102 4908 20154
rect 4920 20102 4972 20154
rect 12092 20102 12144 20154
rect 12156 20102 12208 20154
rect 12220 20102 12272 20154
rect 12284 20102 12336 20154
rect 12348 20102 12400 20154
rect 19520 20102 19572 20154
rect 19584 20102 19636 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 26948 20102 27000 20154
rect 27012 20102 27064 20154
rect 27076 20102 27128 20154
rect 27140 20102 27192 20154
rect 27204 20102 27256 20154
rect 7104 20000 7156 20052
rect 8576 20043 8628 20052
rect 8576 20009 8585 20043
rect 8585 20009 8619 20043
rect 8619 20009 8628 20043
rect 8576 20000 8628 20009
rect 10048 20000 10100 20052
rect 10232 20043 10284 20052
rect 10232 20009 10241 20043
rect 10241 20009 10275 20043
rect 10275 20009 10284 20043
rect 10232 20000 10284 20009
rect 10968 20000 11020 20052
rect 11520 20000 11572 20052
rect 940 19728 992 19780
rect 7656 19864 7708 19916
rect 7380 19796 7432 19848
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 8116 19839 8168 19848
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15844 20043 15896 20052
rect 15844 20009 15853 20043
rect 15853 20009 15887 20043
rect 15887 20009 15896 20043
rect 15844 20000 15896 20009
rect 12072 19975 12124 19984
rect 12072 19941 12081 19975
rect 12081 19941 12115 19975
rect 12115 19941 12124 19975
rect 12072 19932 12124 19941
rect 9496 19864 9548 19873
rect 7840 19728 7892 19780
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 9864 19796 9916 19848
rect 5172 19660 5224 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8760 19660 8812 19712
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 14464 19864 14516 19916
rect 15476 19932 15528 19984
rect 17960 19932 18012 19984
rect 15108 19864 15160 19916
rect 17500 19907 17552 19916
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 11244 19728 11296 19780
rect 11704 19771 11756 19780
rect 11704 19737 11713 19771
rect 11713 19737 11747 19771
rect 11747 19737 11756 19771
rect 11704 19728 11756 19737
rect 12072 19771 12124 19780
rect 12072 19737 12081 19771
rect 12081 19737 12115 19771
rect 12115 19737 12124 19771
rect 12072 19728 12124 19737
rect 12440 19796 12492 19848
rect 12532 19796 12584 19848
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 15568 19796 15620 19848
rect 15752 19796 15804 19848
rect 20812 20000 20864 20052
rect 20996 20043 21048 20052
rect 20996 20009 21005 20043
rect 21005 20009 21039 20043
rect 21039 20009 21048 20043
rect 20996 20000 21048 20009
rect 22376 20000 22428 20052
rect 23296 20000 23348 20052
rect 24032 20000 24084 20052
rect 24768 20000 24820 20052
rect 24860 20000 24912 20052
rect 11980 19660 12032 19712
rect 12348 19660 12400 19712
rect 16028 19728 16080 19780
rect 17040 19728 17092 19780
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 20904 19796 20956 19848
rect 22100 19864 22152 19916
rect 23020 19796 23072 19848
rect 30380 19975 30432 19984
rect 30380 19941 30389 19975
rect 30389 19941 30423 19975
rect 30423 19941 30432 19975
rect 30380 19932 30432 19941
rect 13728 19703 13780 19712
rect 13728 19669 13737 19703
rect 13737 19669 13771 19703
rect 13771 19669 13780 19703
rect 13728 19660 13780 19669
rect 19984 19728 20036 19780
rect 20812 19728 20864 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 21824 19728 21876 19780
rect 24676 19796 24728 19848
rect 25044 19728 25096 19780
rect 22928 19703 22980 19712
rect 22928 19669 22937 19703
rect 22937 19669 22971 19703
rect 22971 19669 22980 19703
rect 22928 19660 22980 19669
rect 5324 19558 5376 19610
rect 5388 19558 5440 19610
rect 5452 19558 5504 19610
rect 5516 19558 5568 19610
rect 5580 19558 5632 19610
rect 12752 19558 12804 19610
rect 12816 19558 12868 19610
rect 12880 19558 12932 19610
rect 12944 19558 12996 19610
rect 13008 19558 13060 19610
rect 20180 19558 20232 19610
rect 20244 19558 20296 19610
rect 20308 19558 20360 19610
rect 20372 19558 20424 19610
rect 20436 19558 20488 19610
rect 27608 19558 27660 19610
rect 27672 19558 27724 19610
rect 27736 19558 27788 19610
rect 27800 19558 27852 19610
rect 27864 19558 27916 19610
rect 4344 19456 4396 19508
rect 4436 19456 4488 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 4620 19320 4672 19372
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 5172 19320 5224 19372
rect 6368 19252 6420 19304
rect 7012 19456 7064 19508
rect 7380 19499 7432 19508
rect 7380 19465 7389 19499
rect 7389 19465 7423 19499
rect 7423 19465 7432 19499
rect 7380 19456 7432 19465
rect 7932 19456 7984 19508
rect 8116 19499 8168 19508
rect 8116 19465 8125 19499
rect 8125 19465 8159 19499
rect 8159 19465 8168 19499
rect 8116 19456 8168 19465
rect 8300 19456 8352 19508
rect 12072 19456 12124 19508
rect 7840 19431 7892 19440
rect 7840 19397 7849 19431
rect 7849 19397 7883 19431
rect 7883 19397 7892 19431
rect 7840 19388 7892 19397
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 15568 19456 15620 19508
rect 10600 19320 10652 19372
rect 10968 19320 11020 19372
rect 11612 19320 11664 19372
rect 12348 19363 12400 19372
rect 12348 19329 12357 19363
rect 12357 19329 12391 19363
rect 12391 19329 12400 19363
rect 12348 19320 12400 19329
rect 12440 19320 12492 19372
rect 12624 19320 12676 19372
rect 13176 19320 13228 19372
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 13728 19252 13780 19304
rect 6552 19184 6604 19236
rect 12440 19184 12492 19236
rect 14004 19320 14056 19372
rect 14280 19320 14332 19372
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 14832 19320 14884 19372
rect 15292 19320 15344 19372
rect 5448 19116 5500 19168
rect 9496 19116 9548 19168
rect 9680 19116 9732 19168
rect 10784 19116 10836 19168
rect 11888 19116 11940 19168
rect 14188 19116 14240 19168
rect 14648 19184 14700 19236
rect 14924 19184 14976 19236
rect 15200 19116 15252 19168
rect 15384 19252 15436 19304
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 16488 19388 16540 19440
rect 17040 19388 17092 19440
rect 17500 19388 17552 19440
rect 18880 19388 18932 19440
rect 19432 19388 19484 19440
rect 19524 19388 19576 19440
rect 20904 19499 20956 19508
rect 20904 19465 20913 19499
rect 20913 19465 20947 19499
rect 20947 19465 20956 19499
rect 20904 19456 20956 19465
rect 21824 19456 21876 19508
rect 22928 19456 22980 19508
rect 23388 19456 23440 19508
rect 22192 19388 22244 19440
rect 24768 19388 24820 19440
rect 25872 19388 25924 19440
rect 26240 19456 26292 19508
rect 30288 19320 30340 19372
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 20904 19252 20956 19304
rect 15844 19227 15896 19236
rect 15844 19193 15853 19227
rect 15853 19193 15887 19227
rect 15887 19193 15896 19227
rect 15844 19184 15896 19193
rect 16396 19159 16448 19168
rect 16396 19125 16405 19159
rect 16405 19125 16439 19159
rect 16439 19125 16448 19159
rect 16396 19116 16448 19125
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 21916 19116 21968 19125
rect 24860 19295 24912 19304
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 24952 19116 25004 19168
rect 4664 19014 4716 19066
rect 4728 19014 4780 19066
rect 4792 19014 4844 19066
rect 4856 19014 4908 19066
rect 4920 19014 4972 19066
rect 12092 19014 12144 19066
rect 12156 19014 12208 19066
rect 12220 19014 12272 19066
rect 12284 19014 12336 19066
rect 12348 19014 12400 19066
rect 19520 19014 19572 19066
rect 19584 19014 19636 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 26948 19014 27000 19066
rect 27012 19014 27064 19066
rect 27076 19014 27128 19066
rect 27140 19014 27192 19066
rect 27204 19014 27256 19066
rect 3608 18912 3660 18964
rect 6552 18912 6604 18964
rect 6644 18912 6696 18964
rect 940 18708 992 18760
rect 4344 18844 4396 18896
rect 5080 18844 5132 18896
rect 5448 18776 5500 18828
rect 4436 18708 4488 18760
rect 5172 18708 5224 18760
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 9956 18844 10008 18896
rect 10048 18844 10100 18896
rect 11152 18912 11204 18964
rect 11704 18912 11756 18964
rect 11796 18912 11848 18964
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 13360 18912 13412 18964
rect 14556 18912 14608 18964
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 21364 18912 21416 18964
rect 24860 18912 24912 18964
rect 6736 18776 6788 18828
rect 6920 18751 6972 18760
rect 6920 18717 6929 18751
rect 6929 18717 6963 18751
rect 6963 18717 6972 18751
rect 6920 18708 6972 18717
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 7196 18708 7248 18760
rect 10140 18708 10192 18760
rect 10784 18776 10836 18828
rect 10968 18708 11020 18760
rect 9680 18640 9732 18692
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 10508 18640 10560 18692
rect 10876 18683 10928 18692
rect 10876 18649 10885 18683
rect 10885 18649 10919 18683
rect 10919 18649 10928 18683
rect 10876 18640 10928 18649
rect 4344 18572 4396 18624
rect 4988 18572 5040 18624
rect 6092 18572 6144 18624
rect 10416 18572 10468 18624
rect 11336 18572 11388 18624
rect 14372 18844 14424 18896
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 14188 18776 14240 18828
rect 15660 18776 15712 18828
rect 13268 18708 13320 18760
rect 12532 18640 12584 18692
rect 12624 18640 12676 18692
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 14832 18708 14884 18760
rect 16396 18708 16448 18760
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 20076 18844 20128 18896
rect 20904 18776 20956 18828
rect 20996 18819 21048 18828
rect 20996 18785 21005 18819
rect 21005 18785 21039 18819
rect 21039 18785 21048 18819
rect 20996 18776 21048 18785
rect 21456 18887 21508 18896
rect 21456 18853 21465 18887
rect 21465 18853 21499 18887
rect 21499 18853 21508 18887
rect 21456 18844 21508 18853
rect 25228 18887 25280 18896
rect 25228 18853 25237 18887
rect 25237 18853 25271 18887
rect 25271 18853 25280 18887
rect 25228 18844 25280 18853
rect 19248 18708 19300 18760
rect 18420 18640 18472 18692
rect 21088 18708 21140 18760
rect 22100 18819 22152 18828
rect 22100 18785 22109 18819
rect 22109 18785 22143 18819
rect 22143 18785 22152 18819
rect 22100 18776 22152 18785
rect 21916 18708 21968 18760
rect 24400 18776 24452 18828
rect 15476 18572 15528 18624
rect 16488 18572 16540 18624
rect 18328 18572 18380 18624
rect 19892 18615 19944 18624
rect 19892 18581 19901 18615
rect 19901 18581 19935 18615
rect 19935 18581 19944 18615
rect 19892 18572 19944 18581
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 22376 18683 22428 18692
rect 22376 18649 22385 18683
rect 22385 18649 22419 18683
rect 22419 18649 22428 18683
rect 22376 18640 22428 18649
rect 24952 18776 25004 18828
rect 25228 18708 25280 18760
rect 26240 18819 26292 18828
rect 26240 18785 26249 18819
rect 26249 18785 26283 18819
rect 26283 18785 26292 18819
rect 26240 18776 26292 18785
rect 26608 18708 26660 18760
rect 24492 18640 24544 18692
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 26424 18615 26476 18624
rect 26424 18581 26433 18615
rect 26433 18581 26467 18615
rect 26467 18581 26476 18615
rect 26424 18572 26476 18581
rect 30380 18615 30432 18624
rect 30380 18581 30389 18615
rect 30389 18581 30423 18615
rect 30423 18581 30432 18615
rect 30380 18572 30432 18581
rect 5324 18470 5376 18522
rect 5388 18470 5440 18522
rect 5452 18470 5504 18522
rect 5516 18470 5568 18522
rect 5580 18470 5632 18522
rect 12752 18470 12804 18522
rect 12816 18470 12868 18522
rect 12880 18470 12932 18522
rect 12944 18470 12996 18522
rect 13008 18470 13060 18522
rect 20180 18470 20232 18522
rect 20244 18470 20296 18522
rect 20308 18470 20360 18522
rect 20372 18470 20424 18522
rect 20436 18470 20488 18522
rect 27608 18470 27660 18522
rect 27672 18470 27724 18522
rect 27736 18470 27788 18522
rect 27800 18470 27852 18522
rect 27864 18470 27916 18522
rect 5080 18300 5132 18352
rect 5908 18300 5960 18352
rect 6552 18368 6604 18420
rect 9404 18368 9456 18420
rect 11612 18368 11664 18420
rect 11704 18368 11756 18420
rect 12256 18368 12308 18420
rect 12624 18411 12676 18420
rect 6736 18300 6788 18352
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 7656 18300 7708 18352
rect 8024 18300 8076 18352
rect 8668 18300 8720 18352
rect 11888 18300 11940 18352
rect 7472 18232 7524 18284
rect 8484 18232 8536 18284
rect 7012 18164 7064 18216
rect 7748 18164 7800 18216
rect 9496 18207 9548 18216
rect 9496 18173 9505 18207
rect 9505 18173 9539 18207
rect 9539 18173 9548 18207
rect 9496 18164 9548 18173
rect 5172 18096 5224 18148
rect 7380 18096 7432 18148
rect 9864 18164 9916 18216
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 10968 18232 11020 18284
rect 10508 18164 10560 18216
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 11612 18232 11664 18284
rect 12624 18377 12633 18411
rect 12633 18377 12667 18411
rect 12667 18377 12676 18411
rect 12624 18368 12676 18377
rect 14372 18368 14424 18420
rect 7288 18028 7340 18080
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 8024 18028 8076 18080
rect 10140 18096 10192 18148
rect 10232 18096 10284 18148
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 11888 18207 11940 18216
rect 11888 18173 11897 18207
rect 11897 18173 11931 18207
rect 11931 18173 11940 18207
rect 11888 18164 11940 18173
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 11612 18028 11664 18080
rect 12256 18096 12308 18148
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 16948 18275 17000 18284
rect 16948 18241 16957 18275
rect 16957 18241 16991 18275
rect 16991 18241 17000 18275
rect 16948 18232 17000 18241
rect 17408 18232 17460 18284
rect 20076 18368 20128 18420
rect 20352 18368 20404 18420
rect 21272 18368 21324 18420
rect 22376 18411 22428 18420
rect 22376 18377 22385 18411
rect 22385 18377 22419 18411
rect 22419 18377 22428 18411
rect 22376 18368 22428 18377
rect 22836 18411 22888 18420
rect 22836 18377 22845 18411
rect 22845 18377 22879 18411
rect 22879 18377 22888 18411
rect 22836 18368 22888 18377
rect 25872 18368 25924 18420
rect 19064 18300 19116 18352
rect 19248 18300 19300 18352
rect 21088 18300 21140 18352
rect 15200 18164 15252 18216
rect 12440 18028 12492 18080
rect 13176 18028 13228 18080
rect 14188 18028 14240 18080
rect 16304 18096 16356 18148
rect 19892 18275 19944 18284
rect 19892 18241 19901 18275
rect 19901 18241 19935 18275
rect 19935 18241 19944 18275
rect 19892 18232 19944 18241
rect 20720 18232 20772 18284
rect 21272 18232 21324 18284
rect 22560 18275 22612 18284
rect 22560 18241 22569 18275
rect 22569 18241 22603 18275
rect 22603 18241 22612 18275
rect 22560 18232 22612 18241
rect 24492 18300 24544 18352
rect 25964 18300 26016 18352
rect 27436 18300 27488 18352
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 25044 18232 25096 18284
rect 20076 18096 20128 18148
rect 23572 18164 23624 18216
rect 23848 18164 23900 18216
rect 16764 18071 16816 18080
rect 16764 18037 16773 18071
rect 16773 18037 16807 18071
rect 16807 18037 16816 18071
rect 16764 18028 16816 18037
rect 17500 18071 17552 18080
rect 17500 18037 17509 18071
rect 17509 18037 17543 18071
rect 17543 18037 17552 18071
rect 17500 18028 17552 18037
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 22652 18028 22704 18080
rect 30288 18028 30340 18080
rect 4664 17926 4716 17978
rect 4728 17926 4780 17978
rect 4792 17926 4844 17978
rect 4856 17926 4908 17978
rect 4920 17926 4972 17978
rect 12092 17926 12144 17978
rect 12156 17926 12208 17978
rect 12220 17926 12272 17978
rect 12284 17926 12336 17978
rect 12348 17926 12400 17978
rect 19520 17926 19572 17978
rect 19584 17926 19636 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 26948 17926 27000 17978
rect 27012 17926 27064 17978
rect 27076 17926 27128 17978
rect 27140 17926 27192 17978
rect 27204 17926 27256 17978
rect 4988 17867 5040 17876
rect 4988 17833 4997 17867
rect 4997 17833 5031 17867
rect 5031 17833 5040 17867
rect 4988 17824 5040 17833
rect 5356 17824 5408 17876
rect 6184 17824 6236 17876
rect 6460 17824 6512 17876
rect 9496 17824 9548 17876
rect 9772 17824 9824 17876
rect 10692 17824 10744 17876
rect 10876 17824 10928 17876
rect 16948 17824 17000 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 21088 17824 21140 17876
rect 21456 17824 21508 17876
rect 5724 17731 5776 17740
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 6644 17756 6696 17808
rect 6736 17756 6788 17808
rect 11244 17756 11296 17808
rect 14188 17756 14240 17808
rect 16672 17756 16724 17808
rect 6000 17688 6052 17740
rect 5908 17663 5960 17672
rect 5908 17629 5917 17663
rect 5917 17629 5951 17663
rect 5951 17629 5960 17663
rect 5908 17620 5960 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 9128 17688 9180 17740
rect 6736 17663 6788 17672
rect 6736 17629 6745 17663
rect 6745 17629 6779 17663
rect 6779 17629 6788 17663
rect 6736 17620 6788 17629
rect 6920 17620 6972 17672
rect 7748 17620 7800 17672
rect 8668 17620 8720 17672
rect 10508 17688 10560 17740
rect 10876 17688 10928 17740
rect 11980 17688 12032 17740
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 17040 17688 17092 17740
rect 18972 17756 19024 17808
rect 17408 17688 17460 17740
rect 9772 17620 9824 17672
rect 4988 17484 5040 17536
rect 6276 17552 6328 17604
rect 9496 17552 9548 17604
rect 10416 17620 10468 17672
rect 13728 17663 13780 17672
rect 13728 17629 13737 17663
rect 13737 17629 13771 17663
rect 13771 17629 13780 17663
rect 13728 17620 13780 17629
rect 16212 17620 16264 17672
rect 10232 17552 10284 17604
rect 6828 17484 6880 17536
rect 7012 17527 7064 17536
rect 7012 17493 7021 17527
rect 7021 17493 7055 17527
rect 7055 17493 7064 17527
rect 7012 17484 7064 17493
rect 8300 17484 8352 17536
rect 9036 17484 9088 17536
rect 13636 17484 13688 17536
rect 15292 17552 15344 17604
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 16672 17663 16724 17672
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 18696 17620 18748 17672
rect 20352 17731 20404 17740
rect 20352 17697 20361 17731
rect 20361 17697 20395 17731
rect 20395 17697 20404 17731
rect 20352 17688 20404 17697
rect 24768 17688 24820 17740
rect 14740 17484 14792 17536
rect 15844 17484 15896 17536
rect 27344 17663 27396 17672
rect 27344 17629 27353 17663
rect 27353 17629 27387 17663
rect 27387 17629 27396 17663
rect 27344 17620 27396 17629
rect 27436 17663 27488 17672
rect 27436 17629 27445 17663
rect 27445 17629 27479 17663
rect 27479 17629 27488 17663
rect 27436 17620 27488 17629
rect 20996 17552 21048 17604
rect 25136 17595 25188 17604
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 17592 17484 17644 17536
rect 19800 17484 19852 17536
rect 19892 17527 19944 17536
rect 19892 17493 19901 17527
rect 19901 17493 19935 17527
rect 19935 17493 19944 17527
rect 19892 17484 19944 17493
rect 26700 17527 26752 17536
rect 26700 17493 26709 17527
rect 26709 17493 26743 17527
rect 26743 17493 26752 17527
rect 26700 17484 26752 17493
rect 5324 17382 5376 17434
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 12752 17382 12804 17434
rect 12816 17382 12868 17434
rect 12880 17382 12932 17434
rect 12944 17382 12996 17434
rect 13008 17382 13060 17434
rect 20180 17382 20232 17434
rect 20244 17382 20296 17434
rect 20308 17382 20360 17434
rect 20372 17382 20424 17434
rect 20436 17382 20488 17434
rect 27608 17382 27660 17434
rect 27672 17382 27724 17434
rect 27736 17382 27788 17434
rect 27800 17382 27852 17434
rect 27864 17382 27916 17434
rect 4988 17323 5040 17332
rect 4988 17289 4997 17323
rect 4997 17289 5031 17323
rect 5031 17289 5040 17323
rect 4988 17280 5040 17289
rect 5172 17280 5224 17332
rect 6460 17280 6512 17332
rect 6552 17280 6604 17332
rect 7196 17280 7248 17332
rect 7012 17212 7064 17264
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 5080 17144 5132 17196
rect 5724 17144 5776 17196
rect 5908 17144 5960 17196
rect 940 17076 992 17128
rect 1676 17119 1728 17128
rect 1676 17085 1685 17119
rect 1685 17085 1719 17119
rect 1719 17085 1728 17119
rect 1676 17076 1728 17085
rect 6276 17144 6328 17196
rect 6460 17119 6512 17128
rect 6460 17085 6469 17119
rect 6469 17085 6503 17119
rect 6503 17085 6512 17119
rect 6460 17076 6512 17085
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 8116 17144 8168 17196
rect 6828 17076 6880 17128
rect 7196 17076 7248 17128
rect 8760 17144 8812 17196
rect 9220 17212 9272 17264
rect 9496 17212 9548 17264
rect 9680 17212 9732 17264
rect 9956 17212 10008 17264
rect 11152 17280 11204 17332
rect 11612 17323 11664 17332
rect 11612 17289 11621 17323
rect 11621 17289 11655 17323
rect 11655 17289 11664 17323
rect 11612 17280 11664 17289
rect 13084 17280 13136 17332
rect 13728 17280 13780 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 15292 17280 15344 17332
rect 15476 17280 15528 17332
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 16580 17280 16632 17332
rect 18972 17280 19024 17332
rect 20076 17323 20128 17332
rect 20076 17289 20085 17323
rect 20085 17289 20119 17323
rect 20119 17289 20128 17323
rect 20076 17280 20128 17289
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 25136 17280 25188 17332
rect 26700 17280 26752 17332
rect 11336 17212 11388 17264
rect 12532 17212 12584 17264
rect 10968 17144 11020 17196
rect 8668 17076 8720 17128
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 9312 17076 9364 17128
rect 6276 17008 6328 17060
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 8760 16940 8812 16992
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 10140 17076 10192 17128
rect 10784 17076 10836 17128
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 12440 17187 12492 17196
rect 12440 17153 12446 17187
rect 12446 17153 12492 17187
rect 12440 17144 12492 17153
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 11980 17076 12032 17128
rect 13636 17144 13688 17196
rect 14464 17144 14516 17196
rect 15752 17212 15804 17264
rect 15844 17212 15896 17264
rect 16488 17212 16540 17264
rect 19340 17212 19392 17264
rect 14556 17076 14608 17128
rect 16028 17144 16080 17196
rect 16396 17144 16448 17196
rect 16948 17144 17000 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 24124 17212 24176 17264
rect 12072 17008 12124 17060
rect 18236 17008 18288 17060
rect 11612 16940 11664 16992
rect 12440 16940 12492 16992
rect 17960 16940 18012 16992
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 18972 17076 19024 17128
rect 21272 17076 21324 17128
rect 22008 17119 22060 17128
rect 22008 17085 22017 17119
rect 22017 17085 22051 17119
rect 22051 17085 22060 17119
rect 22008 17076 22060 17085
rect 22284 17144 22336 17196
rect 22744 17144 22796 17196
rect 23388 17144 23440 17196
rect 23572 17187 23624 17196
rect 23572 17153 23581 17187
rect 23581 17153 23615 17187
rect 23615 17153 23624 17187
rect 23572 17144 23624 17153
rect 24952 17187 25004 17196
rect 24952 17153 24961 17187
rect 24961 17153 24995 17187
rect 24995 17153 25004 17187
rect 24952 17144 25004 17153
rect 27344 17144 27396 17196
rect 22192 17008 22244 17060
rect 19156 16940 19208 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20904 16940 20956 16992
rect 21548 16940 21600 16992
rect 26148 17008 26200 17060
rect 30380 17051 30432 17060
rect 30380 17017 30389 17051
rect 30389 17017 30423 17051
rect 30423 17017 30432 17051
rect 30380 17008 30432 17017
rect 22376 16940 22428 16992
rect 23388 16940 23440 16992
rect 25044 16940 25096 16992
rect 25504 16940 25556 16992
rect 25964 16940 26016 16992
rect 4664 16838 4716 16890
rect 4728 16838 4780 16890
rect 4792 16838 4844 16890
rect 4856 16838 4908 16890
rect 4920 16838 4972 16890
rect 12092 16838 12144 16890
rect 12156 16838 12208 16890
rect 12220 16838 12272 16890
rect 12284 16838 12336 16890
rect 12348 16838 12400 16890
rect 19520 16838 19572 16890
rect 19584 16838 19636 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 26948 16838 27000 16890
rect 27012 16838 27064 16890
rect 27076 16838 27128 16890
rect 27140 16838 27192 16890
rect 27204 16838 27256 16890
rect 1676 16736 1728 16788
rect 6460 16736 6512 16788
rect 6736 16736 6788 16788
rect 7196 16736 7248 16788
rect 8944 16736 8996 16788
rect 9036 16736 9088 16788
rect 9128 16736 9180 16788
rect 9496 16736 9548 16788
rect 11796 16736 11848 16788
rect 4528 16600 4580 16652
rect 5172 16532 5224 16584
rect 8300 16600 8352 16652
rect 9128 16600 9180 16652
rect 7472 16532 7524 16584
rect 9772 16600 9824 16652
rect 10324 16600 10376 16652
rect 11152 16668 11204 16720
rect 12624 16736 12676 16788
rect 13084 16779 13136 16788
rect 13084 16745 13093 16779
rect 13093 16745 13127 16779
rect 13127 16745 13136 16779
rect 13084 16736 13136 16745
rect 15568 16779 15620 16788
rect 15568 16745 15577 16779
rect 15577 16745 15611 16779
rect 15611 16745 15620 16779
rect 15568 16736 15620 16745
rect 19248 16736 19300 16788
rect 19340 16779 19392 16788
rect 19340 16745 19349 16779
rect 19349 16745 19383 16779
rect 19383 16745 19392 16779
rect 19340 16736 19392 16745
rect 18604 16668 18656 16720
rect 10416 16532 10468 16584
rect 10508 16532 10560 16584
rect 3424 16464 3476 16516
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11060 16600 11112 16652
rect 10784 16575 10836 16584
rect 10784 16541 10816 16575
rect 10816 16541 10836 16575
rect 10784 16532 10836 16541
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 12440 16532 12492 16584
rect 12532 16575 12584 16584
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 12532 16532 12584 16541
rect 15292 16532 15344 16584
rect 940 16396 992 16448
rect 4436 16396 4488 16448
rect 10508 16439 10560 16448
rect 10508 16405 10517 16439
rect 10517 16405 10551 16439
rect 10551 16405 10560 16439
rect 10508 16396 10560 16405
rect 11336 16396 11388 16448
rect 13176 16464 13228 16516
rect 13728 16464 13780 16516
rect 13820 16507 13872 16516
rect 13820 16473 13829 16507
rect 13829 16473 13863 16507
rect 13863 16473 13872 16507
rect 13820 16464 13872 16473
rect 14280 16507 14332 16516
rect 14280 16473 14289 16507
rect 14289 16473 14323 16507
rect 14323 16473 14332 16507
rect 14280 16464 14332 16473
rect 14832 16464 14884 16516
rect 15016 16464 15068 16516
rect 18696 16600 18748 16652
rect 18972 16600 19024 16652
rect 19064 16600 19116 16652
rect 19892 16736 19944 16788
rect 20720 16736 20772 16788
rect 22744 16736 22796 16788
rect 22836 16736 22888 16788
rect 19984 16643 20036 16652
rect 19984 16609 19993 16643
rect 19993 16609 20027 16643
rect 20027 16609 20036 16643
rect 20904 16668 20956 16720
rect 20996 16711 21048 16720
rect 20996 16677 21005 16711
rect 21005 16677 21039 16711
rect 21039 16677 21048 16711
rect 20996 16668 21048 16677
rect 19984 16600 20036 16609
rect 20628 16643 20680 16652
rect 20628 16609 20637 16643
rect 20637 16609 20671 16643
rect 20671 16609 20680 16643
rect 20628 16600 20680 16609
rect 21732 16643 21784 16652
rect 21732 16609 21741 16643
rect 21741 16609 21775 16643
rect 21775 16609 21784 16643
rect 21732 16600 21784 16609
rect 22928 16643 22980 16652
rect 22928 16609 22937 16643
rect 22937 16609 22971 16643
rect 22971 16609 22980 16643
rect 22928 16600 22980 16609
rect 24124 16711 24176 16720
rect 24124 16677 24133 16711
rect 24133 16677 24167 16711
rect 24167 16677 24176 16711
rect 24124 16668 24176 16677
rect 25596 16779 25648 16788
rect 25596 16745 25605 16779
rect 25605 16745 25639 16779
rect 25639 16745 25648 16779
rect 25596 16736 25648 16745
rect 20168 16532 20220 16584
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 20812 16575 20864 16584
rect 20812 16541 20821 16575
rect 20821 16541 20855 16575
rect 20855 16541 20864 16575
rect 20812 16532 20864 16541
rect 20904 16532 20956 16584
rect 22192 16575 22244 16584
rect 22192 16541 22201 16575
rect 22201 16541 22235 16575
rect 22235 16541 22244 16575
rect 22192 16532 22244 16541
rect 22376 16575 22428 16584
rect 22376 16541 22385 16575
rect 22385 16541 22419 16575
rect 22419 16541 22428 16575
rect 22376 16532 22428 16541
rect 22652 16575 22704 16584
rect 22652 16541 22687 16575
rect 22687 16541 22704 16575
rect 22652 16532 22704 16541
rect 22836 16575 22888 16584
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 23940 16575 23992 16584
rect 23940 16541 23949 16575
rect 23949 16541 23983 16575
rect 23983 16541 23992 16575
rect 23940 16532 23992 16541
rect 19064 16464 19116 16516
rect 13360 16396 13412 16448
rect 17040 16439 17092 16448
rect 17040 16405 17049 16439
rect 17049 16405 17083 16439
rect 17083 16405 17092 16439
rect 17040 16396 17092 16405
rect 22468 16507 22520 16516
rect 22468 16473 22477 16507
rect 22477 16473 22511 16507
rect 22511 16473 22520 16507
rect 22468 16464 22520 16473
rect 22560 16507 22612 16516
rect 22560 16473 22569 16507
rect 22569 16473 22603 16507
rect 22603 16473 22612 16507
rect 22560 16464 22612 16473
rect 24676 16532 24728 16584
rect 24860 16575 24912 16584
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 25044 16600 25096 16652
rect 25688 16711 25740 16720
rect 25688 16677 25697 16711
rect 25697 16677 25731 16711
rect 25731 16677 25740 16711
rect 26332 16736 26384 16788
rect 25688 16668 25740 16677
rect 25504 16643 25556 16652
rect 25504 16609 25513 16643
rect 25513 16609 25547 16643
rect 25547 16609 25556 16643
rect 25504 16600 25556 16609
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 25780 16575 25832 16584
rect 25780 16541 25789 16575
rect 25789 16541 25823 16575
rect 25823 16541 25832 16575
rect 25780 16532 25832 16541
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 27344 16600 27396 16652
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 24768 16396 24820 16448
rect 30932 16464 30984 16516
rect 5324 16294 5376 16346
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 12752 16294 12804 16346
rect 12816 16294 12868 16346
rect 12880 16294 12932 16346
rect 12944 16294 12996 16346
rect 13008 16294 13060 16346
rect 20180 16294 20232 16346
rect 20244 16294 20296 16346
rect 20308 16294 20360 16346
rect 20372 16294 20424 16346
rect 20436 16294 20488 16346
rect 27608 16294 27660 16346
rect 27672 16294 27724 16346
rect 27736 16294 27788 16346
rect 27800 16294 27852 16346
rect 27864 16294 27916 16346
rect 4436 16192 4488 16244
rect 5172 16192 5224 16244
rect 5448 16192 5500 16244
rect 6092 16192 6144 16244
rect 7472 16235 7524 16244
rect 7472 16201 7481 16235
rect 7481 16201 7515 16235
rect 7515 16201 7524 16235
rect 7472 16192 7524 16201
rect 9220 16192 9272 16244
rect 5908 16099 5960 16108
rect 5908 16065 5917 16099
rect 5917 16065 5951 16099
rect 5951 16065 5960 16099
rect 5908 16056 5960 16065
rect 6092 16099 6144 16108
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 6092 16056 6144 16065
rect 940 15852 992 15904
rect 4436 15988 4488 16040
rect 5080 16031 5132 16040
rect 5080 15997 5089 16031
rect 5089 15997 5123 16031
rect 5123 15997 5132 16031
rect 5080 15988 5132 15997
rect 6276 15988 6328 16040
rect 10508 16192 10560 16244
rect 11980 16192 12032 16244
rect 11428 16124 11480 16176
rect 11612 16124 11664 16176
rect 10416 16056 10468 16108
rect 10784 15988 10836 16040
rect 13636 16056 13688 16108
rect 14832 16056 14884 16108
rect 5908 15920 5960 15972
rect 7012 15920 7064 15972
rect 7472 15920 7524 15972
rect 10692 15920 10744 15972
rect 5356 15852 5408 15904
rect 6000 15895 6052 15904
rect 6000 15861 6009 15895
rect 6009 15861 6043 15895
rect 6043 15861 6052 15895
rect 6000 15852 6052 15861
rect 7196 15852 7248 15904
rect 9312 15895 9364 15904
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 15844 16056 15896 16108
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 16580 16056 16632 16108
rect 17868 16192 17920 16244
rect 18236 16192 18288 16244
rect 20536 16235 20588 16244
rect 20536 16201 20545 16235
rect 20545 16201 20579 16235
rect 20579 16201 20588 16235
rect 20536 16192 20588 16201
rect 20720 16192 20772 16244
rect 21088 16192 21140 16244
rect 17040 16124 17092 16176
rect 22468 16192 22520 16244
rect 19064 16056 19116 16108
rect 20996 16124 21048 16176
rect 21732 16124 21784 16176
rect 22284 16124 22336 16176
rect 22652 16124 22704 16176
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 11428 15920 11480 15972
rect 13820 15920 13872 15972
rect 14924 15920 14976 15972
rect 15384 15920 15436 15972
rect 13636 15852 13688 15904
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 23940 16192 23992 16244
rect 24492 16192 24544 16244
rect 25596 16192 25648 16244
rect 25780 16192 25832 16244
rect 26332 16192 26384 16244
rect 24400 16124 24452 16176
rect 25136 16124 25188 16176
rect 24768 16056 24820 16108
rect 25228 16056 25280 16108
rect 25688 16056 25740 16108
rect 18420 15963 18472 15972
rect 18420 15929 18429 15963
rect 18429 15929 18463 15963
rect 18463 15929 18472 15963
rect 18420 15920 18472 15929
rect 24952 15963 25004 15972
rect 24952 15929 24961 15963
rect 24961 15929 24995 15963
rect 24995 15929 25004 15963
rect 24952 15920 25004 15929
rect 17684 15852 17736 15904
rect 20720 15852 20772 15904
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 24676 15852 24728 15904
rect 25136 15852 25188 15904
rect 25780 15852 25832 15904
rect 25872 15895 25924 15904
rect 25872 15861 25881 15895
rect 25881 15861 25915 15895
rect 25915 15861 25924 15895
rect 25872 15852 25924 15861
rect 26424 15852 26476 15904
rect 30380 15895 30432 15904
rect 30380 15861 30389 15895
rect 30389 15861 30423 15895
rect 30423 15861 30432 15895
rect 30380 15852 30432 15861
rect 4664 15750 4716 15802
rect 4728 15750 4780 15802
rect 4792 15750 4844 15802
rect 4856 15750 4908 15802
rect 4920 15750 4972 15802
rect 12092 15750 12144 15802
rect 12156 15750 12208 15802
rect 12220 15750 12272 15802
rect 12284 15750 12336 15802
rect 12348 15750 12400 15802
rect 19520 15750 19572 15802
rect 19584 15750 19636 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 26948 15750 27000 15802
rect 27012 15750 27064 15802
rect 27076 15750 27128 15802
rect 27140 15750 27192 15802
rect 27204 15750 27256 15802
rect 4436 15648 4488 15700
rect 4896 15648 4948 15700
rect 5448 15648 5500 15700
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 6000 15648 6052 15700
rect 6276 15648 6328 15700
rect 7932 15648 7984 15700
rect 9312 15691 9364 15700
rect 5816 15580 5868 15632
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 6000 15419 6052 15428
rect 6000 15385 6009 15419
rect 6009 15385 6043 15419
rect 6043 15385 6052 15419
rect 6000 15376 6052 15385
rect 6368 15376 6420 15428
rect 7012 15444 7064 15496
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 7472 15444 7524 15496
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 9312 15657 9342 15691
rect 9342 15657 9364 15691
rect 9312 15648 9364 15657
rect 10324 15648 10376 15700
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 15660 15648 15712 15700
rect 18420 15648 18472 15700
rect 24860 15648 24912 15700
rect 25136 15648 25188 15700
rect 25320 15648 25372 15700
rect 25872 15648 25924 15700
rect 10784 15623 10836 15632
rect 10784 15589 10793 15623
rect 10793 15589 10827 15623
rect 10827 15589 10836 15623
rect 10784 15580 10836 15589
rect 9312 15512 9364 15564
rect 12532 15512 12584 15564
rect 13728 15580 13780 15632
rect 8116 15308 8168 15360
rect 11520 15444 11572 15496
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11244 15308 11296 15360
rect 12072 15419 12124 15428
rect 12072 15385 12081 15419
rect 12081 15385 12115 15419
rect 12115 15385 12124 15419
rect 12072 15376 12124 15385
rect 12624 15376 12676 15428
rect 14648 15555 14700 15564
rect 14648 15521 14657 15555
rect 14657 15521 14691 15555
rect 14691 15521 14700 15555
rect 14648 15512 14700 15521
rect 14740 15444 14792 15496
rect 15108 15444 15160 15496
rect 16028 15580 16080 15632
rect 23756 15580 23808 15632
rect 17316 15555 17368 15564
rect 17316 15521 17325 15555
rect 17325 15521 17359 15555
rect 17359 15521 17368 15555
rect 17316 15512 17368 15521
rect 16672 15444 16724 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 21272 15444 21324 15496
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 25044 15444 25096 15496
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 13728 15376 13780 15428
rect 20904 15376 20956 15428
rect 13544 15351 13596 15360
rect 13544 15317 13553 15351
rect 13553 15317 13587 15351
rect 13587 15317 13596 15351
rect 13544 15308 13596 15317
rect 16948 15308 17000 15360
rect 19340 15308 19392 15360
rect 20812 15308 20864 15360
rect 24492 15376 24544 15428
rect 25688 15512 25740 15564
rect 25780 15512 25832 15564
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 24952 15351 25004 15360
rect 24952 15317 24961 15351
rect 24961 15317 24995 15351
rect 24995 15317 25004 15351
rect 24952 15308 25004 15317
rect 25964 15487 26016 15496
rect 25964 15453 25973 15487
rect 25973 15453 26007 15487
rect 26007 15453 26016 15487
rect 25964 15444 26016 15453
rect 30288 15308 30340 15360
rect 5324 15206 5376 15258
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 12752 15206 12804 15258
rect 12816 15206 12868 15258
rect 12880 15206 12932 15258
rect 12944 15206 12996 15258
rect 13008 15206 13060 15258
rect 20180 15206 20232 15258
rect 20244 15206 20296 15258
rect 20308 15206 20360 15258
rect 20372 15206 20424 15258
rect 20436 15206 20488 15258
rect 27608 15206 27660 15258
rect 27672 15206 27724 15258
rect 27736 15206 27788 15258
rect 27800 15206 27852 15258
rect 27864 15206 27916 15258
rect 5724 15104 5776 15156
rect 6184 15104 6236 15156
rect 6368 15036 6420 15088
rect 8024 15036 8076 15088
rect 5080 14968 5132 15020
rect 4896 14832 4948 14884
rect 5264 14968 5316 15020
rect 6000 15011 6052 15020
rect 6000 14977 6009 15011
rect 6009 14977 6043 15011
rect 6043 14977 6052 15011
rect 6000 14968 6052 14977
rect 6276 14968 6328 15020
rect 7472 14968 7524 15020
rect 8300 14968 8352 15020
rect 7104 14900 7156 14952
rect 8116 14900 8168 14952
rect 10600 15079 10652 15088
rect 10600 15045 10609 15079
rect 10609 15045 10643 15079
rect 10643 15045 10652 15079
rect 10600 15036 10652 15045
rect 12072 15104 12124 15156
rect 12624 15104 12676 15156
rect 18880 15104 18932 15156
rect 21548 15104 21600 15156
rect 22008 15104 22060 15156
rect 22100 15104 22152 15156
rect 10324 14968 10376 15020
rect 11428 14968 11480 15020
rect 8576 14900 8628 14952
rect 9220 14900 9272 14952
rect 12532 14900 12584 14952
rect 12624 14900 12676 14952
rect 13268 14968 13320 15020
rect 5632 14832 5684 14884
rect 6092 14832 6144 14884
rect 13544 14968 13596 15020
rect 14648 14968 14700 15020
rect 4528 14764 4580 14816
rect 5172 14764 5224 14816
rect 5908 14764 5960 14816
rect 13544 14832 13596 14884
rect 14556 14832 14608 14884
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 15844 14968 15896 15020
rect 15936 15011 15988 15020
rect 15936 14977 15945 15011
rect 15945 14977 15979 15011
rect 15979 14977 15988 15011
rect 15936 14968 15988 14977
rect 16672 14968 16724 15020
rect 17316 15036 17368 15088
rect 19340 15036 19392 15088
rect 24768 15104 24820 15156
rect 25044 15104 25096 15156
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 8208 14764 8260 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 11152 14764 11204 14816
rect 13636 14764 13688 14816
rect 14280 14807 14332 14816
rect 14280 14773 14289 14807
rect 14289 14773 14323 14807
rect 14323 14773 14332 14807
rect 14280 14764 14332 14773
rect 16304 14943 16356 14952
rect 16304 14909 16313 14943
rect 16313 14909 16347 14943
rect 16347 14909 16356 14943
rect 16304 14900 16356 14909
rect 17684 14900 17736 14952
rect 16028 14764 16080 14816
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 18604 14943 18656 14952
rect 18604 14909 18613 14943
rect 18613 14909 18647 14943
rect 18647 14909 18656 14943
rect 18604 14900 18656 14909
rect 19156 15011 19208 15020
rect 19156 14977 19165 15011
rect 19165 14977 19199 15011
rect 19199 14977 19208 15011
rect 19156 14968 19208 14977
rect 20536 14968 20588 15020
rect 20720 14968 20772 15020
rect 22100 14900 22152 14952
rect 24492 15036 24544 15088
rect 20444 14832 20496 14884
rect 20720 14764 20772 14816
rect 21916 14764 21968 14816
rect 22284 14764 22336 14816
rect 22744 14764 22796 14816
rect 24768 14764 24820 14816
rect 24860 14764 24912 14816
rect 25228 14764 25280 14816
rect 30196 14764 30248 14816
rect 4664 14662 4716 14714
rect 4728 14662 4780 14714
rect 4792 14662 4844 14714
rect 4856 14662 4908 14714
rect 4920 14662 4972 14714
rect 12092 14662 12144 14714
rect 12156 14662 12208 14714
rect 12220 14662 12272 14714
rect 12284 14662 12336 14714
rect 12348 14662 12400 14714
rect 19520 14662 19572 14714
rect 19584 14662 19636 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 26948 14662 27000 14714
rect 27012 14662 27064 14714
rect 27076 14662 27128 14714
rect 27140 14662 27192 14714
rect 27204 14662 27256 14714
rect 5172 14560 5224 14612
rect 5908 14560 5960 14612
rect 6092 14560 6144 14612
rect 6552 14560 6604 14612
rect 5080 14492 5132 14544
rect 8300 14560 8352 14612
rect 9220 14560 9272 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 10968 14560 11020 14612
rect 13728 14560 13780 14612
rect 14280 14560 14332 14612
rect 16304 14560 16356 14612
rect 16580 14560 16632 14612
rect 16856 14560 16908 14612
rect 16948 14560 17000 14612
rect 19156 14560 19208 14612
rect 21916 14560 21968 14612
rect 22100 14560 22152 14612
rect 24492 14560 24544 14612
rect 25044 14560 25096 14612
rect 25320 14560 25372 14612
rect 25504 14560 25556 14612
rect 5632 14467 5684 14476
rect 5632 14433 5641 14467
rect 5641 14433 5675 14467
rect 5675 14433 5684 14467
rect 5632 14424 5684 14433
rect 3240 14356 3292 14408
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 5724 14399 5776 14408
rect 5724 14365 5733 14399
rect 5733 14365 5767 14399
rect 5767 14365 5776 14399
rect 5724 14356 5776 14365
rect 6460 14424 6512 14476
rect 7472 14492 7524 14544
rect 6092 14288 6144 14340
rect 940 14220 992 14272
rect 6276 14288 6328 14340
rect 8576 14492 8628 14544
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 6552 14220 6604 14272
rect 8116 14220 8168 14272
rect 9128 14424 9180 14476
rect 16028 14467 16080 14476
rect 12624 14356 12676 14408
rect 13452 14356 13504 14408
rect 16028 14433 16037 14467
rect 16037 14433 16071 14467
rect 16071 14433 16080 14467
rect 16028 14424 16080 14433
rect 14556 14356 14608 14408
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 18328 14492 18380 14544
rect 20444 14492 20496 14544
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 9220 14220 9272 14272
rect 10508 14220 10560 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 14188 14263 14240 14272
rect 14188 14229 14197 14263
rect 14197 14229 14231 14263
rect 14231 14229 14240 14263
rect 14188 14220 14240 14229
rect 17040 14220 17092 14272
rect 19432 14424 19484 14476
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 20720 14356 20772 14408
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 21272 14356 21324 14408
rect 19340 14288 19392 14340
rect 20812 14288 20864 14340
rect 21456 14288 21508 14340
rect 18788 14220 18840 14272
rect 18972 14263 19024 14272
rect 18972 14229 18981 14263
rect 18981 14229 19015 14263
rect 19015 14229 19024 14263
rect 18972 14220 19024 14229
rect 20720 14220 20772 14272
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 22376 14356 22428 14365
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 22744 14399 22796 14408
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 22284 14331 22336 14340
rect 22284 14297 22293 14331
rect 22293 14297 22327 14331
rect 22327 14297 22336 14331
rect 22284 14288 22336 14297
rect 25228 14424 25280 14476
rect 30380 14535 30432 14544
rect 30380 14501 30389 14535
rect 30389 14501 30423 14535
rect 30423 14501 30432 14535
rect 30380 14492 30432 14501
rect 30196 14399 30248 14408
rect 30196 14365 30205 14399
rect 30205 14365 30239 14399
rect 30239 14365 30248 14399
rect 30196 14356 30248 14365
rect 25872 14331 25924 14340
rect 25872 14297 25881 14331
rect 25881 14297 25915 14331
rect 25915 14297 25924 14331
rect 25872 14288 25924 14297
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 5324 14118 5376 14170
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 12752 14118 12804 14170
rect 12816 14118 12868 14170
rect 12880 14118 12932 14170
rect 12944 14118 12996 14170
rect 13008 14118 13060 14170
rect 20180 14118 20232 14170
rect 20244 14118 20296 14170
rect 20308 14118 20360 14170
rect 20372 14118 20424 14170
rect 20436 14118 20488 14170
rect 27608 14118 27660 14170
rect 27672 14118 27724 14170
rect 27736 14118 27788 14170
rect 27800 14118 27852 14170
rect 27864 14118 27916 14170
rect 5172 14016 5224 14068
rect 4252 13948 4304 14000
rect 4620 13948 4672 14000
rect 5724 14016 5776 14068
rect 6184 14016 6236 14068
rect 6368 14016 6420 14068
rect 8208 14016 8260 14068
rect 9312 14016 9364 14068
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 6092 13948 6144 14000
rect 6460 13948 6512 14000
rect 8668 13948 8720 14000
rect 9128 13948 9180 14000
rect 6276 13880 6328 13932
rect 10508 13948 10560 14000
rect 4988 13855 5040 13864
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 14188 14016 14240 14068
rect 14280 14016 14332 14068
rect 14740 14016 14792 14068
rect 15752 14016 15804 14068
rect 17316 14016 17368 14068
rect 17592 14059 17644 14068
rect 12348 13948 12400 14000
rect 15476 13880 15528 13932
rect 17592 14025 17601 14059
rect 17601 14025 17635 14059
rect 17635 14025 17644 14059
rect 17592 14016 17644 14025
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 18972 14016 19024 14068
rect 20536 14016 20588 14068
rect 18788 13991 18840 14000
rect 18788 13957 18797 13991
rect 18797 13957 18831 13991
rect 18831 13957 18840 13991
rect 18788 13948 18840 13957
rect 18236 13880 18288 13932
rect 18880 13880 18932 13932
rect 4988 13812 5040 13821
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 16028 13812 16080 13864
rect 18788 13812 18840 13864
rect 20812 13948 20864 14000
rect 22652 14016 22704 14068
rect 24400 14016 24452 14068
rect 25320 14016 25372 14068
rect 22744 13948 22796 14000
rect 22928 13948 22980 14000
rect 22100 13880 22152 13932
rect 25136 13948 25188 14000
rect 24768 13923 24820 13932
rect 24768 13889 24777 13923
rect 24777 13889 24811 13923
rect 24811 13889 24820 13923
rect 24768 13880 24820 13889
rect 19432 13787 19484 13796
rect 19432 13753 19441 13787
rect 19441 13753 19475 13787
rect 19475 13753 19484 13787
rect 19432 13744 19484 13753
rect 24492 13812 24544 13864
rect 30196 13812 30248 13864
rect 30288 13812 30340 13864
rect 1676 13676 1728 13728
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 8116 13719 8168 13728
rect 8116 13685 8125 13719
rect 8125 13685 8159 13719
rect 8159 13685 8168 13719
rect 8116 13676 8168 13685
rect 11612 13676 11664 13728
rect 13268 13719 13320 13728
rect 13268 13685 13277 13719
rect 13277 13685 13311 13719
rect 13311 13685 13320 13719
rect 13268 13676 13320 13685
rect 14648 13676 14700 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 19156 13719 19208 13728
rect 19156 13685 19165 13719
rect 19165 13685 19199 13719
rect 19199 13685 19208 13719
rect 19156 13676 19208 13685
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 22284 13676 22336 13728
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 25228 13719 25280 13728
rect 25228 13685 25237 13719
rect 25237 13685 25271 13719
rect 25271 13685 25280 13719
rect 25228 13676 25280 13685
rect 29000 13676 29052 13728
rect 4664 13574 4716 13626
rect 4728 13574 4780 13626
rect 4792 13574 4844 13626
rect 4856 13574 4908 13626
rect 4920 13574 4972 13626
rect 12092 13574 12144 13626
rect 12156 13574 12208 13626
rect 12220 13574 12272 13626
rect 12284 13574 12336 13626
rect 12348 13574 12400 13626
rect 19520 13574 19572 13626
rect 19584 13574 19636 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 26948 13574 27000 13626
rect 27012 13574 27064 13626
rect 27076 13574 27128 13626
rect 27140 13574 27192 13626
rect 27204 13574 27256 13626
rect 4252 13515 4304 13524
rect 4252 13481 4261 13515
rect 4261 13481 4295 13515
rect 4295 13481 4304 13515
rect 4252 13472 4304 13481
rect 6276 13472 6328 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9772 13472 9824 13524
rect 10692 13472 10744 13524
rect 4068 13336 4120 13388
rect 6736 13336 6788 13388
rect 9036 13447 9088 13456
rect 9036 13413 9045 13447
rect 9045 13413 9079 13447
rect 9079 13413 9088 13447
rect 9036 13404 9088 13413
rect 11796 13472 11848 13524
rect 15476 13472 15528 13524
rect 16304 13472 16356 13524
rect 17132 13472 17184 13524
rect 8116 13336 8168 13388
rect 13544 13336 13596 13388
rect 21272 13404 21324 13456
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 6092 13268 6144 13320
rect 7012 13268 7064 13320
rect 7840 13268 7892 13320
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 6000 13243 6052 13252
rect 6000 13209 6009 13243
rect 6009 13209 6043 13243
rect 6043 13209 6052 13243
rect 6000 13200 6052 13209
rect 9404 13243 9456 13252
rect 9404 13209 9413 13243
rect 9413 13209 9447 13243
rect 9447 13209 9456 13243
rect 9404 13200 9456 13209
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 940 13132 992 13184
rect 4160 13132 4212 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 11428 13132 11480 13184
rect 13268 13268 13320 13320
rect 14556 13268 14608 13320
rect 14740 13268 14792 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 16120 13268 16172 13320
rect 19064 13336 19116 13388
rect 21916 13336 21968 13388
rect 22376 13336 22428 13388
rect 22652 13336 22704 13388
rect 23388 13336 23440 13388
rect 17316 13311 17368 13320
rect 17316 13277 17325 13311
rect 17325 13277 17359 13311
rect 17359 13277 17368 13311
rect 17316 13268 17368 13277
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 15384 13243 15436 13252
rect 15384 13209 15393 13243
rect 15393 13209 15427 13243
rect 15427 13209 15436 13243
rect 15384 13200 15436 13209
rect 17040 13200 17092 13252
rect 13084 13132 13136 13184
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 17132 13175 17184 13184
rect 17132 13141 17141 13175
rect 17141 13141 17175 13175
rect 17175 13141 17184 13175
rect 17132 13132 17184 13141
rect 17776 13200 17828 13252
rect 19156 13268 19208 13320
rect 18144 13200 18196 13252
rect 18972 13175 19024 13184
rect 18972 13141 18981 13175
rect 18981 13141 19015 13175
rect 19015 13141 19024 13175
rect 18972 13132 19024 13141
rect 20536 13200 20588 13252
rect 20996 13200 21048 13252
rect 20628 13132 20680 13184
rect 21824 13132 21876 13184
rect 22744 13268 22796 13320
rect 23020 13311 23072 13320
rect 23020 13277 23029 13311
rect 23029 13277 23063 13311
rect 23063 13277 23072 13311
rect 29000 13404 29052 13456
rect 25136 13336 25188 13388
rect 23020 13268 23072 13277
rect 24492 13268 24544 13320
rect 24676 13311 24728 13320
rect 24676 13277 24685 13311
rect 24685 13277 24719 13311
rect 24719 13277 24728 13311
rect 24676 13268 24728 13277
rect 25872 13268 25924 13320
rect 22284 13243 22336 13252
rect 22284 13209 22293 13243
rect 22293 13209 22327 13243
rect 22327 13209 22336 13243
rect 22284 13200 22336 13209
rect 22560 13132 22612 13184
rect 22652 13175 22704 13184
rect 22652 13141 22661 13175
rect 22661 13141 22695 13175
rect 22695 13141 22704 13175
rect 22652 13132 22704 13141
rect 24492 13175 24544 13184
rect 24492 13141 24501 13175
rect 24501 13141 24535 13175
rect 24535 13141 24544 13175
rect 24492 13132 24544 13141
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 30380 13175 30432 13184
rect 30380 13141 30389 13175
rect 30389 13141 30423 13175
rect 30423 13141 30432 13175
rect 30380 13132 30432 13141
rect 5324 13030 5376 13082
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 12752 13030 12804 13082
rect 12816 13030 12868 13082
rect 12880 13030 12932 13082
rect 12944 13030 12996 13082
rect 13008 13030 13060 13082
rect 20180 13030 20232 13082
rect 20244 13030 20296 13082
rect 20308 13030 20360 13082
rect 20372 13030 20424 13082
rect 20436 13030 20488 13082
rect 27608 13030 27660 13082
rect 27672 13030 27724 13082
rect 27736 13030 27788 13082
rect 27800 13030 27852 13082
rect 27864 13030 27916 13082
rect 4068 12928 4120 12980
rect 4344 12928 4396 12980
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 6092 12928 6144 12980
rect 6368 12928 6420 12980
rect 6736 12928 6788 12980
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 5816 12792 5868 12844
rect 6276 12792 6328 12844
rect 6460 12792 6512 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 10508 12928 10560 12980
rect 11428 12928 11480 12980
rect 13360 12928 13412 12980
rect 8300 12860 8352 12912
rect 9404 12860 9456 12912
rect 10416 12903 10468 12912
rect 10416 12869 10425 12903
rect 10425 12869 10459 12903
rect 10459 12869 10468 12903
rect 10416 12860 10468 12869
rect 8392 12792 8444 12844
rect 7932 12724 7984 12776
rect 7748 12656 7800 12708
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 6092 12588 6144 12640
rect 6276 12588 6328 12640
rect 7472 12588 7524 12640
rect 8116 12588 8168 12640
rect 8668 12588 8720 12640
rect 11152 12724 11204 12776
rect 11612 12792 11664 12844
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 14648 12860 14700 12912
rect 15936 12928 15988 12980
rect 16028 12928 16080 12980
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 14004 12724 14056 12776
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15108 12792 15160 12844
rect 14556 12724 14608 12776
rect 16948 12860 17000 12912
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 18604 12928 18656 12980
rect 18972 12928 19024 12980
rect 19432 12928 19484 12980
rect 20536 12971 20588 12980
rect 20536 12937 20545 12971
rect 20545 12937 20579 12971
rect 20579 12937 20588 12971
rect 20536 12928 20588 12937
rect 18052 12792 18104 12844
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 21824 12928 21876 12980
rect 22652 12928 22704 12980
rect 23020 12928 23072 12980
rect 23388 12928 23440 12980
rect 24492 12928 24544 12980
rect 24952 12971 25004 12980
rect 24952 12937 24961 12971
rect 24961 12937 24995 12971
rect 24995 12937 25004 12971
rect 24952 12928 25004 12937
rect 25320 12928 25372 12980
rect 30196 12928 30248 12980
rect 22192 12903 22244 12912
rect 22192 12869 22201 12903
rect 22201 12869 22235 12903
rect 22235 12869 22244 12903
rect 22192 12860 22244 12869
rect 22560 12860 22612 12912
rect 9128 12656 9180 12708
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 10968 12656 11020 12708
rect 19340 12724 19392 12776
rect 21088 12724 21140 12776
rect 22468 12792 22520 12844
rect 22560 12724 22612 12776
rect 22928 12724 22980 12776
rect 19432 12656 19484 12708
rect 20076 12656 20128 12708
rect 20812 12656 20864 12708
rect 21180 12656 21232 12708
rect 24860 12835 24912 12844
rect 24860 12801 24869 12835
rect 24869 12801 24903 12835
rect 24903 12801 24912 12835
rect 24860 12792 24912 12801
rect 25688 12792 25740 12844
rect 30288 12792 30340 12844
rect 24676 12724 24728 12776
rect 25872 12724 25924 12776
rect 11060 12588 11112 12640
rect 11336 12588 11388 12640
rect 11980 12631 12032 12640
rect 11980 12597 11989 12631
rect 11989 12597 12023 12631
rect 12023 12597 12032 12631
rect 11980 12588 12032 12597
rect 12900 12588 12952 12640
rect 13360 12588 13412 12640
rect 16304 12588 16356 12640
rect 18144 12588 18196 12640
rect 18696 12588 18748 12640
rect 19156 12588 19208 12640
rect 22284 12588 22336 12640
rect 22376 12588 22428 12640
rect 23020 12588 23072 12640
rect 25044 12588 25096 12640
rect 4664 12486 4716 12538
rect 4728 12486 4780 12538
rect 4792 12486 4844 12538
rect 4856 12486 4908 12538
rect 4920 12486 4972 12538
rect 12092 12486 12144 12538
rect 12156 12486 12208 12538
rect 12220 12486 12272 12538
rect 12284 12486 12336 12538
rect 12348 12486 12400 12538
rect 19520 12486 19572 12538
rect 19584 12486 19636 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 26948 12486 27000 12538
rect 27012 12486 27064 12538
rect 27076 12486 27128 12538
rect 27140 12486 27192 12538
rect 27204 12486 27256 12538
rect 6368 12427 6420 12436
rect 6368 12393 6377 12427
rect 6377 12393 6411 12427
rect 6411 12393 6420 12427
rect 6368 12384 6420 12393
rect 6644 12384 6696 12436
rect 7840 12316 7892 12368
rect 8300 12384 8352 12436
rect 8392 12384 8444 12436
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 10048 12384 10100 12436
rect 10416 12359 10468 12368
rect 10416 12325 10425 12359
rect 10425 12325 10459 12359
rect 10459 12325 10468 12359
rect 10416 12316 10468 12325
rect 3976 12248 4028 12300
rect 7012 12248 7064 12300
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 8208 12248 8260 12300
rect 9312 12248 9364 12300
rect 10968 12384 11020 12436
rect 11152 12427 11204 12436
rect 11152 12393 11161 12427
rect 11161 12393 11195 12427
rect 11195 12393 11204 12427
rect 11152 12384 11204 12393
rect 13084 12384 13136 12436
rect 13544 12427 13596 12436
rect 13544 12393 13553 12427
rect 13553 12393 13587 12427
rect 13587 12393 13596 12427
rect 13544 12384 13596 12393
rect 14464 12384 14516 12436
rect 16304 12384 16356 12436
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 17224 12384 17276 12436
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 5724 12180 5776 12232
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 6460 12180 6512 12232
rect 7564 12180 7616 12232
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 9680 12180 9732 12232
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10692 12180 10744 12232
rect 6828 12044 6880 12096
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 11336 12180 11388 12232
rect 11888 12180 11940 12232
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 12900 12112 12952 12164
rect 10324 12044 10376 12096
rect 10692 12087 10744 12096
rect 10692 12053 10719 12087
rect 10719 12053 10744 12087
rect 10692 12044 10744 12053
rect 11612 12044 11664 12096
rect 11980 12044 12032 12096
rect 18052 12316 18104 12368
rect 20996 12427 21048 12436
rect 20996 12393 21005 12427
rect 21005 12393 21039 12427
rect 21039 12393 21048 12427
rect 20996 12384 21048 12393
rect 25044 12384 25096 12436
rect 13636 12180 13688 12232
rect 13820 12223 13872 12232
rect 13820 12189 13829 12223
rect 13829 12189 13863 12223
rect 13863 12189 13872 12223
rect 13820 12180 13872 12189
rect 14648 12180 14700 12232
rect 18880 12248 18932 12300
rect 19340 12291 19392 12300
rect 19340 12257 19349 12291
rect 19349 12257 19383 12291
rect 19383 12257 19392 12291
rect 19340 12248 19392 12257
rect 17408 12180 17460 12232
rect 17040 12112 17092 12164
rect 17868 12112 17920 12164
rect 13912 12044 13964 12096
rect 16304 12044 16356 12096
rect 17224 12044 17276 12096
rect 20444 12112 20496 12164
rect 18512 12044 18564 12096
rect 19340 12044 19392 12096
rect 19892 12044 19944 12096
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 24860 12316 24912 12368
rect 21180 12223 21232 12232
rect 21180 12189 21189 12223
rect 21189 12189 21223 12223
rect 21223 12189 21232 12223
rect 21180 12180 21232 12189
rect 21272 12180 21324 12232
rect 22928 12180 22980 12232
rect 25320 12180 25372 12232
rect 24032 12155 24084 12164
rect 24032 12121 24041 12155
rect 24041 12121 24075 12155
rect 24075 12121 24084 12155
rect 24032 12112 24084 12121
rect 24952 12155 25004 12164
rect 24952 12121 24961 12155
rect 24961 12121 24995 12155
rect 24995 12121 25004 12155
rect 24952 12112 25004 12121
rect 25320 12087 25372 12096
rect 25320 12053 25329 12087
rect 25329 12053 25363 12087
rect 25363 12053 25372 12087
rect 25320 12044 25372 12053
rect 25688 12155 25740 12164
rect 25688 12121 25697 12155
rect 25697 12121 25731 12155
rect 25731 12121 25740 12155
rect 25688 12112 25740 12121
rect 5324 11942 5376 11994
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 12752 11942 12804 11994
rect 12816 11942 12868 11994
rect 12880 11942 12932 11994
rect 12944 11942 12996 11994
rect 13008 11942 13060 11994
rect 20180 11942 20232 11994
rect 20244 11942 20296 11994
rect 20308 11942 20360 11994
rect 20372 11942 20424 11994
rect 20436 11942 20488 11994
rect 27608 11942 27660 11994
rect 27672 11942 27724 11994
rect 27736 11942 27788 11994
rect 27800 11942 27852 11994
rect 27864 11942 27916 11994
rect 940 11704 992 11756
rect 4988 11840 5040 11892
rect 7564 11840 7616 11892
rect 8392 11840 8444 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 11612 11840 11664 11892
rect 13084 11840 13136 11892
rect 13544 11840 13596 11892
rect 17684 11840 17736 11892
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 4252 11772 4304 11824
rect 4528 11704 4580 11756
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 4436 11636 4488 11688
rect 4344 11568 4396 11620
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 7748 11704 7800 11756
rect 7288 11568 7340 11620
rect 3976 11500 4028 11552
rect 4528 11500 4580 11552
rect 5264 11500 5316 11552
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 6092 11543 6144 11552
rect 6092 11509 6101 11543
rect 6101 11509 6135 11543
rect 6135 11509 6144 11543
rect 6092 11500 6144 11509
rect 6276 11500 6328 11552
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 8392 11704 8444 11756
rect 8576 11772 8628 11824
rect 9588 11772 9640 11824
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 8760 11636 8812 11688
rect 10784 11704 10836 11756
rect 14004 11772 14056 11824
rect 18328 11772 18380 11824
rect 18512 11772 18564 11824
rect 19248 11883 19300 11892
rect 19248 11849 19257 11883
rect 19257 11849 19291 11883
rect 19291 11849 19300 11883
rect 19248 11840 19300 11849
rect 22652 11840 22704 11892
rect 10692 11636 10744 11688
rect 11980 11636 12032 11688
rect 9220 11568 9272 11620
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 17040 11704 17092 11756
rect 17684 11704 17736 11756
rect 15384 11636 15436 11645
rect 16396 11568 16448 11620
rect 9956 11500 10008 11552
rect 13544 11500 13596 11552
rect 16488 11500 16540 11552
rect 18420 11704 18472 11756
rect 18880 11704 18932 11756
rect 18788 11636 18840 11688
rect 19524 11704 19576 11756
rect 19892 11772 19944 11824
rect 20996 11772 21048 11824
rect 21640 11704 21692 11756
rect 22928 11840 22980 11892
rect 24032 11840 24084 11892
rect 25320 11840 25372 11892
rect 19064 11636 19116 11688
rect 19340 11568 19392 11620
rect 20076 11636 20128 11688
rect 22560 11636 22612 11688
rect 22928 11679 22980 11688
rect 22928 11645 22937 11679
rect 22937 11645 22971 11679
rect 22971 11645 22980 11679
rect 22928 11636 22980 11645
rect 17224 11500 17276 11552
rect 18788 11543 18840 11552
rect 18788 11509 18812 11543
rect 18812 11509 18840 11543
rect 18788 11500 18840 11509
rect 18880 11543 18932 11552
rect 18880 11509 18889 11543
rect 18889 11509 18923 11543
rect 18923 11509 18932 11543
rect 18880 11500 18932 11509
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 19524 11500 19576 11552
rect 20720 11568 20772 11620
rect 23940 11704 23992 11756
rect 24400 11704 24452 11756
rect 24492 11747 24544 11756
rect 24492 11713 24501 11747
rect 24501 11713 24535 11747
rect 24535 11713 24544 11747
rect 24492 11704 24544 11713
rect 24032 11679 24084 11688
rect 24032 11645 24041 11679
rect 24041 11645 24075 11679
rect 24075 11645 24084 11679
rect 24032 11636 24084 11645
rect 24768 11704 24820 11756
rect 25228 11704 25280 11756
rect 25688 11636 25740 11688
rect 22008 11543 22060 11552
rect 22008 11509 22032 11543
rect 22032 11509 22060 11543
rect 22008 11500 22060 11509
rect 22192 11500 22244 11552
rect 23112 11500 23164 11552
rect 23756 11568 23808 11620
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 26148 11636 26200 11688
rect 25688 11500 25740 11552
rect 30380 11611 30432 11620
rect 30380 11577 30389 11611
rect 30389 11577 30423 11611
rect 30423 11577 30432 11611
rect 30380 11568 30432 11577
rect 4664 11398 4716 11450
rect 4728 11398 4780 11450
rect 4792 11398 4844 11450
rect 4856 11398 4908 11450
rect 4920 11398 4972 11450
rect 12092 11398 12144 11450
rect 12156 11398 12208 11450
rect 12220 11398 12272 11450
rect 12284 11398 12336 11450
rect 12348 11398 12400 11450
rect 19520 11398 19572 11450
rect 19584 11398 19636 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 26948 11398 27000 11450
rect 27012 11398 27064 11450
rect 27076 11398 27128 11450
rect 27140 11398 27192 11450
rect 27204 11398 27256 11450
rect 3240 11296 3292 11348
rect 4252 11296 4304 11348
rect 4344 11296 4396 11348
rect 4528 11296 4580 11348
rect 6276 11339 6328 11348
rect 6276 11305 6285 11339
rect 6285 11305 6319 11339
rect 6319 11305 6328 11339
rect 6276 11296 6328 11305
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8392 11296 8444 11348
rect 9312 11296 9364 11348
rect 13544 11296 13596 11348
rect 15384 11296 15436 11348
rect 4252 11135 4304 11144
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4436 11024 4488 11076
rect 5264 11092 5316 11144
rect 6092 11092 6144 11144
rect 6368 11135 6420 11144
rect 6368 11101 6377 11135
rect 6377 11101 6411 11135
rect 6411 11101 6420 11135
rect 6368 11092 6420 11101
rect 7104 11135 7156 11144
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 7748 11092 7800 11144
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 11336 11228 11388 11280
rect 13820 11228 13872 11280
rect 17592 11296 17644 11348
rect 19064 11296 19116 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 22928 11296 22980 11348
rect 23112 11296 23164 11348
rect 23940 11296 23992 11348
rect 24768 11296 24820 11348
rect 27620 11296 27672 11348
rect 25228 11228 25280 11280
rect 25412 11228 25464 11280
rect 16488 11160 16540 11212
rect 6920 11024 6972 11076
rect 11152 11092 11204 11144
rect 11612 11092 11664 11144
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 6736 10956 6788 11008
rect 8208 10956 8260 11008
rect 9864 11024 9916 11076
rect 11428 11024 11480 11076
rect 11060 10956 11112 11008
rect 12072 11024 12124 11076
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 15108 11024 15160 11076
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 19432 11160 19484 11212
rect 21824 11160 21876 11212
rect 18788 11092 18840 11144
rect 18880 11092 18932 11144
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 21916 11024 21968 11076
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 23940 11092 23992 11144
rect 24492 11135 24544 11144
rect 24492 11101 24501 11135
rect 24501 11101 24535 11135
rect 24535 11101 24544 11135
rect 24492 11092 24544 11101
rect 24768 11092 24820 11144
rect 25688 11203 25740 11212
rect 25688 11169 25697 11203
rect 25697 11169 25731 11203
rect 25731 11169 25740 11203
rect 25688 11160 25740 11169
rect 30288 11092 30340 11144
rect 11704 10956 11756 11008
rect 13268 10956 13320 11008
rect 13636 10999 13688 11008
rect 13636 10965 13645 10999
rect 13645 10965 13679 10999
rect 13679 10965 13688 10999
rect 13636 10956 13688 10965
rect 23664 11024 23716 11076
rect 23020 10956 23072 11008
rect 26240 11024 26292 11076
rect 5324 10854 5376 10906
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 12752 10854 12804 10906
rect 12816 10854 12868 10906
rect 12880 10854 12932 10906
rect 12944 10854 12996 10906
rect 13008 10854 13060 10906
rect 20180 10854 20232 10906
rect 20244 10854 20296 10906
rect 20308 10854 20360 10906
rect 20372 10854 20424 10906
rect 20436 10854 20488 10906
rect 27608 10854 27660 10906
rect 27672 10854 27724 10906
rect 27736 10854 27788 10906
rect 27800 10854 27852 10906
rect 27864 10854 27916 10906
rect 6368 10752 6420 10804
rect 6920 10752 6972 10804
rect 8300 10752 8352 10804
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 4528 10616 4580 10668
rect 6736 10684 6788 10736
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 11152 10752 11204 10804
rect 15108 10752 15160 10804
rect 18420 10752 18472 10804
rect 20904 10752 20956 10804
rect 22008 10752 22060 10804
rect 7104 10548 7156 10600
rect 8116 10548 8168 10600
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9772 10616 9824 10668
rect 10140 10616 10192 10668
rect 10416 10684 10468 10736
rect 10324 10659 10376 10668
rect 10324 10625 10333 10659
rect 10333 10625 10367 10659
rect 10367 10625 10376 10659
rect 10324 10616 10376 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11428 10684 11480 10736
rect 11060 10659 11112 10668
rect 11060 10625 11069 10659
rect 11069 10625 11103 10659
rect 11103 10625 11112 10659
rect 11060 10616 11112 10625
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 11612 10616 11664 10668
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 13636 10684 13688 10736
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 13268 10616 13320 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 15752 10616 15804 10668
rect 17408 10616 17460 10668
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 21364 10684 21416 10736
rect 17960 10616 18012 10625
rect 6184 10480 6236 10532
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 940 10412 992 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 8852 10412 8904 10464
rect 9588 10412 9640 10464
rect 11704 10480 11756 10532
rect 11980 10480 12032 10532
rect 13544 10523 13596 10532
rect 13544 10489 13553 10523
rect 13553 10489 13587 10523
rect 13587 10489 13596 10523
rect 13544 10480 13596 10489
rect 14004 10480 14056 10532
rect 18788 10548 18840 10600
rect 11612 10412 11664 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 19984 10412 20036 10464
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 21732 10616 21784 10668
rect 22928 10752 22980 10804
rect 26240 10795 26292 10804
rect 26240 10761 26249 10795
rect 26249 10761 26283 10795
rect 26283 10761 26292 10795
rect 26240 10752 26292 10761
rect 21088 10548 21140 10600
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 23664 10684 23716 10736
rect 24124 10684 24176 10736
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 20812 10480 20864 10532
rect 20720 10412 20772 10464
rect 21364 10412 21416 10464
rect 21916 10480 21968 10532
rect 24032 10548 24084 10600
rect 24860 10616 24912 10668
rect 30932 10616 30984 10668
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 21640 10412 21692 10421
rect 21732 10412 21784 10464
rect 23020 10412 23072 10464
rect 23480 10480 23532 10532
rect 23572 10480 23624 10532
rect 23756 10480 23808 10532
rect 24400 10480 24452 10532
rect 23940 10412 23992 10464
rect 25136 10412 25188 10464
rect 4664 10310 4716 10362
rect 4728 10310 4780 10362
rect 4792 10310 4844 10362
rect 4856 10310 4908 10362
rect 4920 10310 4972 10362
rect 12092 10310 12144 10362
rect 12156 10310 12208 10362
rect 12220 10310 12272 10362
rect 12284 10310 12336 10362
rect 12348 10310 12400 10362
rect 19520 10310 19572 10362
rect 19584 10310 19636 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 26948 10310 27000 10362
rect 27012 10310 27064 10362
rect 27076 10310 27128 10362
rect 27140 10310 27192 10362
rect 27204 10310 27256 10362
rect 6920 10208 6972 10260
rect 8944 10208 8996 10260
rect 10600 10208 10652 10260
rect 11520 10208 11572 10260
rect 8208 10140 8260 10192
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 6184 10072 6236 10124
rect 7840 10072 7892 10124
rect 12624 10140 12676 10192
rect 18236 10208 18288 10260
rect 18788 10208 18840 10260
rect 19340 10208 19392 10260
rect 21548 10208 21600 10260
rect 23204 10208 23256 10260
rect 4988 10004 5040 10056
rect 6644 10004 6696 10056
rect 6736 10004 6788 10056
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 5908 9936 5960 9988
rect 7564 9979 7616 9988
rect 7564 9945 7573 9979
rect 7573 9945 7607 9979
rect 7607 9945 7616 9979
rect 7564 9936 7616 9945
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 8116 9936 8168 9988
rect 8392 9936 8444 9988
rect 9496 10004 9548 10056
rect 9588 10047 9640 10056
rect 9588 10013 9597 10047
rect 9597 10013 9631 10047
rect 9631 10013 9640 10047
rect 9588 10004 9640 10013
rect 9956 10047 10008 10056
rect 9956 10013 9965 10047
rect 9965 10013 9999 10047
rect 9999 10013 10008 10047
rect 9956 10004 10008 10013
rect 10416 10004 10468 10056
rect 11244 10004 11296 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 11704 10004 11756 10056
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 5172 9868 5224 9920
rect 5724 9868 5776 9920
rect 7472 9868 7524 9920
rect 11796 9868 11848 9920
rect 15476 10004 15528 10056
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 14372 9979 14424 9988
rect 14372 9945 14381 9979
rect 14381 9945 14415 9979
rect 14415 9945 14424 9979
rect 14372 9936 14424 9945
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 12624 9868 12676 9920
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 15936 9911 15988 9920
rect 15936 9877 15945 9911
rect 15945 9877 15979 9911
rect 15979 9877 15988 9911
rect 15936 9868 15988 9877
rect 17132 9868 17184 9920
rect 17408 9868 17460 9920
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 20076 10140 20128 10192
rect 20168 10140 20220 10192
rect 20628 10140 20680 10192
rect 21456 10140 21508 10192
rect 23572 10251 23624 10260
rect 23572 10217 23581 10251
rect 23581 10217 23615 10251
rect 23615 10217 23624 10251
rect 23572 10208 23624 10217
rect 23756 10208 23808 10260
rect 23940 10208 23992 10260
rect 19800 10115 19852 10124
rect 19800 10081 19809 10115
rect 19809 10081 19843 10115
rect 19843 10081 19852 10115
rect 19800 10072 19852 10081
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 24952 10140 25004 10192
rect 17684 9868 17736 9920
rect 18144 9868 18196 9920
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 20444 9936 20496 9988
rect 20536 9936 20588 9988
rect 20904 10004 20956 10056
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 22376 10004 22428 10056
rect 22560 10004 22612 10056
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 25320 10115 25372 10124
rect 25320 10081 25329 10115
rect 25329 10081 25363 10115
rect 25363 10081 25372 10115
rect 25320 10072 25372 10081
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 25136 10047 25188 10056
rect 25136 10013 25145 10047
rect 25145 10013 25179 10047
rect 25179 10013 25188 10047
rect 25136 10004 25188 10013
rect 25412 10004 25464 10056
rect 23204 9936 23256 9988
rect 23756 9936 23808 9988
rect 20996 9868 21048 9920
rect 22100 9868 22152 9920
rect 24492 9911 24544 9920
rect 24492 9877 24501 9911
rect 24501 9877 24535 9911
rect 24535 9877 24544 9911
rect 24492 9868 24544 9877
rect 30288 10004 30340 10056
rect 5324 9766 5376 9818
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 12752 9766 12804 9818
rect 12816 9766 12868 9818
rect 12880 9766 12932 9818
rect 12944 9766 12996 9818
rect 13008 9766 13060 9818
rect 20180 9766 20232 9818
rect 20244 9766 20296 9818
rect 20308 9766 20360 9818
rect 20372 9766 20424 9818
rect 20436 9766 20488 9818
rect 27608 9766 27660 9818
rect 27672 9766 27724 9818
rect 27736 9766 27788 9818
rect 27800 9766 27852 9818
rect 27864 9766 27916 9818
rect 5172 9664 5224 9716
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 7564 9664 7616 9716
rect 4528 9596 4580 9648
rect 8116 9664 8168 9716
rect 10600 9707 10652 9716
rect 10600 9673 10609 9707
rect 10609 9673 10643 9707
rect 10643 9673 10652 9707
rect 10600 9664 10652 9673
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 4988 9460 5040 9512
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 6092 9460 6144 9512
rect 6368 9503 6420 9512
rect 6368 9469 6377 9503
rect 6377 9469 6411 9503
rect 6411 9469 6420 9503
rect 6368 9460 6420 9469
rect 6460 9460 6512 9512
rect 5632 9392 5684 9444
rect 6920 9528 6972 9580
rect 6828 9460 6880 9512
rect 7472 9528 7524 9580
rect 7840 9639 7892 9648
rect 7840 9605 7849 9639
rect 7849 9605 7883 9639
rect 7883 9605 7892 9639
rect 7840 9596 7892 9605
rect 8024 9528 8076 9580
rect 8300 9528 8352 9580
rect 11612 9596 11664 9648
rect 11888 9596 11940 9648
rect 12900 9596 12952 9648
rect 13360 9596 13412 9648
rect 15936 9596 15988 9648
rect 16212 9664 16264 9716
rect 18052 9664 18104 9716
rect 19892 9707 19944 9716
rect 19892 9673 19901 9707
rect 19901 9673 19935 9707
rect 19935 9673 19944 9707
rect 19892 9664 19944 9673
rect 17316 9596 17368 9648
rect 8668 9460 8720 9512
rect 10692 9460 10744 9512
rect 11428 9528 11480 9580
rect 13084 9528 13136 9580
rect 14096 9528 14148 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 15476 9528 15528 9580
rect 15752 9528 15804 9580
rect 16948 9528 17000 9580
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 17776 9639 17828 9648
rect 17776 9605 17785 9639
rect 17785 9605 17819 9639
rect 17819 9605 17828 9639
rect 17776 9596 17828 9605
rect 20260 9596 20312 9648
rect 13176 9460 13228 9512
rect 14372 9460 14424 9512
rect 9772 9392 9824 9444
rect 13452 9392 13504 9444
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 19708 9528 19760 9580
rect 20996 9664 21048 9716
rect 22284 9664 22336 9716
rect 22376 9707 22428 9716
rect 22376 9673 22385 9707
rect 22385 9673 22419 9707
rect 22419 9673 22428 9707
rect 22376 9664 22428 9673
rect 24400 9596 24452 9648
rect 20536 9528 20588 9580
rect 18328 9460 18380 9512
rect 21916 9460 21968 9512
rect 18972 9392 19024 9444
rect 19432 9392 19484 9444
rect 21824 9392 21876 9444
rect 23388 9503 23440 9512
rect 23388 9469 23397 9503
rect 23397 9469 23431 9503
rect 23431 9469 23440 9503
rect 23388 9460 23440 9469
rect 24952 9460 25004 9512
rect 25596 9503 25648 9512
rect 25596 9469 25605 9503
rect 25605 9469 25639 9503
rect 25639 9469 25648 9503
rect 25596 9460 25648 9469
rect 6276 9324 6328 9376
rect 10324 9324 10376 9376
rect 20168 9324 20220 9376
rect 21456 9324 21508 9376
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 23572 9324 23624 9376
rect 24952 9367 25004 9376
rect 24952 9333 24961 9367
rect 24961 9333 24995 9367
rect 24995 9333 25004 9367
rect 24952 9324 25004 9333
rect 4664 9222 4716 9274
rect 4728 9222 4780 9274
rect 4792 9222 4844 9274
rect 4856 9222 4908 9274
rect 4920 9222 4972 9274
rect 12092 9222 12144 9274
rect 12156 9222 12208 9274
rect 12220 9222 12272 9274
rect 12284 9222 12336 9274
rect 12348 9222 12400 9274
rect 19520 9222 19572 9274
rect 19584 9222 19636 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 26948 9222 27000 9274
rect 27012 9222 27064 9274
rect 27076 9222 27128 9274
rect 27140 9222 27192 9274
rect 27204 9222 27256 9274
rect 4436 9120 4488 9172
rect 4528 9120 4580 9172
rect 5908 9120 5960 9172
rect 6276 9120 6328 9172
rect 7380 9120 7432 9172
rect 7472 9120 7524 9172
rect 8760 9120 8812 9172
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 11428 9120 11480 9172
rect 17040 9120 17092 9172
rect 18328 9163 18380 9172
rect 18328 9129 18337 9163
rect 18337 9129 18371 9163
rect 18371 9129 18380 9163
rect 18328 9120 18380 9129
rect 18972 9120 19024 9172
rect 20812 9120 20864 9172
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 22284 9120 22336 9172
rect 22376 9120 22428 9172
rect 23388 9120 23440 9172
rect 23756 9163 23808 9172
rect 23756 9129 23765 9163
rect 23765 9129 23799 9163
rect 23799 9129 23808 9163
rect 23756 9120 23808 9129
rect 24492 9120 24544 9172
rect 24952 9120 25004 9172
rect 30380 9163 30432 9172
rect 30380 9129 30389 9163
rect 30389 9129 30423 9163
rect 30423 9129 30432 9163
rect 30380 9120 30432 9129
rect 6368 9052 6420 9104
rect 6828 9052 6880 9104
rect 9036 9052 9088 9104
rect 940 8916 992 8968
rect 4252 8916 4304 8968
rect 4988 8916 5040 8968
rect 6092 8984 6144 9036
rect 5172 8848 5224 8900
rect 5908 8848 5960 8900
rect 6644 8984 6696 9036
rect 9956 9052 10008 9104
rect 8484 8916 8536 8968
rect 9220 8916 9272 8968
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 9956 8916 10008 8968
rect 6092 8780 6144 8832
rect 9404 8891 9456 8900
rect 9404 8857 9413 8891
rect 9413 8857 9447 8891
rect 9447 8857 9456 8891
rect 9404 8848 9456 8857
rect 9496 8891 9548 8900
rect 9496 8857 9505 8891
rect 9505 8857 9539 8891
rect 9539 8857 9548 8891
rect 9496 8848 9548 8857
rect 9680 8848 9732 8900
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 11796 8916 11848 8968
rect 17132 9052 17184 9104
rect 17224 9052 17276 9104
rect 15660 8984 15712 9036
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 13360 8916 13412 8968
rect 7840 8780 7892 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 10416 8780 10468 8832
rect 10968 8780 11020 8832
rect 11244 8780 11296 8832
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 12624 8780 12676 8832
rect 13912 8959 13964 8968
rect 13912 8925 13921 8959
rect 13921 8925 13955 8959
rect 13955 8925 13964 8959
rect 13912 8916 13964 8925
rect 15200 8959 15252 8968
rect 15200 8925 15209 8959
rect 15209 8925 15243 8959
rect 15243 8925 15252 8959
rect 15200 8916 15252 8925
rect 15844 8916 15896 8968
rect 17316 8916 17368 8968
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 17500 8959 17552 8968
rect 17500 8925 17509 8959
rect 17509 8925 17543 8959
rect 17543 8925 17552 8959
rect 17500 8916 17552 8925
rect 18052 8984 18104 9036
rect 20536 9095 20588 9104
rect 20536 9061 20545 9095
rect 20545 9061 20579 9095
rect 20579 9061 20588 9095
rect 20536 9052 20588 9061
rect 20076 9027 20128 9036
rect 20076 8993 20085 9027
rect 20085 8993 20119 9027
rect 20119 8993 20128 9027
rect 20076 8984 20128 8993
rect 17132 8848 17184 8900
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 19432 8916 19484 8968
rect 18604 8848 18656 8900
rect 13452 8780 13504 8832
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 19432 8823 19484 8832
rect 19432 8789 19459 8823
rect 19459 8789 19484 8823
rect 19432 8780 19484 8789
rect 19892 8823 19944 8832
rect 19892 8789 19901 8823
rect 19901 8789 19935 8823
rect 19935 8789 19944 8823
rect 19892 8780 19944 8789
rect 20444 8916 20496 8968
rect 21640 9027 21692 9036
rect 21640 8993 21649 9027
rect 21649 8993 21683 9027
rect 21683 8993 21692 9027
rect 21640 8984 21692 8993
rect 23572 9052 23624 9104
rect 20168 8848 20220 8900
rect 23480 8959 23532 8968
rect 23480 8925 23489 8959
rect 23489 8925 23523 8959
rect 23523 8925 23532 8959
rect 23480 8916 23532 8925
rect 25596 8916 25648 8968
rect 5324 8678 5376 8730
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 12752 8678 12804 8730
rect 12816 8678 12868 8730
rect 12880 8678 12932 8730
rect 12944 8678 12996 8730
rect 13008 8678 13060 8730
rect 20180 8678 20232 8730
rect 20244 8678 20296 8730
rect 20308 8678 20360 8730
rect 20372 8678 20424 8730
rect 20436 8678 20488 8730
rect 27608 8678 27660 8730
rect 27672 8678 27724 8730
rect 27736 8678 27788 8730
rect 27800 8678 27852 8730
rect 27864 8678 27916 8730
rect 5908 8576 5960 8628
rect 7656 8576 7708 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 6552 8508 6604 8560
rect 9404 8576 9456 8628
rect 9496 8576 9548 8628
rect 6000 8372 6052 8424
rect 7472 8440 7524 8492
rect 7656 8483 7708 8492
rect 7656 8449 7681 8483
rect 7681 8449 7708 8483
rect 7656 8440 7708 8449
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 6736 8372 6788 8424
rect 9220 8508 9272 8560
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 8024 8440 8076 8492
rect 8300 8440 8352 8492
rect 9496 8440 9548 8492
rect 9680 8440 9732 8492
rect 10692 8576 10744 8628
rect 10968 8508 11020 8560
rect 13084 8576 13136 8628
rect 13176 8576 13228 8628
rect 15660 8576 15712 8628
rect 16304 8576 16356 8628
rect 17500 8576 17552 8628
rect 19892 8576 19944 8628
rect 20536 8576 20588 8628
rect 20812 8619 20864 8628
rect 20812 8585 20821 8619
rect 20821 8585 20855 8619
rect 20855 8585 20864 8619
rect 20812 8576 20864 8585
rect 21640 8576 21692 8628
rect 24400 8576 24452 8628
rect 13912 8508 13964 8560
rect 8484 8372 8536 8424
rect 6092 8236 6144 8288
rect 8392 8304 8444 8356
rect 9588 8372 9640 8424
rect 9956 8415 10008 8424
rect 9956 8381 9965 8415
rect 9965 8381 9999 8415
rect 9999 8381 10008 8415
rect 9956 8372 10008 8381
rect 11244 8440 11296 8492
rect 7104 8279 7156 8288
rect 7104 8245 7113 8279
rect 7113 8245 7147 8279
rect 7147 8245 7156 8279
rect 7104 8236 7156 8245
rect 7380 8236 7432 8288
rect 9036 8236 9088 8288
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 9312 8236 9364 8288
rect 10416 8304 10468 8356
rect 13452 8440 13504 8492
rect 17224 8440 17276 8492
rect 12624 8372 12676 8424
rect 17868 8440 17920 8492
rect 17960 8440 18012 8492
rect 17408 8372 17460 8424
rect 20628 8372 20680 8424
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 22100 8551 22152 8560
rect 22100 8517 22109 8551
rect 22109 8517 22143 8551
rect 22143 8517 22152 8551
rect 22100 8508 22152 8517
rect 23112 8508 23164 8560
rect 23664 8440 23716 8492
rect 24860 8440 24912 8492
rect 21088 8372 21140 8424
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 22192 8372 22244 8424
rect 23572 8415 23624 8424
rect 23572 8381 23581 8415
rect 23581 8381 23615 8415
rect 23615 8381 23624 8415
rect 23572 8372 23624 8381
rect 30288 8304 30340 8356
rect 19984 8236 20036 8288
rect 4664 8134 4716 8186
rect 4728 8134 4780 8186
rect 4792 8134 4844 8186
rect 4856 8134 4908 8186
rect 4920 8134 4972 8186
rect 12092 8134 12144 8186
rect 12156 8134 12208 8186
rect 12220 8134 12272 8186
rect 12284 8134 12336 8186
rect 12348 8134 12400 8186
rect 19520 8134 19572 8186
rect 19584 8134 19636 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 26948 8134 27000 8186
rect 27012 8134 27064 8186
rect 27076 8134 27128 8186
rect 27140 8134 27192 8186
rect 27204 8134 27256 8186
rect 6368 8032 6420 8084
rect 6552 8032 6604 8084
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 17592 8032 17644 8084
rect 7104 7896 7156 7948
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 5724 7760 5776 7812
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7840 7964 7892 8016
rect 18604 8032 18656 8084
rect 19340 7964 19392 8016
rect 21180 8032 21232 8084
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 21456 8032 21508 8084
rect 22192 8075 22244 8084
rect 22192 8041 22201 8075
rect 22201 8041 22235 8075
rect 22235 8041 22244 8075
rect 22192 8032 22244 8041
rect 23112 8032 23164 8084
rect 12532 7896 12584 7948
rect 13084 7896 13136 7948
rect 16580 7896 16632 7948
rect 17960 7896 18012 7948
rect 17684 7828 17736 7880
rect 17868 7871 17920 7880
rect 17868 7837 17877 7871
rect 17877 7837 17911 7871
rect 17911 7837 17920 7871
rect 17868 7828 17920 7837
rect 18420 7828 18472 7880
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 20996 7828 21048 7880
rect 21916 7964 21968 8016
rect 18236 7760 18288 7812
rect 940 7692 992 7744
rect 6368 7692 6420 7744
rect 11980 7692 12032 7744
rect 12624 7692 12676 7744
rect 17040 7692 17092 7744
rect 19432 7692 19484 7744
rect 21364 7692 21416 7744
rect 21916 7692 21968 7744
rect 22284 7692 22336 7744
rect 23664 7828 23716 7880
rect 5324 7590 5376 7642
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 12752 7590 12804 7642
rect 12816 7590 12868 7642
rect 12880 7590 12932 7642
rect 12944 7590 12996 7642
rect 13008 7590 13060 7642
rect 20180 7590 20232 7642
rect 20244 7590 20296 7642
rect 20308 7590 20360 7642
rect 20372 7590 20424 7642
rect 20436 7590 20488 7642
rect 27608 7590 27660 7642
rect 27672 7590 27724 7642
rect 27736 7590 27788 7642
rect 27800 7590 27852 7642
rect 27864 7590 27916 7642
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 6460 7488 6512 7540
rect 6368 7420 6420 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 5172 7352 5224 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 11520 7488 11572 7540
rect 12440 7488 12492 7540
rect 12624 7488 12676 7540
rect 17040 7420 17092 7472
rect 19432 7420 19484 7472
rect 20076 7420 20128 7472
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12440 7284 12492 7336
rect 18052 7352 18104 7404
rect 21088 7284 21140 7336
rect 10416 7148 10468 7200
rect 18420 7191 18472 7200
rect 18420 7157 18429 7191
rect 18429 7157 18463 7191
rect 18463 7157 18472 7191
rect 18420 7148 18472 7157
rect 20996 7148 21048 7200
rect 4664 7046 4716 7098
rect 4728 7046 4780 7098
rect 4792 7046 4844 7098
rect 4856 7046 4908 7098
rect 4920 7046 4972 7098
rect 12092 7046 12144 7098
rect 12156 7046 12208 7098
rect 12220 7046 12272 7098
rect 12284 7046 12336 7098
rect 12348 7046 12400 7098
rect 19520 7046 19572 7098
rect 19584 7046 19636 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 26948 7046 27000 7098
rect 27012 7046 27064 7098
rect 27076 7046 27128 7098
rect 27140 7046 27192 7098
rect 27204 7046 27256 7098
rect 8300 6944 8352 6996
rect 11796 6944 11848 6996
rect 20076 6987 20128 6996
rect 20076 6953 20085 6987
rect 20085 6953 20119 6987
rect 20119 6953 20128 6987
rect 20076 6944 20128 6953
rect 9128 6808 9180 6860
rect 13084 6808 13136 6860
rect 18052 6808 18104 6860
rect 10416 6740 10468 6792
rect 11980 6740 12032 6792
rect 16948 6740 17000 6792
rect 22284 6740 22336 6792
rect 5324 6502 5376 6554
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 12752 6502 12804 6554
rect 12816 6502 12868 6554
rect 12880 6502 12932 6554
rect 12944 6502 12996 6554
rect 13008 6502 13060 6554
rect 20180 6502 20232 6554
rect 20244 6502 20296 6554
rect 20308 6502 20360 6554
rect 20372 6502 20424 6554
rect 20436 6502 20488 6554
rect 27608 6502 27660 6554
rect 27672 6502 27724 6554
rect 27736 6502 27788 6554
rect 27800 6502 27852 6554
rect 27864 6502 27916 6554
rect 4664 5958 4716 6010
rect 4728 5958 4780 6010
rect 4792 5958 4844 6010
rect 4856 5958 4908 6010
rect 4920 5958 4972 6010
rect 12092 5958 12144 6010
rect 12156 5958 12208 6010
rect 12220 5958 12272 6010
rect 12284 5958 12336 6010
rect 12348 5958 12400 6010
rect 19520 5958 19572 6010
rect 19584 5958 19636 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 26948 5958 27000 6010
rect 27012 5958 27064 6010
rect 27076 5958 27128 6010
rect 27140 5958 27192 6010
rect 27204 5958 27256 6010
rect 5324 5414 5376 5466
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 12752 5414 12804 5466
rect 12816 5414 12868 5466
rect 12880 5414 12932 5466
rect 12944 5414 12996 5466
rect 13008 5414 13060 5466
rect 20180 5414 20232 5466
rect 20244 5414 20296 5466
rect 20308 5414 20360 5466
rect 20372 5414 20424 5466
rect 20436 5414 20488 5466
rect 27608 5414 27660 5466
rect 27672 5414 27724 5466
rect 27736 5414 27788 5466
rect 27800 5414 27852 5466
rect 27864 5414 27916 5466
rect 4664 4870 4716 4922
rect 4728 4870 4780 4922
rect 4792 4870 4844 4922
rect 4856 4870 4908 4922
rect 4920 4870 4972 4922
rect 12092 4870 12144 4922
rect 12156 4870 12208 4922
rect 12220 4870 12272 4922
rect 12284 4870 12336 4922
rect 12348 4870 12400 4922
rect 19520 4870 19572 4922
rect 19584 4870 19636 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 26948 4870 27000 4922
rect 27012 4870 27064 4922
rect 27076 4870 27128 4922
rect 27140 4870 27192 4922
rect 27204 4870 27256 4922
rect 5324 4326 5376 4378
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 12752 4326 12804 4378
rect 12816 4326 12868 4378
rect 12880 4326 12932 4378
rect 12944 4326 12996 4378
rect 13008 4326 13060 4378
rect 20180 4326 20232 4378
rect 20244 4326 20296 4378
rect 20308 4326 20360 4378
rect 20372 4326 20424 4378
rect 20436 4326 20488 4378
rect 27608 4326 27660 4378
rect 27672 4326 27724 4378
rect 27736 4326 27788 4378
rect 27800 4326 27852 4378
rect 27864 4326 27916 4378
rect 4664 3782 4716 3834
rect 4728 3782 4780 3834
rect 4792 3782 4844 3834
rect 4856 3782 4908 3834
rect 4920 3782 4972 3834
rect 12092 3782 12144 3834
rect 12156 3782 12208 3834
rect 12220 3782 12272 3834
rect 12284 3782 12336 3834
rect 12348 3782 12400 3834
rect 19520 3782 19572 3834
rect 19584 3782 19636 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 26948 3782 27000 3834
rect 27012 3782 27064 3834
rect 27076 3782 27128 3834
rect 27140 3782 27192 3834
rect 27204 3782 27256 3834
rect 5324 3238 5376 3290
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 12752 3238 12804 3290
rect 12816 3238 12868 3290
rect 12880 3238 12932 3290
rect 12944 3238 12996 3290
rect 13008 3238 13060 3290
rect 20180 3238 20232 3290
rect 20244 3238 20296 3290
rect 20308 3238 20360 3290
rect 20372 3238 20424 3290
rect 20436 3238 20488 3290
rect 27608 3238 27660 3290
rect 27672 3238 27724 3290
rect 27736 3238 27788 3290
rect 27800 3238 27852 3290
rect 27864 3238 27916 3290
rect 4664 2694 4716 2746
rect 4728 2694 4780 2746
rect 4792 2694 4844 2746
rect 4856 2694 4908 2746
rect 4920 2694 4972 2746
rect 12092 2694 12144 2746
rect 12156 2694 12208 2746
rect 12220 2694 12272 2746
rect 12284 2694 12336 2746
rect 12348 2694 12400 2746
rect 19520 2694 19572 2746
rect 19584 2694 19636 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 26948 2694 27000 2746
rect 27012 2694 27064 2746
rect 27076 2694 27128 2746
rect 27140 2694 27192 2746
rect 27204 2694 27256 2746
rect 9312 2635 9364 2644
rect 9312 2601 9321 2635
rect 9321 2601 9355 2635
rect 9355 2601 9364 2635
rect 9312 2592 9364 2601
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 11060 2592 11112 2644
rect 14004 2592 14056 2644
rect 16120 2592 16172 2644
rect 17132 2592 17184 2644
rect 17868 2592 17920 2644
rect 18972 2635 19024 2644
rect 18972 2601 18981 2635
rect 18981 2601 19015 2635
rect 19015 2601 19024 2635
rect 18972 2592 19024 2601
rect 21456 2592 21508 2644
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 15016 2363 15068 2372
rect 15016 2329 15025 2363
rect 15025 2329 15059 2363
rect 15059 2329 15068 2363
rect 15016 2320 15068 2329
rect 16948 2363 17000 2372
rect 16948 2329 16957 2363
rect 16957 2329 16991 2363
rect 16991 2329 17000 2363
rect 16948 2320 17000 2329
rect 17592 2363 17644 2372
rect 17592 2329 17601 2363
rect 17601 2329 17635 2363
rect 17635 2329 17644 2363
rect 17592 2320 17644 2329
rect 10324 2252 10376 2304
rect 12256 2252 12308 2304
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 15660 2295 15712 2304
rect 15660 2261 15669 2295
rect 15669 2261 15703 2295
rect 15703 2261 15712 2295
rect 15660 2252 15712 2261
rect 16304 2295 16356 2304
rect 16304 2261 16313 2295
rect 16313 2261 16347 2295
rect 16347 2261 16356 2295
rect 16304 2252 16356 2261
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 20628 2252 20680 2304
rect 5324 2150 5376 2202
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 12752 2150 12804 2202
rect 12816 2150 12868 2202
rect 12880 2150 12932 2202
rect 12944 2150 12996 2202
rect 13008 2150 13060 2202
rect 20180 2150 20232 2202
rect 20244 2150 20296 2202
rect 20308 2150 20360 2202
rect 20372 2150 20424 2202
rect 20436 2150 20488 2202
rect 27608 2150 27660 2202
rect 27672 2150 27724 2202
rect 27736 2150 27788 2202
rect 27800 2150 27852 2202
rect 27864 2150 27916 2202
<< metal2 >>
rect 12254 31362 12310 32000
rect 12898 31362 12954 32000
rect 14186 31362 14242 32000
rect 12254 31334 12388 31362
rect 12254 31200 12310 31334
rect 5324 29404 5632 29413
rect 5324 29402 5330 29404
rect 5386 29402 5410 29404
rect 5466 29402 5490 29404
rect 5546 29402 5570 29404
rect 5626 29402 5632 29404
rect 5386 29350 5388 29402
rect 5568 29350 5570 29402
rect 5324 29348 5330 29350
rect 5386 29348 5410 29350
rect 5466 29348 5490 29350
rect 5546 29348 5570 29350
rect 5626 29348 5632 29350
rect 5324 29339 5632 29348
rect 12360 29306 12388 31334
rect 12898 31334 13124 31362
rect 12898 31200 12954 31334
rect 12752 29404 13060 29413
rect 12752 29402 12758 29404
rect 12814 29402 12838 29404
rect 12894 29402 12918 29404
rect 12974 29402 12998 29404
rect 13054 29402 13060 29404
rect 12814 29350 12816 29402
rect 12996 29350 12998 29402
rect 12752 29348 12758 29350
rect 12814 29348 12838 29350
rect 12894 29348 12918 29350
rect 12974 29348 12998 29350
rect 13054 29348 13060 29350
rect 12752 29339 13060 29348
rect 13096 29306 13124 31334
rect 14186 31334 14320 31362
rect 14186 31200 14242 31334
rect 14292 29306 14320 31334
rect 14830 31200 14886 32000
rect 15474 31362 15530 32000
rect 15474 31334 15792 31362
rect 15474 31200 15530 31334
rect 12348 29300 12400 29306
rect 12348 29242 12400 29248
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14844 29238 14872 31200
rect 15764 29306 15792 31334
rect 18694 31200 18750 32000
rect 19338 31362 19394 32000
rect 19338 31334 19656 31362
rect 19338 31200 19394 31334
rect 18708 29306 18736 31200
rect 19628 29306 19656 31334
rect 20626 31200 20682 32000
rect 21914 31200 21970 32000
rect 20180 29404 20488 29413
rect 20180 29402 20186 29404
rect 20242 29402 20266 29404
rect 20322 29402 20346 29404
rect 20402 29402 20426 29404
rect 20482 29402 20488 29404
rect 20242 29350 20244 29402
rect 20424 29350 20426 29402
rect 20180 29348 20186 29350
rect 20242 29348 20266 29350
rect 20322 29348 20346 29350
rect 20402 29348 20426 29350
rect 20482 29348 20488 29350
rect 20180 29339 20488 29348
rect 20640 29306 20668 31200
rect 21928 29306 21956 31200
rect 27608 29404 27916 29413
rect 27608 29402 27614 29404
rect 27670 29402 27694 29404
rect 27750 29402 27774 29404
rect 27830 29402 27854 29404
rect 27910 29402 27916 29404
rect 27670 29350 27672 29402
rect 27852 29350 27854 29402
rect 27608 29348 27614 29350
rect 27670 29348 27694 29350
rect 27750 29348 27774 29350
rect 27830 29348 27854 29350
rect 27910 29348 27916 29350
rect 27608 29339 27916 29348
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 18696 29300 18748 29306
rect 18696 29242 18748 29248
rect 19616 29300 19668 29306
rect 19616 29242 19668 29248
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 14832 29232 14884 29238
rect 14832 29174 14884 29180
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 12532 29028 12584 29034
rect 12532 28970 12584 28976
rect 4664 28860 4972 28869
rect 4664 28858 4670 28860
rect 4726 28858 4750 28860
rect 4806 28858 4830 28860
rect 4886 28858 4910 28860
rect 4966 28858 4972 28860
rect 4726 28806 4728 28858
rect 4908 28806 4910 28858
rect 4664 28804 4670 28806
rect 4726 28804 4750 28806
rect 4806 28804 4830 28806
rect 4886 28804 4910 28806
rect 4966 28804 4972 28806
rect 4664 28795 4972 28804
rect 12092 28860 12400 28869
rect 12092 28858 12098 28860
rect 12154 28858 12178 28860
rect 12234 28858 12258 28860
rect 12314 28858 12338 28860
rect 12394 28858 12400 28860
rect 12154 28806 12156 28858
rect 12336 28806 12338 28858
rect 12092 28804 12098 28806
rect 12154 28804 12178 28806
rect 12234 28804 12258 28806
rect 12314 28804 12338 28806
rect 12394 28804 12400 28806
rect 12092 28795 12400 28804
rect 5324 28316 5632 28325
rect 5324 28314 5330 28316
rect 5386 28314 5410 28316
rect 5466 28314 5490 28316
rect 5546 28314 5570 28316
rect 5626 28314 5632 28316
rect 5386 28262 5388 28314
rect 5568 28262 5570 28314
rect 5324 28260 5330 28262
rect 5386 28260 5410 28262
rect 5466 28260 5490 28262
rect 5546 28260 5570 28262
rect 5626 28260 5632 28262
rect 5324 28251 5632 28260
rect 4664 27772 4972 27781
rect 4664 27770 4670 27772
rect 4726 27770 4750 27772
rect 4806 27770 4830 27772
rect 4886 27770 4910 27772
rect 4966 27770 4972 27772
rect 4726 27718 4728 27770
rect 4908 27718 4910 27770
rect 4664 27716 4670 27718
rect 4726 27716 4750 27718
rect 4806 27716 4830 27718
rect 4886 27716 4910 27718
rect 4966 27716 4972 27718
rect 4664 27707 4972 27716
rect 12092 27772 12400 27781
rect 12092 27770 12098 27772
rect 12154 27770 12178 27772
rect 12234 27770 12258 27772
rect 12314 27770 12338 27772
rect 12394 27770 12400 27772
rect 12154 27718 12156 27770
rect 12336 27718 12338 27770
rect 12092 27716 12098 27718
rect 12154 27716 12178 27718
rect 12234 27716 12258 27718
rect 12314 27716 12338 27718
rect 12394 27716 12400 27718
rect 12092 27707 12400 27716
rect 5324 27228 5632 27237
rect 5324 27226 5330 27228
rect 5386 27226 5410 27228
rect 5466 27226 5490 27228
rect 5546 27226 5570 27228
rect 5626 27226 5632 27228
rect 5386 27174 5388 27226
rect 5568 27174 5570 27226
rect 5324 27172 5330 27174
rect 5386 27172 5410 27174
rect 5466 27172 5490 27174
rect 5546 27172 5570 27174
rect 5626 27172 5632 27174
rect 5324 27163 5632 27172
rect 4664 26684 4972 26693
rect 4664 26682 4670 26684
rect 4726 26682 4750 26684
rect 4806 26682 4830 26684
rect 4886 26682 4910 26684
rect 4966 26682 4972 26684
rect 4726 26630 4728 26682
rect 4908 26630 4910 26682
rect 4664 26628 4670 26630
rect 4726 26628 4750 26630
rect 4806 26628 4830 26630
rect 4886 26628 4910 26630
rect 4966 26628 4972 26630
rect 4664 26619 4972 26628
rect 12092 26684 12400 26693
rect 12092 26682 12098 26684
rect 12154 26682 12178 26684
rect 12234 26682 12258 26684
rect 12314 26682 12338 26684
rect 12394 26682 12400 26684
rect 12154 26630 12156 26682
rect 12336 26630 12338 26682
rect 12092 26628 12098 26630
rect 12154 26628 12178 26630
rect 12234 26628 12258 26630
rect 12314 26628 12338 26630
rect 12394 26628 12400 26630
rect 12092 26619 12400 26628
rect 5324 26140 5632 26149
rect 5324 26138 5330 26140
rect 5386 26138 5410 26140
rect 5466 26138 5490 26140
rect 5546 26138 5570 26140
rect 5626 26138 5632 26140
rect 5386 26086 5388 26138
rect 5568 26086 5570 26138
rect 5324 26084 5330 26086
rect 5386 26084 5410 26086
rect 5466 26084 5490 26086
rect 5546 26084 5570 26086
rect 5626 26084 5632 26086
rect 5324 26075 5632 26084
rect 4664 25596 4972 25605
rect 4664 25594 4670 25596
rect 4726 25594 4750 25596
rect 4806 25594 4830 25596
rect 4886 25594 4910 25596
rect 4966 25594 4972 25596
rect 4726 25542 4728 25594
rect 4908 25542 4910 25594
rect 4664 25540 4670 25542
rect 4726 25540 4750 25542
rect 4806 25540 4830 25542
rect 4886 25540 4910 25542
rect 4966 25540 4972 25542
rect 4664 25531 4972 25540
rect 12092 25596 12400 25605
rect 12092 25594 12098 25596
rect 12154 25594 12178 25596
rect 12234 25594 12258 25596
rect 12314 25594 12338 25596
rect 12394 25594 12400 25596
rect 12154 25542 12156 25594
rect 12336 25542 12338 25594
rect 12092 25540 12098 25542
rect 12154 25540 12178 25542
rect 12234 25540 12258 25542
rect 12314 25540 12338 25542
rect 12394 25540 12400 25542
rect 12092 25531 12400 25540
rect 3422 25256 3478 25265
rect 3422 25191 3478 25200
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1504 23497 1532 23666
rect 1490 23488 1546 23497
rect 1490 23423 1546 23432
rect 938 22536 994 22545
rect 938 22471 940 22480
rect 992 22471 994 22480
rect 940 22442 992 22448
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 940 21888 992 21894
rect 938 21856 940 21865
rect 992 21856 994 21865
rect 938 21791 994 21800
rect 1688 21350 1716 21966
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 952 21185 980 21286
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20641 1532 20742
rect 1490 20632 1546 20641
rect 1490 20567 1546 20576
rect 938 19816 994 19825
rect 938 19751 940 19760
rect 992 19751 994 19760
rect 940 19722 992 19728
rect 3344 19378 3372 20878
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 1412 19281 1440 19314
rect 1398 19272 1454 19281
rect 1398 19207 1454 19216
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 18465 980 18702
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17921 1532 18226
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 940 17128 992 17134
rect 938 17096 940 17105
rect 1676 17128 1728 17134
rect 992 17096 994 17105
rect 1676 17070 1728 17076
rect 938 17031 994 17040
rect 1688 16794 1716 17070
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 3436 16522 3464 25191
rect 5324 25052 5632 25061
rect 5324 25050 5330 25052
rect 5386 25050 5410 25052
rect 5466 25050 5490 25052
rect 5546 25050 5570 25052
rect 5626 25050 5632 25052
rect 5386 24998 5388 25050
rect 5568 24998 5570 25050
rect 5324 24996 5330 24998
rect 5386 24996 5410 24998
rect 5466 24996 5490 24998
rect 5546 24996 5570 24998
rect 5626 24996 5632 24998
rect 5324 24987 5632 24996
rect 4664 24508 4972 24517
rect 4664 24506 4670 24508
rect 4726 24506 4750 24508
rect 4806 24506 4830 24508
rect 4886 24506 4910 24508
rect 4966 24506 4972 24508
rect 4726 24454 4728 24506
rect 4908 24454 4910 24506
rect 4664 24452 4670 24454
rect 4726 24452 4750 24454
rect 4806 24452 4830 24454
rect 4886 24452 4910 24454
rect 4966 24452 4972 24454
rect 4664 24443 4972 24452
rect 12092 24508 12400 24517
rect 12092 24506 12098 24508
rect 12154 24506 12178 24508
rect 12234 24506 12258 24508
rect 12314 24506 12338 24508
rect 12394 24506 12400 24508
rect 12154 24454 12156 24506
rect 12336 24454 12338 24506
rect 12092 24452 12098 24454
rect 12154 24452 12178 24454
rect 12234 24452 12258 24454
rect 12314 24452 12338 24454
rect 12394 24452 12400 24454
rect 12092 24443 12400 24452
rect 5324 23964 5632 23973
rect 5324 23962 5330 23964
rect 5386 23962 5410 23964
rect 5466 23962 5490 23964
rect 5546 23962 5570 23964
rect 5626 23962 5632 23964
rect 5386 23910 5388 23962
rect 5568 23910 5570 23962
rect 5324 23908 5330 23910
rect 5386 23908 5410 23910
rect 5466 23908 5490 23910
rect 5546 23908 5570 23910
rect 5626 23908 5632 23910
rect 5324 23899 5632 23908
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 6920 23588 6972 23594
rect 6920 23530 6972 23536
rect 4664 23420 4972 23429
rect 4664 23418 4670 23420
rect 4726 23418 4750 23420
rect 4806 23418 4830 23420
rect 4886 23418 4910 23420
rect 4966 23418 4972 23420
rect 4726 23366 4728 23418
rect 4908 23366 4910 23418
rect 4664 23364 4670 23366
rect 4726 23364 4750 23366
rect 4806 23364 4830 23366
rect 4886 23364 4910 23366
rect 4966 23364 4972 23366
rect 4664 23355 4972 23364
rect 5324 22876 5632 22885
rect 5324 22874 5330 22876
rect 5386 22874 5410 22876
rect 5466 22874 5490 22876
rect 5546 22874 5570 22876
rect 5626 22874 5632 22876
rect 5386 22822 5388 22874
rect 5568 22822 5570 22874
rect 5324 22820 5330 22822
rect 5386 22820 5410 22822
rect 5466 22820 5490 22822
rect 5546 22820 5570 22822
rect 5626 22820 5632 22822
rect 5324 22811 5632 22820
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 6092 22636 6144 22642
rect 6092 22578 6144 22584
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 20942 3832 21966
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 4448 19514 4476 22578
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4664 22332 4972 22341
rect 4664 22330 4670 22332
rect 4726 22330 4750 22332
rect 4806 22330 4830 22332
rect 4886 22330 4910 22332
rect 4966 22330 4972 22332
rect 4726 22278 4728 22330
rect 4908 22278 4910 22330
rect 4664 22276 4670 22278
rect 4726 22276 4750 22278
rect 4806 22276 4830 22278
rect 4886 22276 4910 22278
rect 4966 22276 4972 22278
rect 4664 22267 4972 22276
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4632 21690 4660 21898
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 5092 21554 5120 22374
rect 5184 22234 5212 22510
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5368 21962 5396 22374
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4664 21244 4972 21253
rect 4664 21242 4670 21244
rect 4726 21242 4750 21244
rect 4806 21242 4830 21244
rect 4886 21242 4910 21244
rect 4966 21242 4972 21244
rect 4726 21190 4728 21242
rect 4908 21190 4910 21242
rect 4664 21188 4670 21190
rect 4726 21188 4750 21190
rect 4806 21188 4830 21190
rect 4886 21188 4910 21190
rect 4966 21188 4972 21190
rect 4664 21179 4972 21188
rect 5184 21146 5212 21830
rect 5324 21788 5632 21797
rect 5324 21786 5330 21788
rect 5386 21786 5410 21788
rect 5466 21786 5490 21788
rect 5546 21786 5570 21788
rect 5626 21786 5632 21788
rect 5386 21734 5388 21786
rect 5568 21734 5570 21786
rect 5324 21732 5330 21734
rect 5386 21732 5410 21734
rect 5466 21732 5490 21734
rect 5546 21732 5570 21734
rect 5626 21732 5632 21734
rect 5324 21723 5632 21732
rect 5736 21570 5764 22170
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5552 21554 5764 21570
rect 5540 21548 5764 21554
rect 5592 21542 5764 21548
rect 5540 21490 5592 21496
rect 5828 21486 5856 21966
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5324 20700 5632 20709
rect 5324 20698 5330 20700
rect 5386 20698 5410 20700
rect 5466 20698 5490 20700
rect 5546 20698 5570 20700
rect 5626 20698 5632 20700
rect 5386 20646 5388 20698
rect 5568 20646 5570 20698
rect 5324 20644 5330 20646
rect 5386 20644 5410 20646
rect 5466 20644 5490 20646
rect 5546 20644 5570 20646
rect 5626 20644 5632 20646
rect 5324 20635 5632 20644
rect 5828 20466 5856 21422
rect 6104 21146 6132 22578
rect 6748 22234 6776 22578
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 21690 6408 21898
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6932 21434 6960 23530
rect 11808 23322 11836 23666
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 9864 23044 9916 23050
rect 9864 22986 9916 22992
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7024 21554 7052 22374
rect 7668 22098 7696 22578
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 8312 21894 8340 22510
rect 9876 22438 9904 22986
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9416 22234 9444 22374
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 7300 21690 7328 21830
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 8496 21554 8524 21830
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 6644 21412 6696 21418
rect 6932 21406 7052 21434
rect 6644 21354 6696 21360
rect 6656 21146 6684 21354
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6932 20602 6960 21286
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 4664 20156 4972 20165
rect 4664 20154 4670 20156
rect 4726 20154 4750 20156
rect 4806 20154 4830 20156
rect 4886 20154 4910 20156
rect 4966 20154 4972 20156
rect 4726 20102 4728 20154
rect 4908 20102 4910 20154
rect 4664 20100 4670 20102
rect 4726 20100 4750 20102
rect 4806 20100 4830 20102
rect 4886 20100 4910 20102
rect 4966 20100 4972 20102
rect 4664 20091 4972 20100
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3620 18970 3648 19246
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 4356 18902 4384 19450
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4448 18766 4476 19450
rect 5184 19378 5212 19654
rect 5324 19612 5632 19621
rect 5324 19610 5330 19612
rect 5386 19610 5410 19612
rect 5466 19610 5490 19612
rect 5546 19610 5570 19612
rect 5626 19610 5632 19612
rect 5386 19558 5388 19610
rect 5568 19558 5570 19610
rect 5324 19556 5330 19558
rect 5386 19556 5410 19558
rect 5466 19556 5490 19558
rect 5546 19556 5570 19558
rect 5626 19556 5632 19558
rect 5324 19547 5632 19556
rect 4620 19372 4672 19378
rect 4540 19332 4620 19360
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 3424 16516 3476 16522
rect 3424 16458 3476 16464
rect 940 16448 992 16454
rect 938 16416 940 16425
rect 992 16416 994 16425
rect 938 16351 994 16360
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 952 15745 980 15846
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 4356 15586 4384 18566
rect 4540 16658 4568 19332
rect 4620 19314 4672 19320
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 4664 19068 4972 19077
rect 4664 19066 4670 19068
rect 4726 19066 4750 19068
rect 4806 19066 4830 19068
rect 4886 19066 4910 19068
rect 4966 19066 4972 19068
rect 4726 19014 4728 19066
rect 4908 19014 4910 19066
rect 4664 19012 4670 19014
rect 4726 19012 4750 19014
rect 4806 19012 4830 19014
rect 4886 19012 4910 19014
rect 4966 19012 4972 19014
rect 4664 19003 4972 19012
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4664 17980 4972 17989
rect 4664 17978 4670 17980
rect 4726 17978 4750 17980
rect 4806 17978 4830 17980
rect 4886 17978 4910 17980
rect 4966 17978 4972 17980
rect 4726 17926 4728 17978
rect 4908 17926 4910 17978
rect 4664 17924 4670 17926
rect 4726 17924 4750 17926
rect 4806 17924 4830 17926
rect 4886 17924 4910 17926
rect 4966 17924 4972 17926
rect 4664 17915 4972 17924
rect 5000 17882 5028 18566
rect 5092 18358 5120 18838
rect 5460 18834 5488 19110
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17338 5028 17478
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5092 17202 5120 18294
rect 5184 18154 5212 18702
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 5324 18524 5632 18533
rect 5324 18522 5330 18524
rect 5386 18522 5410 18524
rect 5466 18522 5490 18524
rect 5546 18522 5570 18524
rect 5626 18522 5632 18524
rect 5386 18470 5388 18522
rect 5568 18470 5570 18522
rect 5324 18468 5330 18470
rect 5386 18468 5410 18470
rect 5466 18468 5490 18470
rect 5546 18468 5570 18470
rect 5626 18468 5632 18470
rect 5324 18459 5632 18468
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5368 17678 5396 17818
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5184 17338 5212 17614
rect 5324 17436 5632 17445
rect 5324 17434 5330 17436
rect 5386 17434 5410 17436
rect 5466 17434 5490 17436
rect 5546 17434 5570 17436
rect 5626 17434 5632 17436
rect 5386 17382 5388 17434
rect 5568 17382 5570 17434
rect 5324 17380 5330 17382
rect 5386 17380 5410 17382
rect 5466 17380 5490 17382
rect 5546 17380 5570 17382
rect 5626 17380 5632 17382
rect 5324 17371 5632 17380
rect 5172 17332 5224 17338
rect 5736 17320 5764 17682
rect 5920 17678 5948 18294
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5736 17292 5948 17320
rect 5172 17274 5224 17280
rect 5722 17232 5778 17241
rect 5080 17196 5132 17202
rect 5920 17202 5948 17292
rect 5722 17167 5724 17176
rect 5080 17138 5132 17144
rect 5776 17167 5778 17176
rect 5908 17196 5960 17202
rect 5724 17138 5776 17144
rect 5908 17138 5960 17144
rect 4664 16892 4972 16901
rect 4664 16890 4670 16892
rect 4726 16890 4750 16892
rect 4806 16890 4830 16892
rect 4886 16890 4910 16892
rect 4966 16890 4972 16892
rect 4726 16838 4728 16890
rect 4908 16838 4910 16890
rect 4664 16836 4670 16838
rect 4726 16836 4750 16838
rect 4806 16836 4830 16838
rect 4886 16836 4910 16838
rect 4966 16836 4972 16838
rect 4664 16827 4972 16836
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16250 4476 16390
rect 5184 16250 5212 16526
rect 5324 16348 5632 16357
rect 5324 16346 5330 16348
rect 5386 16346 5410 16348
rect 5466 16346 5490 16348
rect 5546 16346 5570 16348
rect 5626 16346 5632 16348
rect 5386 16294 5388 16346
rect 5568 16294 5570 16346
rect 5324 16292 5330 16294
rect 5386 16292 5410 16294
rect 5466 16292 5490 16294
rect 5546 16292 5570 16294
rect 5626 16292 5632 16294
rect 5324 16283 5632 16292
rect 4436 16244 4488 16250
rect 4436 16186 4488 16192
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4448 15706 4476 15982
rect 4664 15804 4972 15813
rect 4664 15802 4670 15804
rect 4726 15802 4750 15804
rect 4806 15802 4830 15804
rect 4886 15802 4910 15804
rect 4966 15802 4972 15804
rect 4726 15750 4728 15802
rect 4908 15750 4910 15802
rect 4664 15748 4670 15750
rect 4726 15748 4750 15750
rect 4806 15748 4830 15750
rect 4886 15748 4910 15750
rect 4966 15748 4972 15750
rect 4664 15739 4972 15748
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 4356 15558 4476 15586
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15201 1440 15438
rect 1398 15192 1454 15201
rect 1398 15127 1454 15136
rect 3240 14408 3292 14414
rect 938 14376 994 14385
rect 3240 14350 3292 14356
rect 938 14311 994 14320
rect 952 14278 980 14311
rect 940 14272 992 14278
rect 940 14214 992 14220
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 3252 13734 3280 14350
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 1676 13728 1728 13734
rect 1398 13696 1454 13705
rect 1676 13670 1728 13676
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 1398 13631 1454 13640
rect 1688 13326 1716 13670
rect 4264 13530 4292 13942
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 940 13184 992 13190
rect 940 13126 992 13132
rect 952 13025 980 13126
rect 938 13016 994 13025
rect 4080 12986 4108 13330
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 13002 4200 13126
rect 4172 12986 4384 13002
rect 938 12951 994 12960
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4172 12980 4396 12986
rect 4172 12974 4344 12980
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 3240 11688 3292 11694
rect 938 11656 994 11665
rect 3240 11630 3292 11636
rect 938 11591 994 11600
rect 3252 11354 3280 11630
rect 3988 11558 4016 12242
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 4172 11234 4200 12974
rect 4344 12922 4396 12928
rect 4252 11824 4304 11830
rect 4252 11766 4304 11772
rect 4264 11354 4292 11766
rect 4448 11694 4476 15558
rect 4908 14890 4936 15642
rect 5092 15144 5120 15982
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5264 15496 5316 15502
rect 5368 15450 5396 15846
rect 5460 15706 5488 16186
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5316 15444 5396 15450
rect 5264 15438 5396 15444
rect 5632 15496 5684 15502
rect 5736 15450 5764 17138
rect 6012 17082 6040 17682
rect 5828 17054 6040 17082
rect 5828 15638 5856 17054
rect 6104 16250 6132 18566
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5920 15978 5948 16050
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5684 15444 5764 15450
rect 5632 15438 5764 15444
rect 5276 15422 5396 15438
rect 5644 15422 5764 15438
rect 5324 15260 5632 15269
rect 5324 15258 5330 15260
rect 5386 15258 5410 15260
rect 5466 15258 5490 15260
rect 5546 15258 5570 15260
rect 5626 15258 5632 15260
rect 5386 15206 5388 15258
rect 5568 15206 5570 15258
rect 5324 15204 5330 15206
rect 5386 15204 5410 15206
rect 5466 15204 5490 15206
rect 5546 15204 5570 15206
rect 5626 15204 5632 15206
rect 5324 15195 5632 15204
rect 5736 15162 5764 15422
rect 5000 15116 5120 15144
rect 5724 15156 5776 15162
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14090 4568 14758
rect 4664 14716 4972 14725
rect 4664 14714 4670 14716
rect 4726 14714 4750 14716
rect 4806 14714 4830 14716
rect 4886 14714 4910 14716
rect 4966 14714 4972 14716
rect 4726 14662 4728 14714
rect 4908 14662 4910 14714
rect 4664 14660 4670 14662
rect 4726 14660 4750 14662
rect 4806 14660 4830 14662
rect 4886 14660 4910 14662
rect 4966 14660 4972 14662
rect 4664 14651 4972 14660
rect 4540 14062 4660 14090
rect 4632 14006 4660 14062
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 5000 13870 5028 15116
rect 5724 15098 5776 15104
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5092 14550 5120 14962
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14618 5212 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5080 14544 5132 14550
rect 5276 14498 5304 14962
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5080 14486 5132 14492
rect 5184 14470 5304 14498
rect 5644 14482 5672 14826
rect 5632 14476 5684 14482
rect 5184 14074 5212 14470
rect 5632 14418 5684 14424
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5724 14408 5776 14414
rect 5828 14396 5856 15574
rect 5920 15416 5948 15914
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 6012 15706 6040 15846
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6000 15428 6052 15434
rect 5920 15388 6000 15416
rect 6000 15370 6052 15376
rect 6012 15026 6040 15370
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6104 14890 6132 16050
rect 6196 15162 6224 17818
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 6288 17241 6316 17546
rect 6274 17232 6330 17241
rect 6274 17167 6276 17176
rect 6328 17167 6330 17176
rect 6276 17138 6328 17144
rect 6380 17116 6408 19246
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6564 18970 6592 19178
rect 6656 18970 6684 20334
rect 7024 19514 7052 21406
rect 7656 20596 7708 20602
rect 7656 20538 7708 20544
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7116 20058 7144 20470
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7392 19854 7420 20198
rect 7668 19922 7696 20538
rect 8312 20466 8340 21490
rect 8772 20806 8800 21966
rect 8956 21350 8984 21966
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8956 21146 8984 21286
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9416 21078 9444 22170
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9784 21690 9812 21966
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9876 21554 9904 22374
rect 9968 22030 9996 22510
rect 10060 22030 10088 23122
rect 11992 23118 12020 23734
rect 12092 23420 12400 23429
rect 12092 23418 12098 23420
rect 12154 23418 12178 23420
rect 12234 23418 12258 23420
rect 12314 23418 12338 23420
rect 12394 23418 12400 23420
rect 12154 23366 12156 23418
rect 12336 23366 12338 23418
rect 12092 23364 12098 23366
rect 12154 23364 12178 23366
rect 12234 23364 12258 23366
rect 12314 23364 12338 23366
rect 12394 23364 12400 23366
rect 12092 23355 12400 23364
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 11980 23112 12032 23118
rect 11980 23054 12032 23060
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11624 22234 11652 22510
rect 11612 22228 11664 22234
rect 11612 22170 11664 22176
rect 11992 22098 12020 23054
rect 12268 22710 12296 23258
rect 12256 22704 12308 22710
rect 12256 22646 12308 22652
rect 12092 22332 12400 22341
rect 12092 22330 12098 22332
rect 12154 22330 12178 22332
rect 12234 22330 12258 22332
rect 12314 22330 12338 22332
rect 12394 22330 12400 22332
rect 12154 22278 12156 22330
rect 12336 22278 12338 22330
rect 12092 22276 12098 22278
rect 12154 22276 12178 22278
rect 12234 22276 12258 22278
rect 12314 22276 12338 22278
rect 12394 22276 12400 22278
rect 12092 22267 12400 22276
rect 11980 22094 12032 22098
rect 11532 22092 12032 22094
rect 11532 22066 11980 22092
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21554 9996 21830
rect 10060 21622 10088 21966
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10336 21690 10364 21898
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 11532 21554 11560 22066
rect 11980 22034 12032 22040
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 8496 20602 8524 20742
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6472 17882 6500 18702
rect 6564 18426 6592 18702
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6748 18358 6776 18770
rect 7208 18766 7236 19654
rect 7380 19508 7432 19514
rect 7380 19450 7432 19456
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6472 17338 6500 17614
rect 6564 17338 6592 17614
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6460 17128 6512 17134
rect 6380 17088 6460 17116
rect 6380 17082 6408 17088
rect 6288 17066 6408 17082
rect 6460 17070 6512 17076
rect 6276 17060 6408 17066
rect 6328 17054 6408 17060
rect 6276 17002 6328 17008
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6288 15706 6316 15982
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6368 15428 6420 15434
rect 6472 15416 6500 16730
rect 6420 15388 6500 15416
rect 6368 15370 6420 15376
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14618 5948 14758
rect 6104 14618 6132 14826
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6196 14498 6224 15098
rect 6368 15088 6420 15094
rect 6368 15030 6420 15036
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6012 14470 6224 14498
rect 5776 14368 5948 14396
rect 5724 14350 5776 14356
rect 5552 14260 5580 14350
rect 5552 14232 5764 14260
rect 5324 14172 5632 14181
rect 5324 14170 5330 14172
rect 5386 14170 5410 14172
rect 5466 14170 5490 14172
rect 5546 14170 5570 14172
rect 5626 14170 5632 14172
rect 5386 14118 5388 14170
rect 5568 14118 5570 14170
rect 5324 14116 5330 14118
rect 5386 14116 5410 14118
rect 5466 14116 5490 14118
rect 5546 14116 5570 14118
rect 5626 14116 5632 14118
rect 5324 14107 5632 14116
rect 5736 14074 5764 14232
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4664 13628 4972 13637
rect 4664 13626 4670 13628
rect 4726 13626 4750 13628
rect 4806 13626 4830 13628
rect 4886 13626 4910 13628
rect 4966 13626 4972 13628
rect 4726 13574 4728 13626
rect 4908 13574 4910 13626
rect 4664 13572 4670 13574
rect 4726 13572 4750 13574
rect 4806 13572 4830 13574
rect 4886 13572 4910 13574
rect 4966 13572 4972 13574
rect 4664 13563 4972 13572
rect 5000 12850 5028 13806
rect 5324 13084 5632 13093
rect 5324 13082 5330 13084
rect 5386 13082 5410 13084
rect 5466 13082 5490 13084
rect 5546 13082 5570 13084
rect 5626 13082 5632 13084
rect 5386 13030 5388 13082
rect 5568 13030 5570 13082
rect 5324 13028 5330 13030
rect 5386 13028 5410 13030
rect 5466 13028 5490 13030
rect 5546 13028 5570 13030
rect 5626 13028 5632 13030
rect 5324 13019 5632 13028
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 4664 12540 4972 12549
rect 4664 12538 4670 12540
rect 4726 12538 4750 12540
rect 4806 12538 4830 12540
rect 4886 12538 4910 12540
rect 4966 12538 4972 12540
rect 4726 12486 4728 12538
rect 4908 12486 4910 12538
rect 4664 12484 4670 12486
rect 4726 12484 4750 12486
rect 4806 12484 4830 12486
rect 4886 12484 4910 12486
rect 4966 12484 4972 12486
rect 4664 12475 4972 12484
rect 5000 11898 5028 12786
rect 5552 12434 5580 12786
rect 5552 12406 5764 12434
rect 5736 12238 5764 12406
rect 5828 12238 5856 12786
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5324 11996 5632 12005
rect 5324 11994 5330 11996
rect 5386 11994 5410 11996
rect 5466 11994 5490 11996
rect 5546 11994 5570 11996
rect 5626 11994 5632 11996
rect 5386 11942 5388 11994
rect 5568 11942 5570 11994
rect 5324 11940 5330 11942
rect 5386 11940 5410 11942
rect 5466 11940 5490 11942
rect 5546 11940 5570 11942
rect 5626 11940 5632 11942
rect 5324 11931 5632 11940
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4356 11354 4384 11562
rect 4540 11558 4568 11698
rect 5736 11558 5764 12174
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 4540 11354 4568 11494
rect 4664 11452 4972 11461
rect 4664 11450 4670 11452
rect 4726 11450 4750 11452
rect 4806 11450 4830 11452
rect 4886 11450 4910 11452
rect 4966 11450 4972 11452
rect 4726 11398 4728 11450
rect 4908 11398 4910 11450
rect 4664 11396 4670 11398
rect 4726 11396 4750 11398
rect 4806 11396 4830 11398
rect 4886 11396 4910 11398
rect 4966 11396 4972 11398
rect 4664 11387 4972 11396
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4172 11206 4292 11234
rect 4264 11150 4292 11206
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 940 10464 992 10470
rect 940 10406 992 10412
rect 952 10305 980 10406
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 4264 8974 4292 11086
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 9178 4476 11018
rect 4540 10674 4568 11290
rect 5276 11150 5304 11494
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5324 10908 5632 10917
rect 5324 10906 5330 10908
rect 5386 10906 5410 10908
rect 5466 10906 5490 10908
rect 5546 10906 5570 10908
rect 5626 10906 5632 10908
rect 5386 10854 5388 10906
rect 5568 10854 5570 10906
rect 5324 10852 5330 10854
rect 5386 10852 5410 10854
rect 5466 10852 5490 10854
rect 5546 10852 5570 10854
rect 5626 10852 5632 10854
rect 5324 10843 5632 10852
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4664 10364 4972 10373
rect 4664 10362 4670 10364
rect 4726 10362 4750 10364
rect 4806 10362 4830 10364
rect 4886 10362 4910 10364
rect 4966 10362 4972 10364
rect 4726 10310 4728 10362
rect 4908 10310 4910 10362
rect 4664 10308 4670 10310
rect 4726 10308 4750 10310
rect 4806 10308 4830 10310
rect 4886 10308 4910 10310
rect 4966 10308 4972 10310
rect 4664 10299 4972 10308
rect 5828 10130 5856 12174
rect 5920 10130 5948 14368
rect 6012 13258 6040 14470
rect 6288 14346 6316 14962
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6104 14006 6132 14282
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4540 9178 4568 9590
rect 5000 9518 5028 9998
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5184 9722 5212 9862
rect 5324 9820 5632 9829
rect 5324 9818 5330 9820
rect 5386 9818 5410 9820
rect 5466 9818 5490 9820
rect 5546 9818 5570 9820
rect 5626 9818 5632 9820
rect 5386 9766 5388 9818
rect 5568 9766 5570 9818
rect 5324 9764 5330 9766
rect 5386 9764 5410 9766
rect 5466 9764 5490 9766
rect 5546 9764 5570 9766
rect 5626 9764 5632 9766
rect 5324 9755 5632 9764
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5356 9512 5408 9518
rect 5408 9460 5672 9466
rect 5356 9454 5672 9460
rect 4664 9276 4972 9285
rect 4664 9274 4670 9276
rect 4726 9274 4750 9276
rect 4806 9274 4830 9276
rect 4886 9274 4910 9276
rect 4966 9274 4972 9276
rect 4726 9222 4728 9274
rect 4908 9222 4910 9274
rect 4664 9220 4670 9222
rect 4726 9220 4750 9222
rect 4806 9220 4830 9222
rect 4886 9220 4910 9222
rect 4966 9220 4972 9222
rect 4664 9211 4972 9220
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 5000 8974 5028 9454
rect 5368 9450 5672 9454
rect 5368 9444 5684 9450
rect 5368 9438 5632 9444
rect 5632 9386 5684 9392
rect 5920 9178 5948 9930
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 4252 8968 4304 8974
rect 992 8936 994 8945
rect 4252 8910 4304 8916
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 938 8871 994 8880
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 4664 8188 4972 8197
rect 4664 8186 4670 8188
rect 4726 8186 4750 8188
rect 4806 8186 4830 8188
rect 4886 8186 4910 8188
rect 4966 8186 4972 8188
rect 4726 8134 4728 8186
rect 4908 8134 4910 8186
rect 4664 8132 4670 8134
rect 4726 8132 4750 8134
rect 4806 8132 4830 8134
rect 4886 8132 4910 8134
rect 4966 8132 4972 8134
rect 4664 8123 4972 8132
rect 940 7744 992 7750
rect 940 7686 992 7692
rect 952 7585 980 7686
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 5184 7410 5212 8842
rect 5324 8732 5632 8741
rect 5324 8730 5330 8732
rect 5386 8730 5410 8732
rect 5466 8730 5490 8732
rect 5546 8730 5570 8732
rect 5626 8730 5632 8732
rect 5386 8678 5388 8730
rect 5568 8678 5570 8730
rect 5324 8676 5330 8678
rect 5386 8676 5410 8678
rect 5466 8676 5490 8678
rect 5546 8676 5570 8678
rect 5626 8676 5632 8678
rect 5324 8667 5632 8676
rect 5920 8634 5948 8842
rect 6012 8809 6040 13194
rect 6104 12986 6132 13262
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12646 6132 12922
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6104 11150 6132 11494
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6196 10538 6224 14010
rect 6288 13938 6316 14282
rect 6380 14074 6408 15030
rect 6472 14482 6500 15388
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6472 14006 6500 14418
rect 6564 14278 6592 14554
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6288 13530 6316 13874
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6288 12850 6316 13466
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12986 6408 13126
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 12434 6316 12582
rect 6368 12436 6420 12442
rect 6288 12406 6368 12434
rect 6368 12378 6420 12384
rect 6472 12238 6500 12786
rect 6656 12442 6684 17750
rect 6748 17678 6776 17750
rect 6932 17678 6960 18702
rect 7024 18222 7052 18702
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7392 18154 7420 19450
rect 7852 19446 7880 19722
rect 7944 19514 7972 19858
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8128 19514 8156 19790
rect 8312 19514 8340 20402
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8588 20058 8616 20334
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 9324 19854 9352 20538
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9784 20262 9812 20878
rect 10232 20868 10284 20874
rect 10232 20810 10284 20816
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 10060 20058 10088 20334
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7668 18358 7696 19314
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 8024 18352 8076 18358
rect 8668 18352 8720 18358
rect 8024 18294 8076 18300
rect 8588 18312 8668 18340
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7484 18086 7512 18226
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6748 16794 6776 17614
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6840 17134 6868 17478
rect 7024 17270 7052 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7208 17134 7236 17274
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16794 7236 17070
rect 7300 16998 7328 18022
rect 7760 17678 7788 18158
rect 8036 18086 8064 18294
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7024 15502 7052 15914
rect 7208 15910 7236 16730
rect 7484 16590 7512 17138
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7484 16250 7512 16526
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7472 15972 7524 15978
rect 7472 15914 7524 15920
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15502 7236 15846
rect 7484 15502 7512 15914
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7116 14958 7144 15438
rect 7484 15026 7512 15438
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7484 14550 7512 14962
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6748 12986 6776 13330
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 7024 12850 7052 13262
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6656 11778 6684 12378
rect 7024 12306 7052 12786
rect 7852 12730 7880 13262
rect 7944 12866 7972 15642
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8036 15094 8064 15438
rect 8128 15366 8156 17138
rect 8312 16658 8340 17478
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8024 15088 8076 15094
rect 8024 15030 8076 15036
rect 8128 14958 8156 15302
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8128 14278 8156 14894
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 13734 8156 14214
rect 8220 14074 8248 14758
rect 8312 14618 8340 14962
rect 8496 14906 8524 18226
rect 8588 17116 8616 18312
rect 8668 18294 8720 18300
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 17338 8708 17614
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8772 17202 8800 19654
rect 9416 18426 9444 19654
rect 9508 19174 9536 19858
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18698 9720 19110
rect 9876 18698 9904 19790
rect 10060 18902 10088 19994
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 10048 18896 10100 18902
rect 10048 18838 10100 18844
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9496 18216 9548 18222
rect 9864 18216 9916 18222
rect 9496 18158 9548 18164
rect 9784 18164 9864 18170
rect 9784 18158 9916 18164
rect 9508 17882 9536 18158
rect 9784 18142 9904 18158
rect 9784 17882 9812 18142
rect 9496 17876 9548 17882
rect 9496 17818 9548 17824
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8668 17128 8720 17134
rect 8588 17088 8668 17116
rect 8668 17070 8720 17076
rect 8404 14878 8524 14906
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 7944 12838 8064 12866
rect 7932 12776 7984 12782
rect 7852 12724 7932 12730
rect 7852 12718 7984 12724
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7852 12702 7972 12718
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 12434 7512 12582
rect 7392 12406 7512 12434
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6656 11750 6776 11778
rect 6840 11762 6868 12038
rect 6748 11694 6776 11750
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11354 6316 11494
rect 7300 11354 7328 11562
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6380 10810 6408 11086
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6748 10742 6776 10950
rect 6932 10810 6960 11018
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 10130 6224 10474
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6748 10062 6776 10678
rect 6932 10266 6960 10746
rect 7116 10606 7144 11086
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6104 9042 6132 9454
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 9178 6316 9318
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6380 9110 6408 9454
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6092 8832 6144 8838
rect 5998 8800 6054 8809
rect 6092 8774 6144 8780
rect 5998 8735 6054 8744
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6012 8430 6040 8735
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6104 8294 6132 8774
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6380 8090 6408 8366
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6472 7886 6500 9454
rect 6656 9042 6684 9998
rect 6748 9722 6776 9998
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6840 9518 6868 9998
rect 6932 9586 6960 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 7392 9178 7420 12406
rect 7760 12306 7788 12650
rect 7852 12374 7880 12702
rect 8036 12434 8064 12838
rect 8128 12646 8156 13330
rect 8404 13002 8432 14878
rect 8588 14550 8616 14894
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8680 14006 8708 17070
rect 8772 16998 8800 17138
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8956 16794 8984 17070
rect 9048 16794 9076 17478
rect 9140 16794 9168 17682
rect 9784 17678 9812 17818
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9508 17354 9536 17546
rect 9508 17326 9720 17354
rect 9692 17270 9720 17326
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9140 14482 9168 16594
rect 9232 16250 9260 17206
rect 9312 17128 9364 17134
rect 9364 17076 9444 17082
rect 9312 17070 9444 17076
rect 9324 17054 9444 17070
rect 9416 16674 9444 17054
rect 9508 16794 9536 17206
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9692 16674 9720 17070
rect 9416 16646 9720 16674
rect 9784 16658 9812 17614
rect 9968 17270 9996 18838
rect 10152 18766 10180 20198
rect 10244 20058 10272 20810
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10336 20330 10364 20538
rect 11348 20466 11376 20946
rect 11336 20460 11388 20466
rect 11388 20420 11468 20448
rect 11336 20402 11388 20408
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10980 19378 11008 19994
rect 11256 19786 11284 20198
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10152 18272 10180 18702
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 18290 10456 18566
rect 10416 18284 10468 18290
rect 10152 18244 10272 18272
rect 10244 18154 10272 18244
rect 10416 18226 10468 18232
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 9956 17264 10008 17270
rect 9956 17206 10008 17212
rect 10152 17134 10180 18090
rect 10244 17610 10272 18090
rect 10428 17678 10456 18226
rect 10520 18222 10548 18634
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10520 17746 10548 18158
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 15706 9352 15846
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14618 9260 14894
rect 9324 14822 9352 15506
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8956 13530 8984 14350
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9232 13954 9260 14214
rect 9324 14074 9352 14758
rect 9692 14618 9720 16646
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 15706 10364 16594
rect 10416 16584 10468 16590
rect 10508 16584 10560 16590
rect 10416 16526 10468 16532
rect 10506 16552 10508 16561
rect 10560 16552 10562 16561
rect 10428 16114 10456 16526
rect 10506 16487 10562 16496
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10520 16250 10548 16390
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10612 15094 10640 19314
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18834 10824 19110
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17882 10732 18158
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10796 17218 10824 18770
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10888 17882 10916 18634
rect 10980 18290 11008 18702
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 10704 17190 10824 17218
rect 10704 15978 10732 17190
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10796 16590 10824 17070
rect 10888 16640 10916 17682
rect 11164 17338 11192 18906
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 18290 11376 18566
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11244 17808 11296 17814
rect 11244 17750 11296 17756
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10968 17196 11020 17202
rect 11020 17156 11100 17184
rect 10968 17138 11020 17144
rect 11072 16658 11100 17156
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 10968 16652 11020 16658
rect 10888 16612 10968 16640
rect 10968 16594 11020 16600
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8220 12974 8432 13002
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8036 12406 8156 12434
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7760 11150 7788 11698
rect 8128 11694 8156 12406
rect 8220 12306 8248 12974
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8312 12442 8340 12854
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8404 12442 8432 12786
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8128 11370 8156 11630
rect 7944 11342 8156 11370
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7564 9988 7616 9994
rect 7564 9930 7616 9936
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9586 7512 9862
rect 7576 9722 7604 9930
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7852 9654 7880 10066
rect 7944 10062 7972 11342
rect 8220 11014 8248 12242
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11898 8432 12174
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8576 11824 8628 11830
rect 8576 11766 8628 11772
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8404 11354 8432 11698
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8312 10810 8340 11290
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8404 10674 8432 11154
rect 8588 10810 8616 11766
rect 8680 11762 8708 12582
rect 9048 11898 9076 13398
rect 9140 12714 9168 13942
rect 9232 13926 9352 13954
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 8036 9586 8064 9998
rect 8128 9994 8156 10542
rect 8220 10198 8248 10610
rect 8772 10554 8800 11630
rect 9140 10674 9168 12650
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 11626 9260 12582
rect 9324 12442 9352 13926
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9784 13530 9812 13806
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9416 12918 9444 13194
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12442 10088 12650
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9324 11354 9352 12242
rect 9680 12232 9732 12238
rect 9600 12192 9680 12220
rect 9600 11830 9628 12192
rect 9680 12174 9732 12180
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9876 11898 9904 12174
rect 10336 12102 10364 14962
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10520 14006 10548 14214
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10704 13530 10732 15914
rect 10796 15638 10824 15982
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10980 14618 11008 16594
rect 11072 15706 11100 16594
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11164 14822 11192 16662
rect 11256 15366 11284 17750
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11348 16454 11376 17206
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11440 16182 11468 20420
rect 11532 20058 11560 21490
rect 11888 21480 11940 21486
rect 11940 21428 12020 21434
rect 11888 21422 12020 21428
rect 11900 21406 12020 21422
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11992 19938 12020 21406
rect 12092 21244 12400 21253
rect 12092 21242 12098 21244
rect 12154 21242 12178 21244
rect 12234 21242 12258 21244
rect 12314 21242 12338 21244
rect 12394 21242 12400 21244
rect 12154 21190 12156 21242
rect 12336 21190 12338 21242
rect 12092 21188 12098 21190
rect 12154 21188 12178 21190
rect 12234 21188 12258 21190
rect 12314 21188 12338 21190
rect 12394 21188 12400 21190
rect 12092 21179 12400 21188
rect 12452 21146 12480 21558
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12544 20398 12572 28970
rect 12752 28316 13060 28325
rect 12752 28314 12758 28316
rect 12814 28314 12838 28316
rect 12894 28314 12918 28316
rect 12974 28314 12998 28316
rect 13054 28314 13060 28316
rect 12814 28262 12816 28314
rect 12996 28262 12998 28314
rect 12752 28260 12758 28262
rect 12814 28260 12838 28262
rect 12894 28260 12918 28262
rect 12974 28260 12998 28262
rect 13054 28260 13060 28262
rect 12752 28251 13060 28260
rect 12752 27228 13060 27237
rect 12752 27226 12758 27228
rect 12814 27226 12838 27228
rect 12894 27226 12918 27228
rect 12974 27226 12998 27228
rect 13054 27226 13060 27228
rect 12814 27174 12816 27226
rect 12996 27174 12998 27226
rect 12752 27172 12758 27174
rect 12814 27172 12838 27174
rect 12894 27172 12918 27174
rect 12974 27172 12998 27174
rect 13054 27172 13060 27174
rect 12752 27163 13060 27172
rect 12752 26140 13060 26149
rect 12752 26138 12758 26140
rect 12814 26138 12838 26140
rect 12894 26138 12918 26140
rect 12974 26138 12998 26140
rect 13054 26138 13060 26140
rect 12814 26086 12816 26138
rect 12996 26086 12998 26138
rect 12752 26084 12758 26086
rect 12814 26084 12838 26086
rect 12894 26084 12918 26086
rect 12974 26084 12998 26086
rect 13054 26084 13060 26086
rect 12752 26075 13060 26084
rect 12752 25052 13060 25061
rect 12752 25050 12758 25052
rect 12814 25050 12838 25052
rect 12894 25050 12918 25052
rect 12974 25050 12998 25052
rect 13054 25050 13060 25052
rect 12814 24998 12816 25050
rect 12996 24998 12998 25050
rect 12752 24996 12758 24998
rect 12814 24996 12838 24998
rect 12894 24996 12918 24998
rect 12974 24996 12998 24998
rect 13054 24996 13060 24998
rect 12752 24987 13060 24996
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12636 24410 12664 24686
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12752 23964 13060 23973
rect 12752 23962 12758 23964
rect 12814 23962 12838 23964
rect 12894 23962 12918 23964
rect 12974 23962 12998 23964
rect 13054 23962 13060 23964
rect 12814 23910 12816 23962
rect 12996 23910 12998 23962
rect 12752 23908 12758 23910
rect 12814 23908 12838 23910
rect 12894 23908 12918 23910
rect 12974 23908 12998 23910
rect 13054 23908 13060 23910
rect 12752 23899 13060 23908
rect 13096 23866 13124 24142
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 13280 23594 13308 29038
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 24410 14228 24754
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14188 24404 14240 24410
rect 14188 24346 14240 24352
rect 14384 24206 14412 24686
rect 14476 24410 14504 24686
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22778 12664 22918
rect 12752 22876 13060 22885
rect 12752 22874 12758 22876
rect 12814 22874 12838 22876
rect 12894 22874 12918 22876
rect 12974 22874 12998 22876
rect 13054 22874 13060 22876
rect 12814 22822 12816 22874
rect 12996 22822 12998 22874
rect 12752 22820 12758 22822
rect 12814 22820 12838 22822
rect 12894 22820 12918 22822
rect 12974 22820 12998 22822
rect 13054 22820 13060 22822
rect 12752 22811 13060 22820
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12820 22234 12848 22374
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12752 21788 13060 21797
rect 12752 21786 12758 21788
rect 12814 21786 12838 21788
rect 12894 21786 12918 21788
rect 12974 21786 12998 21788
rect 13054 21786 13060 21788
rect 12814 21734 12816 21786
rect 12996 21734 12998 21786
rect 12752 21732 12758 21734
rect 12814 21732 12838 21734
rect 12894 21732 12918 21734
rect 12974 21732 12998 21734
rect 13054 21732 13060 21734
rect 12752 21723 13060 21732
rect 13832 21690 13860 22510
rect 13924 21894 13952 23734
rect 14292 22030 14320 24006
rect 14384 23730 14412 24142
rect 14568 24138 14596 24550
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14660 23798 14688 29106
rect 15200 29028 15252 29034
rect 15200 28970 15252 28976
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14752 24886 14780 25298
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 14740 24880 14792 24886
rect 14740 24822 14792 24828
rect 14844 24206 14872 25162
rect 14936 24206 14964 25230
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14844 23882 14872 24142
rect 14936 24018 14964 24142
rect 14936 23990 15056 24018
rect 14844 23854 14964 23882
rect 15028 23866 15056 23990
rect 14648 23792 14700 23798
rect 14648 23734 14700 23740
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14844 23186 14872 23666
rect 14936 23526 14964 23854
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 14924 23520 14976 23526
rect 14924 23462 14976 23468
rect 14936 23322 14964 23462
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 14844 22778 14872 23122
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14936 22574 14964 23258
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 15028 22438 15056 23802
rect 15108 23044 15160 23050
rect 15108 22986 15160 22992
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 14016 21486 14044 21966
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13556 21146 13584 21422
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 12752 20700 13060 20709
rect 12752 20698 12758 20700
rect 12814 20698 12838 20700
rect 12894 20698 12918 20700
rect 12974 20698 12998 20700
rect 13054 20698 13060 20700
rect 12814 20646 12816 20698
rect 12996 20646 12998 20698
rect 12752 20644 12758 20646
rect 12814 20644 12838 20646
rect 12894 20644 12918 20646
rect 12974 20644 12998 20646
rect 13054 20644 13060 20646
rect 12752 20635 13060 20644
rect 13556 20466 13584 21082
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12092 20156 12400 20165
rect 12092 20154 12098 20156
rect 12154 20154 12178 20156
rect 12234 20154 12258 20156
rect 12314 20154 12338 20156
rect 12394 20154 12400 20156
rect 12154 20102 12156 20154
rect 12336 20102 12338 20154
rect 12092 20100 12098 20102
rect 12154 20100 12178 20102
rect 12234 20100 12258 20102
rect 12314 20100 12338 20102
rect 12394 20100 12400 20102
rect 12092 20091 12400 20100
rect 12072 19984 12124 19990
rect 11992 19932 12072 19938
rect 11992 19926 12124 19932
rect 11992 19910 12112 19926
rect 12544 19854 12572 20334
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11624 18850 11652 19314
rect 11716 18970 11744 19722
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11624 18822 11744 18850
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11624 18426 11652 18702
rect 11716 18426 11744 18822
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11624 18086 11652 18226
rect 11808 18222 11836 18906
rect 11900 18766 11928 19110
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11888 18352 11940 18358
rect 11992 18329 12020 19654
rect 12084 19514 12112 19722
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12360 19378 12388 19654
rect 12452 19378 12480 19790
rect 12636 19378 12664 20402
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12752 19612 13060 19621
rect 12752 19610 12758 19612
rect 12814 19610 12838 19612
rect 12894 19610 12918 19612
rect 12974 19610 12998 19612
rect 13054 19610 13060 19612
rect 12814 19558 12816 19610
rect 12996 19558 12998 19610
rect 12752 19556 12758 19558
rect 12814 19556 12838 19558
rect 12894 19556 12918 19558
rect 12974 19556 12998 19558
rect 13054 19556 13060 19558
rect 12752 19547 13060 19556
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12092 19068 12400 19077
rect 12092 19066 12098 19068
rect 12154 19066 12178 19068
rect 12234 19066 12258 19068
rect 12314 19066 12338 19068
rect 12394 19066 12400 19068
rect 12154 19014 12156 19066
rect 12336 19014 12338 19066
rect 12092 19012 12098 19014
rect 12154 19012 12178 19014
rect 12234 19012 12258 19014
rect 12314 19012 12338 19014
rect 12394 19012 12400 19014
rect 12092 19003 12400 19012
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 11888 18294 11940 18300
rect 11978 18320 12034 18329
rect 11900 18222 11928 18294
rect 11978 18255 12034 18264
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11992 17746 12020 18158
rect 12268 18154 12296 18362
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12452 18086 12480 19178
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12092 17980 12400 17989
rect 12092 17978 12098 17980
rect 12154 17978 12178 17980
rect 12234 17978 12258 17980
rect 12314 17978 12338 17980
rect 12394 17978 12400 17980
rect 12154 17926 12156 17978
rect 12336 17926 12338 17978
rect 12092 17924 12098 17926
rect 12154 17924 12178 17926
rect 12234 17924 12258 17926
rect 12314 17924 12338 17926
rect 12394 17924 12400 17926
rect 12092 17915 12400 17924
rect 11980 17740 12032 17746
rect 12032 17700 12112 17728
rect 11980 17682 12032 17688
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11624 16998 11652 17274
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11808 16794 11836 17138
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11992 16590 12020 17070
rect 12084 17066 12112 17700
rect 12452 17202 12480 18022
rect 12544 17354 12572 18634
rect 12636 18426 12664 18634
rect 12752 18524 13060 18533
rect 12752 18522 12758 18524
rect 12814 18522 12838 18524
rect 12894 18522 12918 18524
rect 12974 18522 12998 18524
rect 13054 18522 13060 18524
rect 12814 18470 12816 18522
rect 12996 18470 12998 18522
rect 12752 18468 12758 18470
rect 12814 18468 12838 18470
rect 12894 18468 12918 18470
rect 12974 18468 12998 18470
rect 13054 18468 13060 18470
rect 12752 18459 13060 18468
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12752 17436 13060 17445
rect 12752 17434 12758 17436
rect 12814 17434 12838 17436
rect 12894 17434 12918 17436
rect 12974 17434 12998 17436
rect 13054 17434 13060 17436
rect 12814 17382 12816 17434
rect 12996 17382 12998 17434
rect 12752 17380 12758 17382
rect 12814 17380 12838 17382
rect 12894 17380 12918 17382
rect 12974 17380 12998 17382
rect 13054 17380 13060 17382
rect 12752 17371 13060 17380
rect 12544 17326 12664 17354
rect 13096 17338 13124 19858
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13188 18970 13216 19314
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13280 18766 13308 20198
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13372 18970 13400 19314
rect 13740 19310 13768 19654
rect 14016 19378 14044 21422
rect 14292 21078 14320 21966
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21554 14412 21830
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14280 21072 14332 21078
rect 14280 21014 14332 21020
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14292 19378 14320 20334
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 14200 18834 14228 19110
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 18086 13216 18226
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17814 14228 18022
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 14292 17746 14320 19314
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14384 18426 14412 18838
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12092 16892 12400 16901
rect 12092 16890 12098 16892
rect 12154 16890 12178 16892
rect 12234 16890 12258 16892
rect 12314 16890 12338 16892
rect 12394 16890 12400 16892
rect 12154 16838 12156 16890
rect 12336 16838 12338 16890
rect 12092 16836 12098 16838
rect 12154 16836 12178 16838
rect 12234 16836 12258 16838
rect 12314 16836 12338 16838
rect 12394 16836 12400 16838
rect 12092 16827 12400 16836
rect 12452 16590 12480 16934
rect 12544 16590 12572 17206
rect 12636 16794 12664 17326
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13096 16794 13124 17274
rect 13648 17202 13676 17478
rect 13740 17338 13768 17614
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 14476 17202 14504 19858
rect 14568 19378 14596 22374
rect 15120 22250 15148 22986
rect 15028 22222 15148 22250
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21690 14872 21830
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 15028 21622 15056 22222
rect 15212 21842 15240 28970
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15396 23866 15424 24074
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15396 22166 15424 23802
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 15304 21978 15332 22102
rect 15304 21950 15424 21978
rect 15120 21814 15240 21842
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20534 14780 20742
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19378 14872 19790
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14568 18970 14596 19314
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14660 18766 14688 19178
rect 14844 18766 14872 19314
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17338 14780 17478
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 11992 16250 12020 16526
rect 13188 16522 13216 17138
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 12752 16348 13060 16357
rect 12752 16346 12758 16348
rect 12814 16346 12838 16348
rect 12894 16346 12918 16348
rect 12974 16346 12998 16348
rect 13054 16346 13060 16348
rect 12814 16294 12816 16346
rect 12996 16294 12998 16346
rect 12752 16292 12758 16294
rect 12814 16292 12838 16294
rect 12894 16292 12918 16294
rect 12974 16292 12998 16294
rect 13054 16292 13060 16294
rect 12752 16283 13060 16292
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 11428 15972 11480 15978
rect 11428 15914 11480 15920
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11440 15026 11468 15914
rect 11624 15502 11652 16118
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12092 15804 12400 15813
rect 12092 15802 12098 15804
rect 12154 15802 12178 15804
rect 12234 15802 12258 15804
rect 12314 15802 12338 15804
rect 12394 15802 12400 15804
rect 12154 15750 12156 15802
rect 12336 15750 12338 15802
rect 12092 15748 12098 15750
rect 12154 15748 12178 15750
rect 12234 15748 12258 15750
rect 12314 15748 12338 15750
rect 12394 15748 12400 15750
rect 12092 15739 12400 15748
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11532 13870 11560 15438
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12084 15162 12112 15370
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12544 14958 12572 15506
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12636 15162 12664 15370
rect 12752 15260 13060 15269
rect 12752 15258 12758 15260
rect 12814 15258 12838 15260
rect 12894 15258 12918 15260
rect 12974 15258 12998 15260
rect 13054 15258 13060 15260
rect 12814 15206 12816 15258
rect 12996 15206 12998 15258
rect 12752 15204 12758 15206
rect 12814 15204 12838 15206
rect 12894 15204 12918 15206
rect 12974 15204 12998 15206
rect 13054 15204 13060 15206
rect 12752 15195 13060 15204
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 13280 15026 13308 15982
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12092 14716 12400 14725
rect 12092 14714 12098 14716
rect 12154 14714 12178 14716
rect 12234 14714 12258 14716
rect 12314 14714 12338 14716
rect 12394 14714 12400 14716
rect 12154 14662 12156 14714
rect 12336 14662 12338 14714
rect 12092 14660 12098 14662
rect 12154 14660 12178 14662
rect 12234 14660 12258 14662
rect 12314 14660 12338 14662
rect 12394 14660 12400 14662
rect 12092 14651 12400 14660
rect 12636 14414 12664 14894
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 14006 12388 14214
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12986 10548 13262
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11440 12986 11468 13126
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10428 12374 10456 12854
rect 11152 12776 11204 12782
rect 11058 12744 11114 12753
rect 10968 12708 11020 12714
rect 11152 12718 11204 12724
rect 11058 12679 11114 12688
rect 10968 12650 11020 12656
rect 10980 12442 11008 12650
rect 11072 12646 11100 12679
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11164 12442 11192 12718
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9128 10668 9180 10674
rect 9772 10668 9824 10674
rect 9128 10610 9180 10616
rect 9508 10628 9772 10656
rect 8944 10600 8996 10606
rect 8772 10526 8892 10554
rect 8944 10542 8996 10548
rect 8864 10470 8892 10526
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8404 9994 8432 10406
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8128 9722 8156 9930
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 6828 9104 6880 9110
rect 6828 9046 6880 9052
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6564 8090 6592 8502
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6748 7886 6776 8366
rect 7392 8294 7420 9114
rect 7484 8498 7512 9114
rect 7840 8832 7892 8838
rect 7892 8792 7972 8820
rect 7840 8774 7892 8780
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7668 8498 7696 8570
rect 7944 8498 7972 8792
rect 8312 8498 8340 9522
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7116 7954 7144 8230
rect 7944 8090 7972 8434
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7840 8016 7892 8022
rect 8036 7970 8064 8434
rect 8312 8090 8340 8434
rect 8404 8362 8432 9930
rect 8680 9518 8708 9998
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8772 9178 8800 10406
rect 8956 10266 8984 10542
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9508 10062 9536 10628
rect 9772 10610 9824 10616
rect 9588 10464 9640 10470
rect 9876 10418 9904 11018
rect 9588 10406 9640 10412
rect 9600 10062 9628 10406
rect 9784 10390 9904 10418
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9784 9450 9812 10390
rect 9968 10062 9996 11494
rect 10428 10742 10456 12310
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 12102 10732 12174
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11694 10732 12038
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10140 10668 10192 10674
rect 10324 10668 10376 10674
rect 10192 10628 10324 10656
rect 10140 10610 10192 10616
rect 10324 10610 10376 10616
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8496 8430 8524 8910
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 9048 8294 9076 9046
rect 9784 8974 9812 9386
rect 10336 9382 10364 10610
rect 10428 10062 10456 10678
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10554 10640 10610
rect 10796 10554 10824 11698
rect 11164 11150 11192 12378
rect 11348 12238 11376 12582
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11348 11286 11376 12174
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11072 10674 11100 10950
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10612 10526 10824 10554
rect 10612 10266 10640 10526
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10612 9722 10640 10202
rect 11164 9722 11192 10746
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10062 11284 10610
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 9178 10364 9318
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9968 8974 9996 9046
rect 10704 8974 10732 9454
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7892 7964 8064 7970
rect 7840 7958 8064 7964
rect 7104 7948 7156 7954
rect 7852 7942 8064 7958
rect 7104 7890 7156 7896
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5324 7644 5632 7653
rect 5324 7642 5330 7644
rect 5386 7642 5410 7644
rect 5466 7642 5490 7644
rect 5546 7642 5570 7644
rect 5626 7642 5632 7644
rect 5386 7590 5388 7642
rect 5568 7590 5570 7642
rect 5324 7588 5330 7590
rect 5386 7588 5410 7590
rect 5466 7588 5490 7590
rect 5546 7588 5570 7590
rect 5626 7588 5632 7590
rect 5324 7579 5632 7588
rect 5736 7546 5764 7754
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 6380 7478 6408 7686
rect 6472 7546 6500 7822
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 1412 6905 1440 7346
rect 4664 7100 4972 7109
rect 4664 7098 4670 7100
rect 4726 7098 4750 7100
rect 4806 7098 4830 7100
rect 4886 7098 4910 7100
rect 4966 7098 4972 7100
rect 4726 7046 4728 7098
rect 4908 7046 4910 7098
rect 4664 7044 4670 7046
rect 4726 7044 4750 7046
rect 4806 7044 4830 7046
rect 4886 7044 4910 7046
rect 4966 7044 4972 7046
rect 4664 7035 4972 7044
rect 8312 7002 8340 7346
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 1398 6896 1454 6905
rect 9140 6866 9168 8774
rect 9232 8566 9260 8910
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9416 8634 9444 8842
rect 9508 8809 9536 8842
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9508 8498 9536 8570
rect 9692 8498 9720 8842
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9968 8430 9996 8910
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 9588 8424 9640 8430
rect 9232 8372 9588 8378
rect 9232 8366 9640 8372
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9232 8350 9628 8366
rect 9232 8294 9260 8350
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 1398 6831 1454 6840
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 5324 6556 5632 6565
rect 5324 6554 5330 6556
rect 5386 6554 5410 6556
rect 5466 6554 5490 6556
rect 5546 6554 5570 6556
rect 5626 6554 5632 6556
rect 5386 6502 5388 6554
rect 5568 6502 5570 6554
rect 5324 6500 5330 6502
rect 5386 6500 5410 6502
rect 5466 6500 5490 6502
rect 5546 6500 5570 6502
rect 5626 6500 5632 6502
rect 5324 6491 5632 6500
rect 4664 6012 4972 6021
rect 4664 6010 4670 6012
rect 4726 6010 4750 6012
rect 4806 6010 4830 6012
rect 4886 6010 4910 6012
rect 4966 6010 4972 6012
rect 4726 5958 4728 6010
rect 4908 5958 4910 6010
rect 4664 5956 4670 5958
rect 4726 5956 4750 5958
rect 4806 5956 4830 5958
rect 4886 5956 4910 5958
rect 4966 5956 4972 5958
rect 4664 5947 4972 5956
rect 5324 5468 5632 5477
rect 5324 5466 5330 5468
rect 5386 5466 5410 5468
rect 5466 5466 5490 5468
rect 5546 5466 5570 5468
rect 5626 5466 5632 5468
rect 5386 5414 5388 5466
rect 5568 5414 5570 5466
rect 5324 5412 5330 5414
rect 5386 5412 5410 5414
rect 5466 5412 5490 5414
rect 5546 5412 5570 5414
rect 5626 5412 5632 5414
rect 5324 5403 5632 5412
rect 4664 4924 4972 4933
rect 4664 4922 4670 4924
rect 4726 4922 4750 4924
rect 4806 4922 4830 4924
rect 4886 4922 4910 4924
rect 4966 4922 4972 4924
rect 4726 4870 4728 4922
rect 4908 4870 4910 4922
rect 4664 4868 4670 4870
rect 4726 4868 4750 4870
rect 4806 4868 4830 4870
rect 4886 4868 4910 4870
rect 4966 4868 4972 4870
rect 4664 4859 4972 4868
rect 5324 4380 5632 4389
rect 5324 4378 5330 4380
rect 5386 4378 5410 4380
rect 5466 4378 5490 4380
rect 5546 4378 5570 4380
rect 5626 4378 5632 4380
rect 5386 4326 5388 4378
rect 5568 4326 5570 4378
rect 5324 4324 5330 4326
rect 5386 4324 5410 4326
rect 5466 4324 5490 4326
rect 5546 4324 5570 4326
rect 5626 4324 5632 4326
rect 5324 4315 5632 4324
rect 4664 3836 4972 3845
rect 4664 3834 4670 3836
rect 4726 3834 4750 3836
rect 4806 3834 4830 3836
rect 4886 3834 4910 3836
rect 4966 3834 4972 3836
rect 4726 3782 4728 3834
rect 4908 3782 4910 3834
rect 4664 3780 4670 3782
rect 4726 3780 4750 3782
rect 4806 3780 4830 3782
rect 4886 3780 4910 3782
rect 4966 3780 4972 3782
rect 4664 3771 4972 3780
rect 5324 3292 5632 3301
rect 5324 3290 5330 3292
rect 5386 3290 5410 3292
rect 5466 3290 5490 3292
rect 5546 3290 5570 3292
rect 5626 3290 5632 3292
rect 5386 3238 5388 3290
rect 5568 3238 5570 3290
rect 5324 3236 5330 3238
rect 5386 3236 5410 3238
rect 5466 3236 5490 3238
rect 5546 3236 5570 3238
rect 5626 3236 5632 3238
rect 5324 3227 5632 3236
rect 4664 2748 4972 2757
rect 4664 2746 4670 2748
rect 4726 2746 4750 2748
rect 4806 2746 4830 2748
rect 4886 2746 4910 2748
rect 4966 2746 4972 2748
rect 4726 2694 4728 2746
rect 4908 2694 4910 2746
rect 4664 2692 4670 2694
rect 4726 2692 4750 2694
rect 4806 2692 4830 2694
rect 4886 2692 4910 2694
rect 4966 2692 4972 2694
rect 4664 2683 4972 2692
rect 9324 2650 9352 8230
rect 9968 2650 9996 8366
rect 10428 8362 10456 8774
rect 10704 8634 10732 8910
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10980 8566 11008 8774
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 11256 8498 11284 8774
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 7206 10456 8298
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10428 6798 10456 7142
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10428 2446 10456 6734
rect 11348 2774 11376 11222
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11440 10742 11468 11018
rect 11428 10736 11480 10742
rect 11428 10678 11480 10684
rect 11532 10266 11560 13806
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13326 11652 13670
rect 11808 13530 11836 13806
rect 12092 13628 12400 13637
rect 12092 13626 12098 13628
rect 12154 13626 12178 13628
rect 12234 13626 12258 13628
rect 12314 13626 12338 13628
rect 12394 13626 12400 13628
rect 12154 13574 12156 13626
rect 12336 13574 12338 13626
rect 12092 13572 12098 13574
rect 12154 13572 12178 13574
rect 12234 13572 12258 13574
rect 12314 13572 12338 13574
rect 12394 13572 12400 13574
rect 12092 13563 12400 13572
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11898 11652 12038
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11900 11098 11928 12174
rect 11992 12102 12020 12582
rect 12092 12540 12400 12549
rect 12092 12538 12098 12540
rect 12154 12538 12178 12540
rect 12234 12538 12258 12540
rect 12314 12538 12338 12540
rect 12394 12538 12400 12540
rect 12154 12486 12156 12538
rect 12336 12486 12338 12538
rect 12092 12484 12098 12486
rect 12154 12484 12178 12486
rect 12234 12484 12258 12486
rect 12314 12484 12338 12486
rect 12394 12484 12400 12486
rect 12092 12475 12400 12484
rect 12636 12434 12664 14350
rect 12752 14172 13060 14181
rect 12752 14170 12758 14172
rect 12814 14170 12838 14172
rect 12894 14170 12918 14172
rect 12974 14170 12998 14172
rect 13054 14170 13060 14172
rect 12814 14118 12816 14170
rect 12996 14118 12998 14170
rect 12752 14116 12758 14118
rect 12814 14116 12838 14118
rect 12894 14116 12918 14118
rect 12974 14116 12998 14118
rect 13054 14116 13060 14118
rect 12752 14107 13060 14116
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13326 13308 13670
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12752 13084 13060 13093
rect 12752 13082 12758 13084
rect 12814 13082 12838 13084
rect 12894 13082 12918 13084
rect 12974 13082 12998 13084
rect 13054 13082 13060 13084
rect 12814 13030 12816 13082
rect 12996 13030 12998 13082
rect 12752 13028 12758 13030
rect 12814 13028 12838 13030
rect 12894 13028 12918 13030
rect 12974 13028 12998 13030
rect 13054 13028 13060 13030
rect 12752 13019 13060 13028
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12452 12406 12664 12434
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11694 12020 12038
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 11234 12020 11630
rect 12092 11452 12400 11461
rect 12092 11450 12098 11452
rect 12154 11450 12178 11452
rect 12234 11450 12258 11452
rect 12314 11450 12338 11452
rect 12394 11450 12400 11452
rect 12154 11398 12156 11450
rect 12336 11398 12338 11450
rect 12092 11396 12098 11398
rect 12154 11396 12178 11398
rect 12234 11396 12258 11398
rect 12314 11396 12338 11398
rect 12394 11396 12400 11398
rect 12092 11387 12400 11396
rect 11992 11206 12112 11234
rect 11624 10674 11652 11086
rect 11900 11070 12020 11098
rect 12084 11082 12112 11206
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10470 11652 10610
rect 11716 10538 11744 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11440 9178 11468 9522
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11532 7546 11560 10202
rect 11716 10062 11744 10474
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11624 9654 11652 9998
rect 11808 9926 11836 10542
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11808 8974 11836 9862
rect 11900 9654 11928 10610
rect 11992 10538 12020 11070
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10674 12112 11018
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11992 10062 12020 10474
rect 12092 10364 12400 10373
rect 12092 10362 12098 10364
rect 12154 10362 12178 10364
rect 12234 10362 12258 10364
rect 12314 10362 12338 10364
rect 12394 10362 12400 10364
rect 12154 10310 12156 10362
rect 12336 10310 12338 10362
rect 12092 10308 12098 10310
rect 12154 10308 12178 10310
rect 12234 10308 12258 10310
rect 12314 10308 12338 10310
rect 12394 10308 12400 10310
rect 12092 10299 12400 10308
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 12092 9276 12400 9285
rect 12092 9274 12098 9276
rect 12154 9274 12178 9276
rect 12234 9274 12258 9276
rect 12314 9274 12338 9276
rect 12394 9274 12400 9276
rect 12154 9222 12156 9274
rect 12336 9222 12338 9274
rect 12092 9220 12098 9222
rect 12154 9220 12178 9222
rect 12234 9220 12258 9222
rect 12314 9220 12338 9222
rect 12394 9220 12400 9222
rect 12092 9211 12400 9220
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 12092 8188 12400 8197
rect 12092 8186 12098 8188
rect 12154 8186 12178 8188
rect 12234 8186 12258 8188
rect 12314 8186 12338 8188
rect 12394 8186 12400 8188
rect 12154 8134 12156 8186
rect 12336 8134 12338 8186
rect 12092 8132 12098 8134
rect 12154 8132 12178 8134
rect 12234 8132 12258 8134
rect 12314 8132 12338 8134
rect 12394 8132 12400 8134
rect 12092 8123 12400 8132
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11532 7410 11560 7482
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11808 7002 11836 7278
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11992 6798 12020 7686
rect 12452 7546 12480 12406
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 10674 12664 12174
rect 12912 12170 12940 12582
rect 13096 12442 13124 13126
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 13004 12084 13032 12174
rect 13004 12056 13124 12084
rect 12752 11996 13060 12005
rect 12752 11994 12758 11996
rect 12814 11994 12838 11996
rect 12894 11994 12918 11996
rect 12974 11994 12998 11996
rect 13054 11994 13060 11996
rect 12814 11942 12816 11994
rect 12996 11942 12998 11994
rect 12752 11940 12758 11942
rect 12814 11940 12838 11942
rect 12894 11940 12918 11942
rect 12974 11940 12998 11942
rect 13054 11940 13060 11942
rect 12752 11931 13060 11940
rect 13096 11898 13124 12056
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13280 11014 13308 13262
rect 13372 12986 13400 16390
rect 13648 16114 13676 17138
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14278 16552 14334 16561
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13820 16516 13872 16522
rect 14278 16487 14280 16496
rect 13820 16458 13872 16464
rect 14332 16487 14334 16496
rect 14280 16458 14332 16464
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13556 15026 13584 15302
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13648 14906 13676 15846
rect 13740 15638 13768 16458
rect 13832 15978 13860 16458
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15434 13768 15574
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13556 14890 13676 14906
rect 14568 14890 14596 17070
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 14844 16114 14872 16458
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14936 15978 14964 19178
rect 15028 16522 15056 21558
rect 15120 19922 15148 21814
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15212 21434 15240 21626
rect 15304 21554 15332 21830
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15396 21486 15424 21950
rect 15384 21480 15436 21486
rect 15212 21406 15332 21434
rect 15384 21422 15436 21428
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15212 20058 15240 20878
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14660 15026 14688 15506
rect 15120 15502 15148 19858
rect 15304 19378 15332 21406
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15396 19310 15424 21422
rect 15488 20942 15516 22918
rect 15580 22438 15608 22918
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15580 21350 15608 21830
rect 15672 21690 15700 29106
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24886 15792 25094
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15948 24750 15976 25230
rect 16212 25220 16264 25226
rect 16212 25162 16264 25168
rect 17224 25220 17276 25226
rect 17224 25162 17276 25168
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 16028 25152 16080 25158
rect 16028 25094 16080 25100
rect 16040 24818 16068 25094
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15936 24744 15988 24750
rect 15936 24686 15988 24692
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 16132 24138 16160 24686
rect 16224 24410 16252 25162
rect 17236 24954 17264 25162
rect 17224 24948 17276 24954
rect 17224 24890 17276 24896
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16120 24132 16172 24138
rect 16120 24074 16172 24080
rect 16132 23594 16160 24074
rect 16120 23588 16172 23594
rect 16120 23530 16172 23536
rect 16132 23254 16160 23530
rect 16224 23322 16252 24346
rect 17236 24274 17540 24290
rect 17880 24274 17908 25162
rect 18144 25152 18196 25158
rect 18144 25094 18196 25100
rect 18156 24818 18184 25094
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17972 24410 18000 24550
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17236 24268 17552 24274
rect 17236 24262 17500 24268
rect 17236 24206 17264 24262
rect 17500 24210 17552 24216
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23526 16988 24006
rect 17236 23866 17264 24142
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17512 23866 17540 24006
rect 18156 23866 18184 24074
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 16212 23316 16264 23322
rect 16212 23258 16264 23264
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16120 23248 16172 23254
rect 16120 23190 16172 23196
rect 16316 22982 16344 23258
rect 17040 23112 17092 23118
rect 17144 23066 17172 23462
rect 17236 23254 17264 23802
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17972 23322 18000 23666
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17092 23060 17172 23066
rect 17040 23054 17172 23060
rect 17052 23038 17172 23054
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 21962 16160 22374
rect 16500 22234 16528 22918
rect 17052 22438 17080 23038
rect 18340 22778 18368 24754
rect 18432 24750 18460 25298
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18420 24744 18472 24750
rect 18420 24686 18472 24692
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18708 24410 18736 24686
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18524 23730 18552 24142
rect 18616 23866 18644 24278
rect 18800 24138 18828 25094
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18892 23866 18920 24142
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18616 22574 18644 23462
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 17592 22432 17644 22438
rect 17592 22374 17644 22380
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16224 22094 16436 22114
rect 16224 22086 16712 22094
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15660 21684 15712 21690
rect 15660 21626 15712 21632
rect 15764 21486 15792 21830
rect 16132 21622 16160 21898
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 16224 21486 16252 22086
rect 16408 22066 16712 22086
rect 16304 22024 16356 22030
rect 16580 22024 16632 22030
rect 16304 21966 16356 21972
rect 16500 21984 16580 22012
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16316 21418 16344 21966
rect 16500 21486 16528 21984
rect 16580 21966 16632 21972
rect 16684 21962 16712 22066
rect 16672 21956 16724 21962
rect 16672 21898 16724 21904
rect 16868 21894 16896 22170
rect 17052 22098 17080 22374
rect 17604 22234 17632 22374
rect 17592 22228 17644 22234
rect 17592 22170 17644 22176
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 17328 21622 17356 22102
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18236 22024 18288 22030
rect 18064 21984 18236 22012
rect 18064 21894 18092 21984
rect 18236 21966 18288 21972
rect 18432 21962 18460 22034
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 16304 21412 16356 21418
rect 16304 21354 16356 21360
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 19990 15516 20742
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15580 19854 15608 21286
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 18222 15240 19110
rect 15476 18624 15528 18630
rect 15476 18566 15528 18572
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15304 17338 15332 17546
rect 15488 17338 15516 18566
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15580 16794 15608 19450
rect 15672 19378 15700 21354
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15764 19854 15792 21014
rect 16500 20534 16528 21422
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15856 20058 15884 20402
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18834 15700 19314
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15764 17270 15792 19790
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15856 17542 15884 19178
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15304 16046 15332 16526
rect 15856 16114 15884 17206
rect 16040 17202 16068 19722
rect 16500 19446 16528 20470
rect 17052 19786 17080 20742
rect 17236 20602 17264 20810
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17972 19990 18000 20334
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 17052 19446 17080 19722
rect 17512 19446 17540 19858
rect 16488 19440 16540 19446
rect 16488 19382 16540 19388
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16408 18766 16436 19110
rect 16960 18970 16988 19246
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16224 17338 16252 17614
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 13544 14884 13676 14890
rect 13596 14878 13676 14884
rect 14556 14884 14608 14890
rect 13544 14826 13596 14832
rect 14556 14826 14608 14832
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13372 12646 13400 12922
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 12752 10908 13060 10917
rect 12752 10906 12758 10908
rect 12814 10906 12838 10908
rect 12894 10906 12918 10908
rect 12974 10906 12998 10908
rect 13054 10906 13060 10908
rect 12814 10854 12816 10906
rect 12996 10854 12998 10906
rect 12752 10852 12758 10854
rect 12814 10852 12838 10854
rect 12894 10852 12918 10854
rect 12974 10852 12998 10854
rect 13054 10852 13060 10854
rect 12752 10843 13060 10852
rect 13280 10674 13308 10950
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12636 10198 12664 10610
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 8838 12664 9862
rect 12752 9820 13060 9829
rect 12752 9818 12758 9820
rect 12814 9818 12838 9820
rect 12894 9818 12918 9820
rect 12974 9818 12998 9820
rect 13054 9818 13060 9820
rect 12814 9766 12816 9818
rect 12996 9766 12998 9818
rect 12752 9764 12758 9766
rect 12814 9764 12838 9766
rect 12894 9764 12918 9766
rect 12974 9764 12998 9766
rect 13054 9764 13060 9766
rect 12752 9755 13060 9764
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12912 8974 12940 9590
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12544 7954 12572 8774
rect 12752 8732 13060 8741
rect 12752 8730 12758 8732
rect 12814 8730 12838 8732
rect 12894 8730 12918 8732
rect 12974 8730 12998 8732
rect 13054 8730 13060 8732
rect 12814 8678 12816 8730
rect 12996 8678 12998 8730
rect 12752 8676 12758 8678
rect 12814 8676 12838 8678
rect 12894 8676 12918 8678
rect 12974 8676 12998 8678
rect 13054 8676 13060 8678
rect 12752 8667 13060 8676
rect 13096 8634 13124 9522
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 8634 13216 9454
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12636 7750 12664 8366
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12752 7644 13060 7653
rect 12752 7642 12758 7644
rect 12814 7642 12838 7644
rect 12894 7642 12918 7644
rect 12974 7642 12998 7644
rect 13054 7642 13060 7644
rect 12814 7590 12816 7642
rect 12996 7590 12998 7642
rect 12752 7588 12758 7590
rect 12814 7588 12838 7590
rect 12894 7588 12918 7590
rect 12974 7588 12998 7590
rect 13054 7588 13060 7590
rect 12752 7579 13060 7588
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12452 7342 12480 7482
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12092 7100 12400 7109
rect 12092 7098 12098 7100
rect 12154 7098 12178 7100
rect 12234 7098 12258 7100
rect 12314 7098 12338 7100
rect 12394 7098 12400 7100
rect 12154 7046 12156 7098
rect 12336 7046 12338 7098
rect 12092 7044 12098 7046
rect 12154 7044 12178 7046
rect 12234 7044 12258 7046
rect 12314 7044 12338 7046
rect 12394 7044 12400 7046
rect 12092 7035 12400 7044
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12092 6012 12400 6021
rect 12092 6010 12098 6012
rect 12154 6010 12178 6012
rect 12234 6010 12258 6012
rect 12314 6010 12338 6012
rect 12394 6010 12400 6012
rect 12154 5958 12156 6010
rect 12336 5958 12338 6010
rect 12092 5956 12098 5958
rect 12154 5956 12178 5958
rect 12234 5956 12258 5958
rect 12314 5956 12338 5958
rect 12394 5956 12400 5958
rect 12092 5947 12400 5956
rect 12092 4924 12400 4933
rect 12092 4922 12098 4924
rect 12154 4922 12178 4924
rect 12234 4922 12258 4924
rect 12314 4922 12338 4924
rect 12394 4922 12400 4924
rect 12154 4870 12156 4922
rect 12336 4870 12338 4922
rect 12092 4868 12098 4870
rect 12154 4868 12178 4870
rect 12234 4868 12258 4870
rect 12314 4868 12338 4870
rect 12394 4868 12400 4870
rect 12092 4859 12400 4868
rect 12092 3836 12400 3845
rect 12092 3834 12098 3836
rect 12154 3834 12178 3836
rect 12234 3834 12258 3836
rect 12314 3834 12338 3836
rect 12394 3834 12400 3836
rect 12154 3782 12156 3834
rect 12336 3782 12338 3834
rect 12092 3780 12098 3782
rect 12154 3780 12178 3782
rect 12234 3780 12258 3782
rect 12314 3780 12338 3782
rect 12394 3780 12400 3782
rect 12092 3771 12400 3780
rect 11072 2746 11376 2774
rect 12092 2748 12400 2757
rect 12092 2746 12098 2748
rect 12154 2746 12178 2748
rect 12234 2746 12258 2748
rect 12314 2746 12338 2748
rect 12394 2746 12400 2748
rect 11072 2650 11100 2746
rect 12154 2694 12156 2746
rect 12336 2694 12338 2746
rect 12092 2692 12098 2694
rect 12154 2692 12178 2694
rect 12234 2692 12258 2694
rect 12314 2692 12338 2694
rect 12394 2692 12400 2694
rect 12092 2683 12400 2692
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 12636 2446 12664 7482
rect 13096 6866 13124 7890
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 12752 6556 13060 6565
rect 12752 6554 12758 6556
rect 12814 6554 12838 6556
rect 12894 6554 12918 6556
rect 12974 6554 12998 6556
rect 13054 6554 13060 6556
rect 12814 6502 12816 6554
rect 12996 6502 12998 6554
rect 12752 6500 12758 6502
rect 12814 6500 12838 6502
rect 12894 6500 12918 6502
rect 12974 6500 12998 6502
rect 13054 6500 13060 6502
rect 12752 6491 13060 6500
rect 12752 5468 13060 5477
rect 12752 5466 12758 5468
rect 12814 5466 12838 5468
rect 12894 5466 12918 5468
rect 12974 5466 12998 5468
rect 13054 5466 13060 5468
rect 12814 5414 12816 5466
rect 12996 5414 12998 5466
rect 12752 5412 12758 5414
rect 12814 5412 12838 5414
rect 12894 5412 12918 5414
rect 12974 5412 12998 5414
rect 13054 5412 13060 5414
rect 12752 5403 13060 5412
rect 12752 4380 13060 4389
rect 12752 4378 12758 4380
rect 12814 4378 12838 4380
rect 12894 4378 12918 4380
rect 12974 4378 12998 4380
rect 13054 4378 13060 4380
rect 12814 4326 12816 4378
rect 12996 4326 12998 4378
rect 12752 4324 12758 4326
rect 12814 4324 12838 4326
rect 12894 4324 12918 4326
rect 12974 4324 12998 4326
rect 13054 4324 13060 4326
rect 12752 4315 13060 4324
rect 12752 3292 13060 3301
rect 12752 3290 12758 3292
rect 12814 3290 12838 3292
rect 12894 3290 12918 3292
rect 12974 3290 12998 3292
rect 13054 3290 13060 3292
rect 12814 3238 12816 3290
rect 12996 3238 12998 3290
rect 12752 3236 12758 3238
rect 12814 3236 12838 3238
rect 12894 3236 12918 3238
rect 12974 3236 12998 3238
rect 13054 3236 13060 3238
rect 12752 3227 13060 3236
rect 13280 2446 13308 10610
rect 13372 9654 13400 12582
rect 13464 12306 13492 14350
rect 13556 13394 13584 14826
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13648 12782 13676 14758
rect 14292 14618 14320 14758
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 13740 12866 13768 14554
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14200 14074 14228 14214
rect 14292 14074 14320 14554
rect 14568 14414 14596 14826
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14568 13326 14596 14350
rect 14660 13734 14688 14962
rect 14752 14414 14780 15438
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 14074 14780 14350
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14752 13326 14780 14010
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12918 14688 13126
rect 14648 12912 14700 12918
rect 13740 12850 14136 12866
rect 14648 12854 14700 12860
rect 13728 12844 14136 12850
rect 13780 12838 14136 12844
rect 13728 12786 13780 12792
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13556 12442 13584 12718
rect 13544 12436 13596 12442
rect 13924 12434 13952 12718
rect 13544 12378 13596 12384
rect 13832 12406 13952 12434
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13464 9450 13492 12242
rect 13556 11898 13584 12378
rect 13832 12238 13860 12406
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 11552 13596 11558
rect 13648 11540 13676 12174
rect 13596 11512 13676 11540
rect 13544 11494 13596 11500
rect 13556 11354 13584 11494
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13556 10538 13584 11290
rect 13832 11286 13860 12174
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13648 10742 13676 10950
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13464 9058 13492 9386
rect 13372 9030 13492 9058
rect 13372 8974 13400 9030
rect 13924 8974 13952 12038
rect 14016 11830 14044 12718
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 8498 13492 8774
rect 13924 8566 13952 8910
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 14016 2650 14044 10474
rect 14108 9586 14136 12838
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14464 12436 14516 12442
rect 14568 12434 14596 12718
rect 14516 12406 14596 12434
rect 14464 12378 14516 12384
rect 14660 12238 14688 12854
rect 15120 12850 15148 13262
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14936 12345 14964 12786
rect 14922 12336 14978 12345
rect 14922 12271 14978 12280
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15120 10810 15148 11018
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15304 10674 15332 15982
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15396 13258 15424 15914
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15706 15700 15846
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15856 15026 15884 16050
rect 16040 15638 16068 16050
rect 16028 15632 16080 15638
rect 16080 15580 16160 15586
rect 16028 15574 16160 15580
rect 16040 15558 16160 15574
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15764 14074 15792 14962
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13530 15516 13874
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15948 12986 15976 14962
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14482 16068 14758
rect 16028 14476 16080 14482
rect 16028 14418 16080 14424
rect 16132 14414 16160 15558
rect 16316 15042 16344 18090
rect 16500 17270 16528 18566
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16764 18080 16816 18086
rect 16764 18022 16816 18028
rect 16776 17864 16804 18022
rect 16960 17882 16988 18226
rect 16948 17876 17000 17882
rect 16776 17836 16896 17864
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16684 17678 16712 17750
rect 16868 17678 16896 17836
rect 16948 17818 17000 17824
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16592 17338 16620 17614
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16960 17202 16988 17818
rect 17052 17746 17080 19382
rect 17972 18834 18000 19926
rect 18432 19174 18460 21898
rect 18616 21842 18644 22510
rect 18708 22098 18736 22918
rect 18800 22778 18828 23598
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18892 22658 18920 23598
rect 18984 23050 19012 25434
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18972 22704 19024 22710
rect 18892 22652 18972 22658
rect 18892 22646 19024 22652
rect 18892 22630 19012 22646
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18800 22234 18828 22510
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 18892 22030 18920 22630
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 19076 22166 19104 22442
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18616 21814 18828 21842
rect 18800 21622 18828 21814
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 19168 21554 19196 22034
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18708 21010 18736 21286
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18892 19446 18920 19790
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 18432 18698 18460 19110
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17590 18320 17646 18329
rect 17408 18284 17460 18290
rect 17590 18255 17646 18264
rect 17408 18226 17460 18232
rect 17420 17746 17448 18226
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17512 17202 17540 18022
rect 17604 17542 17632 18255
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 16408 16674 16436 17138
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 16408 16646 16528 16674
rect 16224 15014 16344 15042
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16040 12986 16068 13806
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11354 15424 11630
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14384 9518 14412 9930
rect 15488 9586 15516 9998
rect 15764 9586 15792 10610
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 15212 8974 15240 9522
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15672 8634 15700 8978
rect 15856 8974 15884 9862
rect 15948 9654 15976 9862
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 15856 2446 15884 8910
rect 16132 2650 16160 13262
rect 16224 10062 16252 15014
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 14618 16344 14894
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16304 14408 16356 14414
rect 16500 14385 16528 16646
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16182 17080 16390
rect 17868 16244 17920 16250
rect 17972 16232 18000 16934
rect 18248 16250 18276 17002
rect 17920 16204 18000 16232
rect 18236 16244 18288 16250
rect 17868 16186 17920 16192
rect 18236 16186 18288 16192
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 14618 16620 16050
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16684 15026 16712 15438
rect 16960 15366 16988 15982
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17328 15094 17356 15506
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14618 16896 14758
rect 16960 14618 16988 14962
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 17328 14414 17356 15030
rect 17696 14958 17724 15846
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 18340 14550 18368 18566
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18708 17678 18736 18022
rect 18984 17814 19012 20470
rect 19168 20330 19196 21490
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 20602 19288 20742
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18358 19288 18702
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18984 17134 19012 17274
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18616 16726 18644 17070
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18984 16658 19012 17070
rect 19076 16658 19104 18294
rect 19352 17882 19380 29106
rect 19520 28860 19828 28869
rect 19520 28858 19526 28860
rect 19582 28858 19606 28860
rect 19662 28858 19686 28860
rect 19742 28858 19766 28860
rect 19822 28858 19828 28860
rect 19582 28806 19584 28858
rect 19764 28806 19766 28858
rect 19520 28804 19526 28806
rect 19582 28804 19606 28806
rect 19662 28804 19686 28806
rect 19742 28804 19766 28806
rect 19822 28804 19828 28806
rect 19520 28795 19828 28804
rect 19520 27772 19828 27781
rect 19520 27770 19526 27772
rect 19582 27770 19606 27772
rect 19662 27770 19686 27772
rect 19742 27770 19766 27772
rect 19822 27770 19828 27772
rect 19582 27718 19584 27770
rect 19764 27718 19766 27770
rect 19520 27716 19526 27718
rect 19582 27716 19606 27718
rect 19662 27716 19686 27718
rect 19742 27716 19766 27718
rect 19822 27716 19828 27718
rect 19520 27707 19828 27716
rect 19520 26684 19828 26693
rect 19520 26682 19526 26684
rect 19582 26682 19606 26684
rect 19662 26682 19686 26684
rect 19742 26682 19766 26684
rect 19822 26682 19828 26684
rect 19582 26630 19584 26682
rect 19764 26630 19766 26682
rect 19520 26628 19526 26630
rect 19582 26628 19606 26630
rect 19662 26628 19686 26630
rect 19742 26628 19766 26630
rect 19822 26628 19828 26630
rect 19520 26619 19828 26628
rect 19520 25596 19828 25605
rect 19520 25594 19526 25596
rect 19582 25594 19606 25596
rect 19662 25594 19686 25596
rect 19742 25594 19766 25596
rect 19822 25594 19828 25596
rect 19582 25542 19584 25594
rect 19764 25542 19766 25594
rect 19520 25540 19526 25542
rect 19582 25540 19606 25542
rect 19662 25540 19686 25542
rect 19742 25540 19766 25542
rect 19822 25540 19828 25542
rect 19520 25531 19828 25540
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 24886 19472 25094
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19520 24508 19828 24517
rect 19520 24506 19526 24508
rect 19582 24506 19606 24508
rect 19662 24506 19686 24508
rect 19742 24506 19766 24508
rect 19822 24506 19828 24508
rect 19582 24454 19584 24506
rect 19764 24454 19766 24506
rect 19520 24452 19526 24454
rect 19582 24452 19606 24454
rect 19662 24452 19686 24454
rect 19742 24452 19766 24454
rect 19822 24452 19828 24454
rect 19520 24443 19828 24452
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23186 19472 23666
rect 19520 23420 19828 23429
rect 19520 23418 19526 23420
rect 19582 23418 19606 23420
rect 19662 23418 19686 23420
rect 19742 23418 19766 23420
rect 19822 23418 19828 23420
rect 19582 23366 19584 23418
rect 19764 23366 19766 23418
rect 19520 23364 19526 23366
rect 19582 23364 19606 23366
rect 19662 23364 19686 23366
rect 19742 23364 19766 23366
rect 19822 23364 19828 23366
rect 19520 23355 19828 23364
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19520 22332 19828 22341
rect 19520 22330 19526 22332
rect 19582 22330 19606 22332
rect 19662 22330 19686 22332
rect 19742 22330 19766 22332
rect 19822 22330 19828 22332
rect 19582 22278 19584 22330
rect 19764 22278 19766 22330
rect 19520 22276 19526 22278
rect 19582 22276 19606 22278
rect 19662 22276 19686 22278
rect 19742 22276 19766 22278
rect 19822 22276 19828 22278
rect 19520 22267 19828 22276
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 19812 21434 19840 22034
rect 19904 21690 19932 29106
rect 20180 28316 20488 28325
rect 20180 28314 20186 28316
rect 20242 28314 20266 28316
rect 20322 28314 20346 28316
rect 20402 28314 20426 28316
rect 20482 28314 20488 28316
rect 20242 28262 20244 28314
rect 20424 28262 20426 28314
rect 20180 28260 20186 28262
rect 20242 28260 20266 28262
rect 20322 28260 20346 28262
rect 20402 28260 20426 28262
rect 20482 28260 20488 28262
rect 20180 28251 20488 28260
rect 20180 27228 20488 27237
rect 20180 27226 20186 27228
rect 20242 27226 20266 27228
rect 20322 27226 20346 27228
rect 20402 27226 20426 27228
rect 20482 27226 20488 27228
rect 20242 27174 20244 27226
rect 20424 27174 20426 27226
rect 20180 27172 20186 27174
rect 20242 27172 20266 27174
rect 20322 27172 20346 27174
rect 20402 27172 20426 27174
rect 20482 27172 20488 27174
rect 20180 27163 20488 27172
rect 20180 26140 20488 26149
rect 20180 26138 20186 26140
rect 20242 26138 20266 26140
rect 20322 26138 20346 26140
rect 20402 26138 20426 26140
rect 20482 26138 20488 26140
rect 20242 26086 20244 26138
rect 20424 26086 20426 26138
rect 20180 26084 20186 26086
rect 20242 26084 20266 26086
rect 20322 26084 20346 26086
rect 20402 26084 20426 26086
rect 20482 26084 20488 26086
rect 20180 26075 20488 26084
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25294 20116 25842
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20180 25052 20488 25061
rect 20180 25050 20186 25052
rect 20242 25050 20266 25052
rect 20322 25050 20346 25052
rect 20402 25050 20426 25052
rect 20482 25050 20488 25052
rect 20242 24998 20244 25050
rect 20424 24998 20426 25050
rect 20180 24996 20186 24998
rect 20242 24996 20266 24998
rect 20322 24996 20346 24998
rect 20402 24996 20426 24998
rect 20482 24996 20488 24998
rect 20180 24987 20488 24996
rect 20548 24954 20576 25162
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 19996 24206 20024 24550
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19996 23798 20024 24142
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19996 21690 20024 23734
rect 20088 23662 20116 24346
rect 20456 24342 20484 24550
rect 20640 24410 20668 24754
rect 20720 24744 20772 24750
rect 20720 24686 20772 24692
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20444 24336 20496 24342
rect 20732 24290 20760 24686
rect 20444 24278 20496 24284
rect 20640 24274 20760 24290
rect 20628 24268 20760 24274
rect 20680 24262 20760 24268
rect 20628 24210 20680 24216
rect 20720 24132 20772 24138
rect 20720 24074 20772 24080
rect 20180 23964 20488 23973
rect 20180 23962 20186 23964
rect 20242 23962 20266 23964
rect 20322 23962 20346 23964
rect 20402 23962 20426 23964
rect 20482 23962 20488 23964
rect 20242 23910 20244 23962
rect 20424 23910 20426 23962
rect 20180 23908 20186 23910
rect 20242 23908 20266 23910
rect 20322 23908 20346 23910
rect 20402 23908 20426 23910
rect 20482 23908 20488 23910
rect 20180 23899 20488 23908
rect 20732 23866 20760 24074
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 20352 23520 20404 23526
rect 20640 23474 20668 23802
rect 20352 23462 20404 23468
rect 20364 23118 20392 23462
rect 20456 23446 20760 23474
rect 20456 23118 20484 23446
rect 20732 23186 20760 23446
rect 20720 23180 20772 23186
rect 20720 23122 20772 23128
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20180 22876 20488 22885
rect 20180 22874 20186 22876
rect 20242 22874 20266 22876
rect 20322 22874 20346 22876
rect 20402 22874 20426 22876
rect 20482 22874 20488 22876
rect 20242 22822 20244 22874
rect 20424 22822 20426 22874
rect 20180 22820 20186 22822
rect 20242 22820 20266 22822
rect 20322 22820 20346 22822
rect 20402 22820 20426 22822
rect 20482 22820 20488 22822
rect 20180 22811 20488 22820
rect 20548 22778 20576 22918
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 20088 22094 20116 22374
rect 20548 22234 20576 22578
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20088 22066 20208 22094
rect 20180 22030 20208 22066
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19984 21684 20036 21690
rect 20088 21672 20116 21966
rect 20180 21788 20488 21797
rect 20180 21786 20186 21788
rect 20242 21786 20266 21788
rect 20322 21786 20346 21788
rect 20402 21786 20426 21788
rect 20482 21786 20488 21788
rect 20242 21734 20244 21786
rect 20424 21734 20426 21786
rect 20180 21732 20186 21734
rect 20242 21732 20266 21734
rect 20322 21732 20346 21734
rect 20402 21732 20426 21734
rect 20482 21732 20488 21734
rect 20180 21723 20488 21732
rect 20168 21684 20220 21690
rect 20088 21644 20168 21672
rect 19984 21626 20036 21632
rect 20168 21626 20220 21632
rect 20548 21554 20576 21966
rect 20732 21962 20760 23122
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 19444 21418 19840 21434
rect 19904 21418 19932 21490
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19444 21412 19852 21418
rect 19444 21406 19800 21412
rect 19444 21026 19472 21406
rect 19800 21354 19852 21360
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19520 21244 19828 21253
rect 19520 21242 19526 21244
rect 19582 21242 19606 21244
rect 19662 21242 19686 21244
rect 19742 21242 19766 21244
rect 19822 21242 19828 21244
rect 19582 21190 19584 21242
rect 19764 21190 19766 21242
rect 19520 21188 19526 21190
rect 19582 21188 19606 21190
rect 19662 21188 19686 21190
rect 19742 21188 19766 21190
rect 19822 21188 19828 21190
rect 19520 21179 19828 21188
rect 19444 20998 19564 21026
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20466 19472 20878
rect 19536 20602 19564 20998
rect 19904 20942 19932 21354
rect 19996 20942 20024 21422
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19444 19802 19472 20402
rect 19520 20156 19828 20165
rect 19520 20154 19526 20156
rect 19582 20154 19606 20156
rect 19662 20154 19686 20156
rect 19742 20154 19766 20156
rect 19822 20154 19828 20156
rect 19582 20102 19584 20154
rect 19764 20102 19766 20154
rect 19520 20100 19526 20102
rect 19582 20100 19606 20102
rect 19662 20100 19686 20102
rect 19742 20100 19766 20102
rect 19822 20100 19828 20102
rect 19520 20091 19828 20100
rect 19444 19774 19564 19802
rect 19536 19446 19564 19774
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19444 18970 19472 19382
rect 19520 19068 19828 19077
rect 19520 19066 19526 19068
rect 19582 19066 19606 19068
rect 19662 19066 19686 19068
rect 19742 19066 19766 19068
rect 19822 19066 19828 19068
rect 19582 19014 19584 19066
rect 19764 19014 19766 19066
rect 19520 19012 19526 19014
rect 19582 19012 19606 19014
rect 19662 19012 19686 19014
rect 19742 19012 19766 19014
rect 19822 19012 19828 19014
rect 19520 19003 19828 19012
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19904 18630 19932 20878
rect 19996 20602 20024 20878
rect 20088 20602 20116 21286
rect 20364 21146 20392 21490
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20180 20700 20488 20709
rect 20180 20698 20186 20700
rect 20242 20698 20266 20700
rect 20322 20698 20346 20700
rect 20402 20698 20426 20700
rect 20482 20698 20488 20700
rect 20242 20646 20244 20698
rect 20424 20646 20426 20698
rect 20180 20644 20186 20646
rect 20242 20644 20266 20646
rect 20322 20644 20346 20646
rect 20402 20644 20426 20646
rect 20482 20644 20488 20646
rect 20180 20635 20488 20644
rect 20824 20602 20852 29106
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21192 25226 21220 25638
rect 21180 25220 21232 25226
rect 21180 25162 21232 25168
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21376 24818 21404 25094
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 20904 24268 20956 24274
rect 21088 24268 21140 24274
rect 20956 24228 21036 24256
rect 20904 24210 20956 24216
rect 21008 24070 21036 24228
rect 21088 24210 21140 24216
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20904 23860 20956 23866
rect 21100 23848 21128 24210
rect 21376 24138 21404 24754
rect 21836 24410 21864 24754
rect 21916 24608 21968 24614
rect 21916 24550 21968 24556
rect 21928 24410 21956 24550
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 20956 23820 21128 23848
rect 20904 23802 20956 23808
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20916 23526 20944 23666
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 20904 23520 20956 23526
rect 20904 23462 20956 23468
rect 21192 23118 21220 23530
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 21088 22976 21140 22982
rect 21088 22918 21140 22924
rect 21100 22710 21128 22918
rect 21088 22704 21140 22710
rect 20994 22672 21050 22681
rect 21088 22646 21140 22652
rect 20994 22607 20996 22616
rect 21048 22607 21050 22616
rect 20996 22578 21048 22584
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20916 22438 20944 22510
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20916 21146 20944 21898
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21690 21036 21830
rect 21100 21690 21128 22646
rect 21192 22030 21220 23054
rect 21284 22778 21312 24074
rect 21376 23526 21404 24074
rect 21468 23730 21496 24074
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 23520 21416 23526
rect 21364 23462 21416 23468
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 21008 21298 21036 21490
rect 21100 21418 21128 21626
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21192 21298 21220 21966
rect 21284 21690 21312 22578
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21468 22234 21496 22510
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21560 22030 21588 23462
rect 21744 22778 21772 24142
rect 22112 23202 22140 29106
rect 26948 28860 27256 28869
rect 26948 28858 26954 28860
rect 27010 28858 27034 28860
rect 27090 28858 27114 28860
rect 27170 28858 27194 28860
rect 27250 28858 27256 28860
rect 27010 28806 27012 28858
rect 27192 28806 27194 28858
rect 26948 28804 26954 28806
rect 27010 28804 27034 28806
rect 27090 28804 27114 28806
rect 27170 28804 27194 28806
rect 27250 28804 27256 28806
rect 26948 28795 27256 28804
rect 27608 28316 27916 28325
rect 27608 28314 27614 28316
rect 27670 28314 27694 28316
rect 27750 28314 27774 28316
rect 27830 28314 27854 28316
rect 27910 28314 27916 28316
rect 27670 28262 27672 28314
rect 27852 28262 27854 28314
rect 27608 28260 27614 28262
rect 27670 28260 27694 28262
rect 27750 28260 27774 28262
rect 27830 28260 27854 28262
rect 27910 28260 27916 28262
rect 27608 28251 27916 28260
rect 26948 27772 27256 27781
rect 26948 27770 26954 27772
rect 27010 27770 27034 27772
rect 27090 27770 27114 27772
rect 27170 27770 27194 27772
rect 27250 27770 27256 27772
rect 27010 27718 27012 27770
rect 27192 27718 27194 27770
rect 26948 27716 26954 27718
rect 27010 27716 27034 27718
rect 27090 27716 27114 27718
rect 27170 27716 27194 27718
rect 27250 27716 27256 27718
rect 26948 27707 27256 27716
rect 27608 27228 27916 27237
rect 27608 27226 27614 27228
rect 27670 27226 27694 27228
rect 27750 27226 27774 27228
rect 27830 27226 27854 27228
rect 27910 27226 27916 27228
rect 27670 27174 27672 27226
rect 27852 27174 27854 27226
rect 27608 27172 27614 27174
rect 27670 27172 27694 27174
rect 27750 27172 27774 27174
rect 27830 27172 27854 27174
rect 27910 27172 27916 27174
rect 27608 27163 27916 27172
rect 26948 26684 27256 26693
rect 26948 26682 26954 26684
rect 27010 26682 27034 26684
rect 27090 26682 27114 26684
rect 27170 26682 27194 26684
rect 27250 26682 27256 26684
rect 27010 26630 27012 26682
rect 27192 26630 27194 26682
rect 26948 26628 26954 26630
rect 27010 26628 27034 26630
rect 27090 26628 27114 26630
rect 27170 26628 27194 26630
rect 27250 26628 27256 26630
rect 26948 26619 27256 26628
rect 27608 26140 27916 26149
rect 27608 26138 27614 26140
rect 27670 26138 27694 26140
rect 27750 26138 27774 26140
rect 27830 26138 27854 26140
rect 27910 26138 27916 26140
rect 27670 26086 27672 26138
rect 27852 26086 27854 26138
rect 27608 26084 27614 26086
rect 27670 26084 27694 26086
rect 27750 26084 27774 26086
rect 27830 26084 27854 26086
rect 27910 26084 27916 26086
rect 27608 26075 27916 26084
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22296 24614 22324 25094
rect 22572 24954 22600 25094
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22376 24812 22428 24818
rect 22756 24800 22784 25842
rect 26948 25596 27256 25605
rect 26948 25594 26954 25596
rect 27010 25594 27034 25596
rect 27090 25594 27114 25596
rect 27170 25594 27194 25596
rect 27250 25594 27256 25596
rect 27010 25542 27012 25594
rect 27192 25542 27194 25594
rect 26948 25540 26954 25542
rect 27010 25540 27034 25542
rect 27090 25540 27114 25542
rect 27170 25540 27194 25542
rect 27250 25540 27256 25542
rect 26948 25531 27256 25540
rect 24216 25356 24268 25362
rect 24216 25298 24268 25304
rect 22836 25220 22888 25226
rect 22836 25162 22888 25168
rect 22848 24954 22876 25162
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 22836 24812 22888 24818
rect 22756 24772 22836 24800
rect 22376 24754 22428 24760
rect 22836 24754 22888 24760
rect 24124 24812 24176 24818
rect 24228 24800 24256 25298
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 24688 24954 24716 25162
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 24176 24772 24256 24800
rect 24124 24754 24176 24760
rect 22284 24608 22336 24614
rect 22284 24550 22336 24556
rect 22296 24206 22324 24550
rect 22388 24410 22416 24754
rect 22848 24410 22876 24754
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23216 24614 23244 24686
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 23798 22324 24142
rect 23308 24138 23336 24550
rect 23664 24336 23716 24342
rect 23664 24278 23716 24284
rect 23296 24132 23348 24138
rect 23296 24074 23348 24080
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 22284 23792 22336 23798
rect 22284 23734 22336 23740
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22204 23322 22232 23530
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22296 23202 22324 23734
rect 23032 23594 23060 24006
rect 23400 23798 23428 24006
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23492 23730 23520 24006
rect 23676 23730 23704 24278
rect 23480 23724 23532 23730
rect 23664 23724 23716 23730
rect 23532 23684 23612 23712
rect 23480 23666 23532 23672
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 22020 23186 22140 23202
rect 22008 23180 22140 23186
rect 22060 23174 22140 23180
rect 22204 23174 22324 23202
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 22008 23122 22060 23128
rect 22204 22930 22232 23174
rect 22112 22902 22232 22930
rect 22284 22976 22336 22982
rect 22336 22924 22600 22930
rect 22284 22918 22600 22924
rect 22296 22902 22600 22918
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22008 22568 22060 22574
rect 22006 22536 22008 22545
rect 22060 22536 22062 22545
rect 22006 22471 22062 22480
rect 22112 22030 22140 22902
rect 22572 22778 22600 22902
rect 22560 22772 22612 22778
rect 22560 22714 22612 22720
rect 23204 22704 23256 22710
rect 22558 22672 22614 22681
rect 22284 22636 22336 22642
rect 23204 22646 23256 22652
rect 22558 22607 22560 22616
rect 22284 22578 22336 22584
rect 22612 22607 22614 22616
rect 22560 22578 22612 22584
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22204 22114 22232 22442
rect 22296 22234 22324 22578
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22204 22086 22324 22114
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21560 21622 21588 21966
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21008 21270 21220 21298
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 22112 20942 22140 21966
rect 22296 21418 22324 22086
rect 22756 22094 22784 22510
rect 23216 22506 23244 22646
rect 23400 22642 23428 23190
rect 23492 23118 23520 23462
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23584 22760 23612 23684
rect 23664 23666 23716 23672
rect 23676 23322 23704 23666
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23492 22732 23612 22760
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23204 22500 23256 22506
rect 23204 22442 23256 22448
rect 23216 22098 23244 22442
rect 22756 22066 22876 22094
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22204 21146 22232 21286
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22388 21010 22416 21558
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22664 21146 22692 21490
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22744 21004 22796 21010
rect 22744 20946 22796 20952
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20088 20466 20116 20538
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19996 20346 20024 20402
rect 19996 20318 20116 20346
rect 20088 20262 20116 20318
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 19996 19786 20024 20198
rect 21008 20058 21036 20198
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20824 19786 20852 19994
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20180 19612 20488 19621
rect 20180 19610 20186 19612
rect 20242 19610 20266 19612
rect 20322 19610 20346 19612
rect 20402 19610 20426 19612
rect 20482 19610 20488 19612
rect 20242 19558 20244 19610
rect 20424 19558 20426 19610
rect 20180 19556 20186 19558
rect 20242 19556 20266 19558
rect 20322 19556 20346 19558
rect 20402 19556 20426 19558
rect 20482 19556 20488 19558
rect 20180 19547 20488 19556
rect 20916 19514 20944 19790
rect 20904 19508 20956 19514
rect 20904 19450 20956 19456
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 18290 19932 18566
rect 20088 18426 20116 18838
rect 20916 18834 20944 19246
rect 21008 18834 21036 19994
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21376 18970 21404 19722
rect 21836 19514 21864 19722
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21456 18896 21508 18902
rect 21456 18838 21508 18844
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 20180 18524 20488 18533
rect 20180 18522 20186 18524
rect 20242 18522 20266 18524
rect 20322 18522 20346 18524
rect 20402 18522 20426 18524
rect 20482 18522 20488 18524
rect 20242 18470 20244 18522
rect 20424 18470 20426 18522
rect 20180 18468 20186 18470
rect 20242 18468 20266 18470
rect 20322 18468 20346 18470
rect 20402 18468 20426 18470
rect 20482 18468 20488 18470
rect 20180 18459 20488 18468
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19520 17980 19828 17989
rect 19520 17978 19526 17980
rect 19582 17978 19606 17980
rect 19662 17978 19686 17980
rect 19742 17978 19766 17980
rect 19822 17978 19828 17980
rect 19582 17926 19584 17978
rect 19764 17926 19766 17978
rect 19520 17924 19526 17926
rect 19582 17924 19606 17926
rect 19662 17924 19686 17926
rect 19742 17924 19766 17926
rect 19822 17924 19828 17926
rect 19520 17915 19828 17924
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 19812 17598 20024 17626
rect 19812 17542 19840 17598
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 18432 15706 18460 15914
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18604 14952 18656 14958
rect 18604 14894 18656 14900
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 17316 14408 17368 14414
rect 16304 14350 16356 14356
rect 16486 14376 16542 14385
rect 16316 13530 16344 14350
rect 18340 14362 18368 14486
rect 17316 14350 17368 14356
rect 16486 14311 16542 14320
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16302 12744 16358 12753
rect 16302 12679 16358 12688
rect 16316 12646 16344 12679
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12442 16344 12582
rect 16304 12436 16356 12442
rect 16500 12434 16528 14311
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16960 12918 16988 13670
rect 17052 13258 17080 14214
rect 17328 14074 17356 14350
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 18248 14334 18368 14362
rect 17604 14074 17632 14282
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13530 17172 13670
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17328 13326 17356 14010
rect 18248 13938 18276 14334
rect 17776 13932 17828 13938
rect 17776 13874 17828 13880
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 17052 12442 17080 13194
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 17144 12850 17172 13126
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17236 12442 17264 12786
rect 17040 12436 17092 12442
rect 16500 12406 16620 12434
rect 16304 12378 16356 12384
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11150 16344 12038
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16224 9722 16252 9998
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 8634 16344 9998
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16408 2774 16436 11562
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11218 16528 11494
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16592 10062 16620 12406
rect 17040 12378 17092 12384
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17052 12170 17080 12378
rect 17040 12164 17092 12170
rect 17040 12106 17092 12112
rect 17236 12102 17264 12378
rect 17420 12238 17448 13262
rect 17788 13258 17816 13874
rect 17776 13252 17828 13258
rect 17696 13212 17776 13240
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17696 11898 17724 13212
rect 17776 13194 17828 13200
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17696 11762 17724 11834
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17052 11540 17080 11698
rect 17224 11552 17276 11558
rect 17052 11512 17224 11540
rect 17224 11494 17276 11500
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 7954 16620 9998
rect 17420 9926 17448 10610
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16960 6798 16988 9522
rect 17052 9178 17080 9522
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 17144 9110 17172 9862
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 17144 8906 17172 9046
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 7478 17080 7686
rect 17040 7472 17092 7478
rect 17040 7414 17092 7420
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16408 2746 16528 2774
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16500 2446 16528 2746
rect 17144 2650 17172 8842
rect 17236 8498 17264 9046
rect 17328 8974 17356 9590
rect 17420 9518 17448 9862
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17420 8430 17448 8910
rect 17512 8634 17540 8910
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17604 8090 17632 11290
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17696 7886 17724 9862
rect 17788 9654 17816 12378
rect 18064 12374 18092 12786
rect 18156 12646 18184 13194
rect 18616 12986 18644 14894
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18708 12646 18736 16594
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 19076 16114 19104 16458
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 15162 18920 15438
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18972 14272 19024 14278
rect 19076 14260 19104 16050
rect 19168 15026 19196 16934
rect 19352 16794 19380 17206
rect 19520 16892 19828 16901
rect 19520 16890 19526 16892
rect 19582 16890 19606 16892
rect 19662 16890 19686 16892
rect 19742 16890 19766 16892
rect 19822 16890 19828 16892
rect 19582 16838 19584 16890
rect 19764 16838 19766 16890
rect 19520 16836 19526 16838
rect 19582 16836 19606 16838
rect 19662 16836 19686 16838
rect 19742 16836 19766 16838
rect 19822 16836 19828 16838
rect 19520 16827 19828 16836
rect 19904 16794 19932 17478
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 19168 14618 19196 14962
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19260 14414 19288 16730
rect 19996 16658 20024 17598
rect 20088 17338 20116 18090
rect 20364 17746 20392 18362
rect 21100 18358 21128 18702
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18426 21312 18566
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 20180 17436 20488 17445
rect 20180 17434 20186 17436
rect 20242 17434 20266 17436
rect 20322 17434 20346 17436
rect 20402 17434 20426 17436
rect 20482 17434 20488 17436
rect 20242 17382 20244 17434
rect 20424 17382 20426 17434
rect 20180 17380 20186 17382
rect 20242 17380 20266 17382
rect 20322 17380 20346 17382
rect 20402 17380 20426 17382
rect 20482 17380 20488 17382
rect 20180 17371 20488 17380
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 20180 16590 20208 16934
rect 20732 16794 20760 18226
rect 21100 17882 21128 18294
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 20996 17604 21048 17610
rect 20996 17546 21048 17552
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20180 16348 20488 16357
rect 20180 16346 20186 16348
rect 20242 16346 20266 16348
rect 20322 16346 20346 16348
rect 20402 16346 20426 16348
rect 20482 16346 20488 16348
rect 20242 16294 20244 16346
rect 20424 16294 20426 16346
rect 20180 16292 20186 16294
rect 20242 16292 20266 16294
rect 20322 16292 20346 16294
rect 20402 16292 20426 16294
rect 20482 16292 20488 16294
rect 20180 16283 20488 16292
rect 20548 16250 20576 16526
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20640 16130 20668 16594
rect 20732 16250 20760 16730
rect 20916 16726 20944 16934
rect 21008 16726 21036 17546
rect 21284 17134 21312 18226
rect 21468 17882 21496 18838
rect 21928 18766 21956 19110
rect 22112 18834 22140 19858
rect 22204 19446 22232 20810
rect 22756 20466 22784 20946
rect 22848 20874 22876 22066
rect 23204 22092 23256 22098
rect 23204 22034 23256 22040
rect 23400 22030 23428 22578
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23400 21690 23428 21966
rect 23492 21894 23520 22732
rect 23768 22234 23796 24686
rect 24136 24070 24164 24754
rect 24872 24070 24900 25094
rect 25240 24954 25268 25162
rect 27608 25052 27916 25061
rect 27608 25050 27614 25052
rect 27670 25050 27694 25052
rect 27750 25050 27774 25052
rect 27830 25050 27854 25052
rect 27910 25050 27916 25052
rect 27670 24998 27672 25050
rect 27852 24998 27854 25050
rect 27608 24996 27614 24998
rect 27670 24996 27694 24998
rect 27750 24996 27774 24998
rect 27830 24996 27854 24998
rect 27910 24996 27916 24998
rect 27608 24987 27916 24996
rect 25228 24948 25280 24954
rect 25228 24890 25280 24896
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25148 24342 25176 24754
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25136 24336 25188 24342
rect 25136 24278 25188 24284
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24136 23866 24164 24006
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24136 23662 24164 23802
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24032 23656 24084 23662
rect 24032 23598 24084 23604
rect 24124 23656 24176 23662
rect 24124 23598 24176 23604
rect 23952 23322 23980 23598
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 23860 22234 23888 23054
rect 24044 22710 24072 23598
rect 24124 23520 24176 23526
rect 24124 23462 24176 23468
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 24030 22536 24086 22545
rect 24030 22471 24086 22480
rect 24044 22438 24072 22471
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 24044 22030 24072 22374
rect 24136 22030 24164 23462
rect 24504 23118 24532 24006
rect 24872 23474 24900 24006
rect 24964 23866 24992 24142
rect 25516 24070 25544 24210
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25516 23866 25544 24006
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25504 23860 25556 23866
rect 25504 23802 25556 23808
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 24780 23446 24900 23474
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23492 21622 23520 21830
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 23860 21146 23888 21966
rect 24584 21956 24636 21962
rect 24584 21898 24636 21904
rect 24596 21690 24624 21898
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23952 20942 23980 21490
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24412 20942 24440 21286
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 22836 20868 22888 20874
rect 22836 20810 22888 20816
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 22940 20534 22968 20810
rect 23124 20602 23152 20810
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 22928 20528 22980 20534
rect 22928 20470 22980 20476
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22388 20058 22416 20402
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 23032 19854 23060 20334
rect 23308 20058 23336 20334
rect 24044 20058 24072 20470
rect 24504 20398 24532 21490
rect 24596 20874 24624 21490
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 24676 20868 24728 20874
rect 24676 20810 24728 20816
rect 24688 20534 24716 20810
rect 24676 20528 24728 20534
rect 24676 20470 24728 20476
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24688 19854 24716 20198
rect 24780 20058 24808 23446
rect 25424 23322 25452 23598
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24872 22574 24900 22986
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 24872 22030 24900 22510
rect 24964 22438 24992 22986
rect 25516 22574 25544 23802
rect 25608 23662 25636 24550
rect 25976 23730 26004 24754
rect 26948 24508 27256 24517
rect 26948 24506 26954 24508
rect 27010 24506 27034 24508
rect 27090 24506 27114 24508
rect 27170 24506 27194 24508
rect 27250 24506 27256 24508
rect 27010 24454 27012 24506
rect 27192 24454 27194 24506
rect 26948 24452 26954 24454
rect 27010 24452 27034 24454
rect 27090 24452 27114 24454
rect 27170 24452 27194 24454
rect 27250 24452 27256 24454
rect 26948 24443 27256 24452
rect 26056 24132 26108 24138
rect 26056 24074 26108 24080
rect 26068 23866 26096 24074
rect 27608 23964 27916 23973
rect 27608 23962 27614 23964
rect 27670 23962 27694 23964
rect 27750 23962 27774 23964
rect 27830 23962 27854 23964
rect 27910 23962 27916 23964
rect 27670 23910 27672 23962
rect 27852 23910 27854 23962
rect 27608 23908 27614 23910
rect 27670 23908 27694 23910
rect 27750 23908 27774 23910
rect 27830 23908 27854 23910
rect 27910 23908 27916 23910
rect 27608 23899 27916 23908
rect 26056 23860 26108 23866
rect 26056 23802 26108 23808
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 25596 23656 25648 23662
rect 25596 23598 25648 23604
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25608 22642 25636 22918
rect 25884 22778 25912 23054
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25504 22568 25556 22574
rect 25504 22510 25556 22516
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 25516 22094 25544 22510
rect 25332 22066 25544 22094
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25056 21690 25084 21966
rect 25044 21684 25096 21690
rect 25044 21626 25096 21632
rect 25332 21622 25360 22066
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24872 21078 24900 21490
rect 24860 21072 24912 21078
rect 24860 21014 24912 21020
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20398 24900 20810
rect 25608 20534 25636 22578
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20602 25728 20742
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25596 20528 25648 20534
rect 25596 20470 25648 20476
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24872 20058 24900 20198
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 22928 19712 22980 19718
rect 22928 19654 22980 19660
rect 22940 19514 22968 19654
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 22376 18692 22428 18698
rect 22376 18634 22428 18640
rect 22388 18426 22416 18634
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 21456 17876 21508 17882
rect 21456 17818 21508 17824
rect 22572 17338 22600 18226
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 22008 17128 22060 17134
rect 22060 17076 22140 17082
rect 22008 17070 22140 17076
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 20812 16584 20864 16590
rect 20810 16552 20812 16561
rect 20904 16584 20956 16590
rect 20864 16552 20866 16561
rect 20904 16526 20956 16532
rect 20810 16487 20866 16496
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20640 16102 20760 16130
rect 20732 15910 20760 16102
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 19520 15804 19828 15813
rect 19520 15802 19526 15804
rect 19582 15802 19606 15804
rect 19662 15802 19686 15804
rect 19742 15802 19766 15804
rect 19822 15802 19828 15804
rect 19582 15750 19584 15802
rect 19764 15750 19766 15802
rect 19520 15748 19526 15750
rect 19582 15748 19606 15750
rect 19662 15748 19686 15750
rect 19742 15748 19766 15750
rect 19822 15748 19828 15750
rect 19520 15739 19828 15748
rect 20916 15434 20944 16526
rect 21008 16182 21036 16662
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 21100 15910 21128 16186
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21284 15502 21312 17070
rect 22020 17054 22140 17070
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 20904 15428 20956 15434
rect 20904 15370 20956 15376
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 19352 15094 19380 15302
rect 20180 15260 20488 15269
rect 20180 15258 20186 15260
rect 20242 15258 20266 15260
rect 20322 15258 20346 15260
rect 20402 15258 20426 15260
rect 20482 15258 20488 15260
rect 20242 15206 20244 15258
rect 20424 15206 20426 15258
rect 20180 15204 20186 15206
rect 20242 15204 20266 15206
rect 20322 15204 20346 15206
rect 20402 15204 20426 15206
rect 20482 15204 20488 15206
rect 20180 15195 20488 15204
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20444 14884 20496 14890
rect 20444 14826 20496 14832
rect 19520 14716 19828 14725
rect 19520 14714 19526 14716
rect 19582 14714 19606 14716
rect 19662 14714 19686 14716
rect 19742 14714 19766 14716
rect 19822 14714 19828 14716
rect 19582 14662 19584 14714
rect 19764 14662 19766 14714
rect 19520 14660 19526 14662
rect 19582 14660 19606 14662
rect 19662 14660 19686 14662
rect 19742 14660 19766 14662
rect 19822 14660 19828 14662
rect 19520 14651 19828 14660
rect 20456 14550 20484 14826
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19076 14232 19288 14260
rect 18972 14214 19024 14220
rect 18800 14006 18828 14214
rect 18984 14074 19012 14214
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18800 13870 18828 13942
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12434 18736 12582
rect 18248 12406 18736 12434
rect 18052 12368 18104 12374
rect 18248 12345 18276 12406
rect 18234 12336 18290 12345
rect 18052 12310 18104 12316
rect 18156 12294 18234 12322
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17880 11898 17908 12106
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17776 9648 17828 9654
rect 17776 9590 17828 9596
rect 17972 8498 18000 10610
rect 18156 9926 18184 12294
rect 18892 12306 18920 13874
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12986 19012 13126
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19076 12850 19104 13330
rect 19168 13326 19196 13670
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19260 12866 19288 14232
rect 19352 13002 19380 14282
rect 19444 13802 19472 14418
rect 20180 14172 20488 14181
rect 20180 14170 20186 14172
rect 20242 14170 20266 14172
rect 20322 14170 20346 14172
rect 20402 14170 20426 14172
rect 20482 14170 20488 14172
rect 20242 14118 20244 14170
rect 20424 14118 20426 14170
rect 20180 14116 20186 14118
rect 20242 14116 20266 14118
rect 20322 14116 20346 14118
rect 20402 14116 20426 14118
rect 20482 14116 20488 14118
rect 20180 14107 20488 14116
rect 20548 14074 20576 14962
rect 20732 14822 20760 14962
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14414 20760 14758
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20824 14346 20852 15302
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 20732 13716 20760 14214
rect 20824 14006 20852 14282
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20640 13688 20760 13716
rect 19520 13628 19828 13637
rect 19520 13626 19526 13628
rect 19582 13626 19606 13628
rect 19662 13626 19686 13628
rect 19742 13626 19766 13628
rect 19822 13626 19828 13628
rect 19582 13574 19584 13626
rect 19764 13574 19766 13626
rect 19520 13572 19526 13574
rect 19582 13572 19606 13574
rect 19662 13572 19686 13574
rect 19742 13572 19766 13574
rect 19822 13572 19828 13574
rect 19520 13563 19828 13572
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20180 13084 20488 13093
rect 20180 13082 20186 13084
rect 20242 13082 20266 13084
rect 20322 13082 20346 13084
rect 20402 13082 20426 13084
rect 20482 13082 20488 13084
rect 20242 13030 20244 13082
rect 20424 13030 20426 13082
rect 20180 13028 20186 13030
rect 20242 13028 20266 13030
rect 20322 13028 20346 13030
rect 20402 13028 20426 13030
rect 20482 13028 20488 13030
rect 20180 13019 20488 13028
rect 19352 12986 19472 13002
rect 20548 12986 20576 13194
rect 20640 13190 20668 13688
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 19352 12980 19484 12986
rect 19352 12974 19432 12980
rect 19432 12922 19484 12928
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19156 12844 19208 12850
rect 19260 12838 19472 12866
rect 19156 12786 19208 12792
rect 18234 12271 18290 12280
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11830 18552 12038
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10266 18276 10406
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18236 10056 18288 10062
rect 18340 10044 18368 11766
rect 18892 11762 18920 12242
rect 19076 11778 19104 12786
rect 19168 12646 19196 12786
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19352 12306 19380 12718
rect 19444 12714 19472 12838
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 19520 12540 19828 12549
rect 19520 12538 19526 12540
rect 19582 12538 19606 12540
rect 19662 12538 19686 12540
rect 19742 12538 19766 12540
rect 19822 12538 19828 12540
rect 19582 12486 19584 12538
rect 19764 12486 19766 12538
rect 19520 12484 19526 12486
rect 19582 12484 19606 12486
rect 19662 12484 19686 12486
rect 19742 12484 19766 12486
rect 19822 12484 19828 12486
rect 19520 12475 19828 12484
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19260 11778 19288 11834
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18880 11756 18932 11762
rect 19076 11750 19288 11778
rect 18880 11698 18932 11704
rect 18432 11150 18460 11698
rect 18788 11688 18840 11694
rect 19064 11688 19116 11694
rect 18840 11636 18920 11642
rect 18788 11630 18920 11636
rect 19064 11630 19116 11636
rect 18800 11614 18920 11630
rect 18892 11558 18920 11614
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18880 11552 18932 11558
rect 18880 11494 18932 11500
rect 18800 11150 18828 11494
rect 18892 11150 18920 11494
rect 19076 11354 19104 11630
rect 19352 11626 19380 12038
rect 19904 11830 19932 12038
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19536 11558 19564 11698
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19444 11218 19472 11494
rect 19520 11452 19828 11461
rect 19520 11450 19526 11452
rect 19582 11450 19606 11452
rect 19662 11450 19686 11452
rect 19742 11450 19766 11452
rect 19822 11450 19828 11452
rect 19582 11398 19584 11450
rect 19764 11398 19766 11450
rect 19520 11396 19526 11398
rect 19582 11396 19606 11398
rect 19662 11396 19686 11398
rect 19742 11396 19766 11398
rect 19822 11396 19828 11398
rect 19520 11387 19828 11396
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18432 10810 18460 11086
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18800 10606 18828 11086
rect 18788 10600 18840 10606
rect 18788 10542 18840 10548
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18800 10266 18828 10406
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18288 10016 18368 10044
rect 18236 9998 18288 10004
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18064 9042 18092 9658
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18340 9178 18368 9454
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17880 7886 17908 8434
rect 17972 7954 18000 8434
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17972 7732 18000 7890
rect 18248 7818 18276 8774
rect 18616 8090 18644 8842
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 17880 7704 18000 7732
rect 17880 2650 17908 7704
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18064 6866 18092 7346
rect 18432 7206 18460 7822
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 18432 2446 18460 7142
rect 18892 2774 18920 11086
rect 19520 10364 19828 10373
rect 19520 10362 19526 10364
rect 19582 10362 19606 10364
rect 19662 10362 19686 10364
rect 19742 10362 19766 10364
rect 19822 10362 19828 10364
rect 19582 10310 19584 10362
rect 19764 10310 19766 10362
rect 19520 10308 19526 10310
rect 19582 10308 19606 10310
rect 19662 10308 19686 10310
rect 19742 10308 19766 10310
rect 19822 10308 19828 10310
rect 19520 10299 19828 10308
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18984 9178 19012 9386
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18984 8974 19012 9114
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19352 8022 19380 10202
rect 19798 10160 19854 10169
rect 19798 10095 19800 10104
rect 19852 10095 19854 10104
rect 19800 10066 19852 10072
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9586 19748 9998
rect 19904 9722 19932 11766
rect 20088 11694 20116 12650
rect 20442 12200 20498 12209
rect 20442 12135 20444 12144
rect 20496 12135 20498 12144
rect 20444 12106 20496 12112
rect 20180 11996 20488 12005
rect 20180 11994 20186 11996
rect 20242 11994 20266 11996
rect 20322 11994 20346 11996
rect 20402 11994 20426 11996
rect 20482 11994 20488 11996
rect 20242 11942 20244 11994
rect 20424 11942 20426 11994
rect 20180 11940 20186 11942
rect 20242 11940 20266 11942
rect 20322 11940 20346 11942
rect 20402 11940 20426 11942
rect 20482 11940 20488 11942
rect 20180 11931 20488 11940
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19444 8974 19472 9386
rect 19520 9276 19828 9285
rect 19520 9274 19526 9276
rect 19582 9274 19606 9276
rect 19662 9274 19686 9276
rect 19742 9274 19766 9276
rect 19822 9274 19828 9276
rect 19582 9222 19584 9274
rect 19764 9222 19766 9274
rect 19520 9220 19526 9222
rect 19582 9220 19606 9222
rect 19662 9220 19686 9222
rect 19742 9220 19766 9222
rect 19822 9220 19828 9222
rect 19520 9211 19828 9220
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19444 8838 19472 8910
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19904 8634 19932 8774
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19996 8514 20024 10406
rect 20088 10198 20116 11630
rect 20180 10908 20488 10917
rect 20180 10906 20186 10908
rect 20242 10906 20266 10908
rect 20322 10906 20346 10908
rect 20402 10906 20426 10908
rect 20482 10906 20488 10908
rect 20242 10854 20244 10906
rect 20424 10854 20426 10906
rect 20180 10852 20186 10854
rect 20242 10852 20266 10854
rect 20322 10852 20346 10854
rect 20402 10852 20426 10854
rect 20482 10852 20488 10854
rect 20180 10843 20488 10852
rect 20640 10690 20668 13126
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20824 12238 20852 12650
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11620 20772 11626
rect 20720 11562 20772 11568
rect 20456 10662 20668 10690
rect 20076 10192 20128 10198
rect 20168 10192 20220 10198
rect 20076 10134 20128 10140
rect 20166 10160 20168 10169
rect 20220 10160 20222 10169
rect 20166 10095 20222 10104
rect 20260 10056 20312 10062
rect 20088 10016 20260 10044
rect 20088 9042 20116 10016
rect 20260 9998 20312 10004
rect 20456 9994 20484 10662
rect 20732 10470 20760 11562
rect 20916 10810 20944 15370
rect 21284 14414 21312 15438
rect 21560 15162 21588 16934
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21744 16182 21772 16594
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22020 15162 22048 15438
rect 22112 15162 22140 17054
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22204 16590 22232 17002
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 22296 16182 22324 17138
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16590 22416 16934
rect 22664 16590 22692 18022
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22756 16794 22784 17138
rect 22848 16794 22876 18362
rect 23400 18290 23428 19450
rect 24780 19446 24808 19994
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24400 18828 24452 18834
rect 24400 18770 24452 18776
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23400 17202 23428 18226
rect 23860 18222 23888 18566
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23584 17202 23612 18158
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 23400 16998 23428 17138
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22480 16250 22508 16458
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21454 14376 21510 14385
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13258 21036 13670
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21100 12782 21128 14350
rect 21454 14311 21456 14320
rect 21508 14311 21510 14320
rect 21456 14282 21508 14288
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21284 12986 21312 13398
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21008 11830 21036 12378
rect 21192 12238 21220 12650
rect 21180 12232 21232 12238
rect 21272 12232 21324 12238
rect 21180 12174 21232 12180
rect 21270 12200 21272 12209
rect 21324 12200 21326 12209
rect 21270 12135 21326 12144
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20824 10538 20852 10610
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20180 9820 20488 9829
rect 20180 9818 20186 9820
rect 20242 9818 20266 9820
rect 20322 9818 20346 9820
rect 20402 9818 20426 9820
rect 20482 9818 20488 9820
rect 20242 9766 20244 9818
rect 20424 9766 20426 9818
rect 20180 9764 20186 9766
rect 20242 9764 20266 9766
rect 20322 9764 20346 9766
rect 20402 9764 20426 9766
rect 20482 9764 20488 9766
rect 20180 9755 20488 9764
rect 20260 9648 20312 9654
rect 20312 9608 20484 9636
rect 20260 9590 20312 9596
rect 20456 9466 20484 9608
rect 20548 9586 20576 9930
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20534 9480 20590 9489
rect 20456 9438 20534 9466
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20180 8906 20208 9318
rect 20456 8974 20484 9438
rect 20534 9415 20590 9424
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20444 8968 20496 8974
rect 20444 8910 20496 8916
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20180 8732 20488 8741
rect 20180 8730 20186 8732
rect 20242 8730 20266 8732
rect 20322 8730 20346 8732
rect 20402 8730 20426 8732
rect 20482 8730 20488 8732
rect 20242 8678 20244 8730
rect 20424 8678 20426 8730
rect 20180 8676 20186 8678
rect 20242 8676 20266 8678
rect 20322 8676 20346 8678
rect 20402 8676 20426 8678
rect 20482 8676 20488 8678
rect 20180 8667 20488 8676
rect 20548 8634 20576 9046
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 19904 8486 20024 8514
rect 19520 8188 19828 8197
rect 19520 8186 19526 8188
rect 19582 8186 19606 8188
rect 19662 8186 19686 8188
rect 19742 8186 19766 8188
rect 19822 8186 19828 8188
rect 19582 8134 19584 8186
rect 19764 8134 19766 8186
rect 19520 8132 19526 8134
rect 19582 8132 19606 8134
rect 19662 8132 19686 8134
rect 19742 8132 19766 8134
rect 19822 8132 19828 8134
rect 19520 8123 19828 8132
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19904 7886 19932 8486
rect 20640 8430 20668 10134
rect 20904 10056 20956 10062
rect 21008 10044 21036 11766
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21088 10600 21140 10606
rect 21284 10588 21312 11018
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21140 10560 21312 10588
rect 21088 10542 21140 10548
rect 20956 10016 21036 10044
rect 20904 9998 20956 10004
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 21008 9722 21036 9862
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20824 8634 20852 9114
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 7886 20024 8230
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 7478 19472 7686
rect 20180 7644 20488 7653
rect 20180 7642 20186 7644
rect 20242 7642 20266 7644
rect 20322 7642 20346 7644
rect 20402 7642 20426 7644
rect 20482 7642 20488 7644
rect 20242 7590 20244 7642
rect 20424 7590 20426 7642
rect 20180 7588 20186 7590
rect 20242 7588 20266 7590
rect 20322 7588 20346 7590
rect 20402 7588 20426 7590
rect 20482 7588 20488 7590
rect 20180 7579 20488 7588
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 19520 7100 19828 7109
rect 19520 7098 19526 7100
rect 19582 7098 19606 7100
rect 19662 7098 19686 7100
rect 19742 7098 19766 7100
rect 19822 7098 19828 7100
rect 19582 7046 19584 7098
rect 19764 7046 19766 7098
rect 19520 7044 19526 7046
rect 19582 7044 19606 7046
rect 19662 7044 19686 7046
rect 19742 7044 19766 7046
rect 19822 7044 19828 7046
rect 19520 7035 19828 7044
rect 20088 7002 20116 7414
rect 21008 7206 21036 7822
rect 21100 7342 21128 8366
rect 21192 8090 21220 8434
rect 21180 8084 21232 8090
rect 21284 8072 21312 10560
rect 21376 10470 21404 10678
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21468 10198 21496 14282
rect 21560 10266 21588 15098
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 21928 14618 21956 14758
rect 22112 14618 22140 14894
rect 22296 14822 22324 15438
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 21928 13394 21956 14554
rect 22572 14498 22600 16458
rect 22652 16176 22704 16182
rect 22756 16164 22784 16730
rect 22848 16590 22876 16730
rect 24136 16726 24164 17206
rect 24124 16720 24176 16726
rect 24124 16662 24176 16668
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22704 16136 22784 16164
rect 22652 16118 22704 16124
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22388 14470 22600 14498
rect 22388 14414 22416 14470
rect 22756 14414 22784 14758
rect 22940 14414 22968 16594
rect 23664 16584 23716 16590
rect 23662 16552 23664 16561
rect 23940 16584 23992 16590
rect 23716 16552 23718 16561
rect 23940 16526 23992 16532
rect 23662 16487 23718 16496
rect 23952 16250 23980 16526
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 24412 16182 24440 18770
rect 24492 18692 24544 18698
rect 24492 18634 24544 18640
rect 24504 18358 24532 18634
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24504 16250 24532 18294
rect 24780 17746 24808 19382
rect 24860 19304 24912 19310
rect 24860 19246 24912 19252
rect 24872 18970 24900 19246
rect 24964 19174 24992 20266
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24964 18834 24992 19110
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 25056 18290 25084 19722
rect 25228 18896 25280 18902
rect 25228 18838 25280 18844
rect 25240 18766 25268 18838
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 17338 25176 17546
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24676 16584 24728 16590
rect 24860 16584 24912 16590
rect 24728 16544 24808 16572
rect 24676 16526 24728 16532
rect 24780 16454 24808 16544
rect 24860 16526 24912 16532
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24400 16176 24452 16182
rect 24400 16118 24452 16124
rect 24688 15910 24716 16390
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 23768 15638 23796 15846
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24504 15094 24532 15370
rect 24780 15162 24808 16050
rect 24872 15706 24900 16526
rect 24964 15978 24992 17138
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16658 25084 16934
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 25056 15502 25084 16594
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25148 16182 25176 16526
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25240 16114 25268 16526
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25136 15904 25188 15910
rect 25332 15858 25360 20470
rect 25872 19440 25924 19446
rect 25872 19382 25924 19388
rect 25884 18426 25912 19382
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25976 18358 26004 23666
rect 26056 23588 26108 23594
rect 26056 23530 26108 23536
rect 26068 22642 26096 23530
rect 26948 23420 27256 23429
rect 26948 23418 26954 23420
rect 27010 23418 27034 23420
rect 27090 23418 27114 23420
rect 27170 23418 27194 23420
rect 27250 23418 27256 23420
rect 27010 23366 27012 23418
rect 27192 23366 27194 23418
rect 26948 23364 26954 23366
rect 27010 23364 27034 23366
rect 27090 23364 27114 23366
rect 27170 23364 27194 23366
rect 27250 23364 27256 23366
rect 26948 23355 27256 23364
rect 30300 23225 30328 23666
rect 30286 23216 30342 23225
rect 30286 23151 30342 23160
rect 27608 22876 27916 22885
rect 27608 22874 27614 22876
rect 27670 22874 27694 22876
rect 27750 22874 27774 22876
rect 27830 22874 27854 22876
rect 27910 22874 27916 22876
rect 27670 22822 27672 22874
rect 27852 22822 27854 22874
rect 27608 22820 27614 22822
rect 27670 22820 27694 22822
rect 27750 22820 27774 22822
rect 27830 22820 27854 22822
rect 27910 22820 27916 22822
rect 27608 22811 27916 22820
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 26252 21690 26280 22578
rect 30944 22545 30972 22578
rect 30930 22536 30986 22545
rect 30930 22471 30986 22480
rect 26948 22332 27256 22341
rect 26948 22330 26954 22332
rect 27010 22330 27034 22332
rect 27090 22330 27114 22332
rect 27170 22330 27194 22332
rect 27250 22330 27256 22332
rect 27010 22278 27012 22330
rect 27192 22278 27194 22330
rect 26948 22276 26954 22278
rect 27010 22276 27034 22278
rect 27090 22276 27114 22278
rect 27170 22276 27194 22278
rect 27250 22276 27256 22278
rect 26948 22267 27256 22276
rect 26608 21956 26660 21962
rect 26608 21898 26660 21904
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 26068 21010 26096 21354
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26160 20806 26188 21490
rect 26620 21486 26648 21898
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30470 21856 30526 21865
rect 27608 21788 27916 21797
rect 27608 21786 27614 21788
rect 27670 21786 27694 21788
rect 27750 21786 27774 21788
rect 27830 21786 27854 21788
rect 27910 21786 27916 21788
rect 27670 21734 27672 21786
rect 27852 21734 27854 21786
rect 27608 21732 27614 21734
rect 27670 21732 27694 21734
rect 27750 21732 27774 21734
rect 27830 21732 27854 21734
rect 27910 21732 27916 21734
rect 27608 21723 27916 21732
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 26160 20602 26188 20742
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26252 19514 26280 21286
rect 26344 20874 26372 21422
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 26344 20602 26372 20810
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26620 20534 26648 21422
rect 26948 21244 27256 21253
rect 26948 21242 26954 21244
rect 27010 21242 27034 21244
rect 27090 21242 27114 21244
rect 27170 21242 27194 21244
rect 27250 21242 27256 21244
rect 27010 21190 27012 21242
rect 27192 21190 27194 21242
rect 26948 21188 26954 21190
rect 27010 21188 27034 21190
rect 27090 21188 27114 21190
rect 27170 21188 27194 21190
rect 27250 21188 27256 21190
rect 26948 21179 27256 21188
rect 30392 21185 30420 21830
rect 30470 21791 30526 21800
rect 30484 21554 30512 21791
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 30378 21176 30434 21185
rect 30378 21111 30434 21120
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 27608 20700 27916 20709
rect 27608 20698 27614 20700
rect 27670 20698 27694 20700
rect 27750 20698 27774 20700
rect 27830 20698 27854 20700
rect 27910 20698 27916 20700
rect 27670 20646 27672 20698
rect 27852 20646 27854 20698
rect 27608 20644 27614 20646
rect 27670 20644 27694 20646
rect 27750 20644 27774 20646
rect 27830 20644 27854 20646
rect 27910 20644 27916 20646
rect 27608 20635 27916 20644
rect 26608 20528 26660 20534
rect 30300 20505 30328 20742
rect 26608 20470 26660 20476
rect 30286 20496 30342 20505
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26252 18834 26280 19450
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26620 18766 26648 20470
rect 30286 20431 30342 20440
rect 26948 20156 27256 20165
rect 26948 20154 26954 20156
rect 27010 20154 27034 20156
rect 27090 20154 27114 20156
rect 27170 20154 27194 20156
rect 27250 20154 27256 20156
rect 27010 20102 27012 20154
rect 27192 20102 27194 20154
rect 26948 20100 26954 20102
rect 27010 20100 27034 20102
rect 27090 20100 27114 20102
rect 27170 20100 27194 20102
rect 27250 20100 27256 20102
rect 26948 20091 27256 20100
rect 30380 19984 30432 19990
rect 30380 19926 30432 19932
rect 30392 19825 30420 19926
rect 30378 19816 30434 19825
rect 30378 19751 30434 19760
rect 27608 19612 27916 19621
rect 27608 19610 27614 19612
rect 27670 19610 27694 19612
rect 27750 19610 27774 19612
rect 27830 19610 27854 19612
rect 27910 19610 27916 19612
rect 27670 19558 27672 19610
rect 27852 19558 27854 19610
rect 27608 19556 27614 19558
rect 27670 19556 27694 19558
rect 27750 19556 27774 19558
rect 27830 19556 27854 19558
rect 27910 19556 27916 19558
rect 27608 19547 27916 19556
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30300 19145 30328 19314
rect 30286 19136 30342 19145
rect 26948 19068 27256 19077
rect 30286 19071 30342 19080
rect 26948 19066 26954 19068
rect 27010 19066 27034 19068
rect 27090 19066 27114 19068
rect 27170 19066 27194 19068
rect 27250 19066 27256 19068
rect 27010 19014 27012 19066
rect 27192 19014 27194 19066
rect 26948 19012 26954 19014
rect 27010 19012 27034 19014
rect 27090 19012 27114 19014
rect 27170 19012 27194 19014
rect 27250 19012 27256 19014
rect 26948 19003 27256 19012
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25516 16658 25544 16934
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25504 16652 25556 16658
rect 25504 16594 25556 16600
rect 25608 16250 25636 16730
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 25596 16244 25648 16250
rect 25596 16186 25648 16192
rect 25700 16114 25728 16662
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25792 16250 25820 16526
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25136 15846 25188 15852
rect 25148 15706 25176 15846
rect 25240 15830 25360 15858
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25148 15502 25176 15642
rect 25044 15496 25096 15502
rect 25044 15438 25096 15444
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24492 15088 24544 15094
rect 24492 15030 24544 15036
rect 24504 14618 24532 15030
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21836 12986 21864 13126
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21928 12434 21956 13330
rect 21836 12406 21956 12434
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21652 11354 21680 11698
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21836 11218 21864 12406
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21744 10470 21772 10610
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21652 10062 21680 10406
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21836 9450 21864 11154
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21928 10538 21956 11018
rect 22020 10810 22048 11494
rect 22112 11234 22140 13874
rect 22296 13734 22324 14282
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22388 13546 22416 14350
rect 22664 14074 22692 14350
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22296 13518 22416 13546
rect 22296 13258 22324 13518
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22192 12912 22244 12918
rect 22192 12854 22244 12860
rect 22204 11558 22232 12854
rect 22296 12646 22324 13194
rect 22388 12646 22416 13330
rect 22480 12850 22508 13670
rect 22664 13394 22692 14010
rect 22756 14006 22784 14350
rect 22940 14006 22968 14350
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24412 14074 24440 14214
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 22744 14000 22796 14006
rect 22744 13942 22796 13948
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22756 13326 22784 13942
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22572 12918 22600 13126
rect 22664 12986 22692 13126
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22940 12782 22968 13942
rect 24780 13938 24808 14758
rect 24872 14414 24900 14758
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 23388 13388 23440 13394
rect 23388 13330 23440 13336
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 12986 23060 13262
rect 23400 12986 23428 13330
rect 24504 13326 24532 13806
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24504 12986 24532 13126
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24688 12782 24716 13262
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24872 12850 24900 13126
rect 24964 12986 24992 15302
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25056 14618 25084 15098
rect 25240 14822 25268 15830
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25228 14816 25280 14822
rect 25228 14758 25280 14764
rect 25332 14618 25360 15642
rect 25700 15570 25728 16050
rect 25780 15904 25832 15910
rect 25780 15846 25832 15852
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25792 15570 25820 15846
rect 25884 15706 25912 15846
rect 25872 15700 25924 15706
rect 25872 15642 25924 15648
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25976 15502 26004 16934
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 25516 14618 25544 15438
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 25320 14612 25372 14618
rect 25320 14554 25372 14560
rect 25504 14612 25556 14618
rect 25504 14554 25556 14560
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25056 12866 25084 14554
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25148 13394 25176 13942
rect 25240 13734 25268 14418
rect 25332 14074 25360 14554
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25884 13326 25912 14282
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24964 12838 25084 12866
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 22284 12640 22336 12646
rect 22284 12582 22336 12588
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22572 11694 22600 12718
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 22928 12232 22980 12238
rect 22928 12174 22980 12180
rect 22940 11898 22968 12174
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22112 11206 22232 11234
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21928 9518 21956 10474
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21468 8090 21496 9318
rect 21640 9036 21692 9042
rect 21640 8978 21692 8984
rect 21652 8634 21680 8978
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21836 8430 21864 9386
rect 21928 9178 21956 9454
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22112 8566 22140 9862
rect 22100 8560 22152 8566
rect 22100 8502 22152 8508
rect 22204 8514 22232 11206
rect 22664 10674 22692 11834
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22940 11354 22968 11630
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22940 10810 22968 11290
rect 23032 11014 23060 12582
rect 24872 12374 24900 12786
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24964 12170 24992 12838
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 25056 12442 25084 12582
rect 25044 12436 25096 12442
rect 25044 12378 25096 12384
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 24952 12164 25004 12170
rect 24952 12106 25004 12112
rect 24044 11898 24072 12106
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23124 11354 23152 11494
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23020 11008 23072 11014
rect 23124 10996 23152 11086
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 23072 10968 23152 10996
rect 23020 10950 23072 10956
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 23032 10674 23060 10950
rect 23676 10742 23704 11018
rect 23664 10736 23716 10742
rect 23664 10678 23716 10684
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22572 10062 22600 10610
rect 23032 10470 23060 10610
rect 23768 10538 23796 11562
rect 23952 11354 23980 11698
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 23952 11150 23980 11290
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 24044 10606 24072 11630
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 23204 10260 23256 10266
rect 23204 10202 23256 10208
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22388 9722 22416 9998
rect 23216 9994 23244 10202
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22296 9466 22324 9658
rect 23388 9512 23440 9518
rect 22296 9438 22416 9466
rect 23388 9454 23440 9460
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9178 22324 9318
rect 22388 9178 22416 9438
rect 23400 9178 23428 9454
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23492 8974 23520 10474
rect 23584 10266 23612 10474
rect 23768 10266 23796 10474
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23952 10266 23980 10406
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23756 10260 23808 10266
rect 23756 10202 23808 10208
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 24136 10062 24164 10678
rect 24412 10538 24440 11698
rect 24504 11150 24532 11698
rect 24780 11354 24808 11698
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24780 11150 24808 11290
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24400 10532 24452 10538
rect 24400 10474 24452 10480
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23584 9110 23612 9318
rect 23768 9178 23796 9930
rect 24492 9920 24544 9926
rect 24492 9862 24544 9868
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23112 8560 23164 8566
rect 22204 8486 22324 8514
rect 23112 8502 23164 8508
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22204 8090 22232 8366
rect 21364 8084 21416 8090
rect 21284 8044 21364 8072
rect 21180 8026 21232 8032
rect 21364 8026 21416 8032
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 21376 7750 21404 8026
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21928 7750 21956 7958
rect 22296 7750 22324 8486
rect 23124 8090 23152 8502
rect 23584 8430 23612 9046
rect 24412 8634 24440 9590
rect 24504 9178 24532 9862
rect 24492 9172 24544 9178
rect 24492 9114 24544 9120
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24872 8498 24900 10610
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24964 9518 24992 10134
rect 25056 10062 25084 12378
rect 25332 12238 25360 12922
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25700 12170 25728 12786
rect 25884 12782 25912 13262
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25320 12096 25372 12102
rect 25320 12038 25372 12044
rect 25332 11898 25360 12038
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25240 11286 25268 11698
rect 25700 11694 25728 12106
rect 26160 11694 26188 17002
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26344 16250 26372 16730
rect 26436 16658 26464 18566
rect 27608 18524 27916 18533
rect 27608 18522 27614 18524
rect 27670 18522 27694 18524
rect 27750 18522 27774 18524
rect 27830 18522 27854 18524
rect 27910 18522 27916 18524
rect 27670 18470 27672 18522
rect 27852 18470 27854 18522
rect 27608 18468 27614 18470
rect 27670 18468 27694 18470
rect 27750 18468 27774 18470
rect 27830 18468 27854 18470
rect 27910 18468 27916 18470
rect 27608 18459 27916 18468
rect 30392 18465 30420 18566
rect 30378 18456 30434 18465
rect 30378 18391 30434 18400
rect 27436 18352 27488 18358
rect 27436 18294 27488 18300
rect 26948 17980 27256 17989
rect 26948 17978 26954 17980
rect 27010 17978 27034 17980
rect 27090 17978 27114 17980
rect 27170 17978 27194 17980
rect 27250 17978 27256 17980
rect 27010 17926 27012 17978
rect 27192 17926 27194 17978
rect 26948 17924 26954 17926
rect 27010 17924 27034 17926
rect 27090 17924 27114 17926
rect 27170 17924 27194 17926
rect 27250 17924 27256 17926
rect 26948 17915 27256 17924
rect 27448 17678 27476 18294
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30300 17785 30328 18022
rect 30286 17776 30342 17785
rect 30286 17711 30342 17720
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 26700 17536 26752 17542
rect 26700 17478 26752 17484
rect 26712 17338 26740 17478
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 27356 17202 27384 17614
rect 27608 17436 27916 17445
rect 27608 17434 27614 17436
rect 27670 17434 27694 17436
rect 27750 17434 27774 17436
rect 27830 17434 27854 17436
rect 27910 17434 27916 17436
rect 27670 17382 27672 17434
rect 27852 17382 27854 17434
rect 27608 17380 27614 17382
rect 27670 17380 27694 17382
rect 27750 17380 27774 17382
rect 27830 17380 27854 17382
rect 27910 17380 27916 17382
rect 27608 17371 27916 17380
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 26948 16892 27256 16901
rect 26948 16890 26954 16892
rect 27010 16890 27034 16892
rect 27090 16890 27114 16892
rect 27170 16890 27194 16892
rect 27250 16890 27256 16892
rect 27010 16838 27012 16890
rect 27192 16838 27194 16890
rect 26948 16836 26954 16838
rect 27010 16836 27034 16838
rect 27090 16836 27114 16838
rect 27170 16836 27194 16838
rect 27250 16836 27256 16838
rect 26948 16827 27256 16836
rect 27356 16658 27384 17138
rect 30378 17096 30434 17105
rect 30378 17031 30380 17040
rect 30432 17031 30434 17040
rect 30380 17002 30432 17008
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26436 15910 26464 16594
rect 30932 16516 30984 16522
rect 30932 16458 30984 16464
rect 30944 16425 30972 16458
rect 30930 16416 30986 16425
rect 27608 16348 27916 16357
rect 30930 16351 30986 16360
rect 27608 16346 27614 16348
rect 27670 16346 27694 16348
rect 27750 16346 27774 16348
rect 27830 16346 27854 16348
rect 27910 16346 27916 16348
rect 27670 16294 27672 16346
rect 27852 16294 27854 16346
rect 27608 16292 27614 16294
rect 27670 16292 27694 16294
rect 27750 16292 27774 16294
rect 27830 16292 27854 16294
rect 27910 16292 27916 16294
rect 27608 16283 27916 16292
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 26948 15804 27256 15813
rect 26948 15802 26954 15804
rect 27010 15802 27034 15804
rect 27090 15802 27114 15804
rect 27170 15802 27194 15804
rect 27250 15802 27256 15804
rect 27010 15750 27012 15802
rect 27192 15750 27194 15802
rect 26948 15748 26954 15750
rect 27010 15748 27034 15750
rect 27090 15748 27114 15750
rect 27170 15748 27194 15750
rect 27250 15748 27256 15750
rect 26948 15739 27256 15748
rect 30392 15745 30420 15846
rect 30378 15736 30434 15745
rect 30378 15671 30434 15680
rect 30288 15360 30340 15366
rect 30288 15302 30340 15308
rect 27608 15260 27916 15269
rect 27608 15258 27614 15260
rect 27670 15258 27694 15260
rect 27750 15258 27774 15260
rect 27830 15258 27854 15260
rect 27910 15258 27916 15260
rect 27670 15206 27672 15258
rect 27852 15206 27854 15258
rect 27608 15204 27614 15206
rect 27670 15204 27694 15206
rect 27750 15204 27774 15206
rect 27830 15204 27854 15206
rect 27910 15204 27916 15206
rect 27608 15195 27916 15204
rect 30300 15065 30328 15302
rect 30286 15056 30342 15065
rect 30286 14991 30342 15000
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 26948 14716 27256 14725
rect 26948 14714 26954 14716
rect 27010 14714 27034 14716
rect 27090 14714 27114 14716
rect 27170 14714 27194 14716
rect 27250 14714 27256 14716
rect 27010 14662 27012 14714
rect 27192 14662 27194 14714
rect 26948 14660 26954 14662
rect 27010 14660 27034 14662
rect 27090 14660 27114 14662
rect 27170 14660 27194 14662
rect 27250 14660 27256 14662
rect 26948 14651 27256 14660
rect 30208 14414 30236 14758
rect 30380 14544 30432 14550
rect 30380 14486 30432 14492
rect 30196 14408 30248 14414
rect 30392 14385 30420 14486
rect 30196 14350 30248 14356
rect 30378 14376 30434 14385
rect 30378 14311 30434 14320
rect 27608 14172 27916 14181
rect 27608 14170 27614 14172
rect 27670 14170 27694 14172
rect 27750 14170 27774 14172
rect 27830 14170 27854 14172
rect 27910 14170 27916 14172
rect 27670 14118 27672 14170
rect 27852 14118 27854 14170
rect 27608 14116 27614 14118
rect 27670 14116 27694 14118
rect 27750 14116 27774 14118
rect 27830 14116 27854 14118
rect 27910 14116 27916 14118
rect 27608 14107 27916 14116
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 30288 13864 30340 13870
rect 30288 13806 30340 13812
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 26948 13628 27256 13637
rect 26948 13626 26954 13628
rect 27010 13626 27034 13628
rect 27090 13626 27114 13628
rect 27170 13626 27194 13628
rect 27250 13626 27256 13628
rect 27010 13574 27012 13626
rect 27192 13574 27194 13626
rect 26948 13572 26954 13574
rect 27010 13572 27034 13574
rect 27090 13572 27114 13574
rect 27170 13572 27194 13574
rect 27250 13572 27256 13574
rect 26948 13563 27256 13572
rect 29012 13462 29040 13670
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 27608 13084 27916 13093
rect 27608 13082 27614 13084
rect 27670 13082 27694 13084
rect 27750 13082 27774 13084
rect 27830 13082 27854 13084
rect 27910 13082 27916 13084
rect 27670 13030 27672 13082
rect 27852 13030 27854 13082
rect 27608 13028 27614 13030
rect 27670 13028 27694 13030
rect 27750 13028 27774 13030
rect 27830 13028 27854 13030
rect 27910 13028 27916 13030
rect 27608 13019 27916 13028
rect 30208 12986 30236 13806
rect 30300 13705 30328 13806
rect 30286 13696 30342 13705
rect 30286 13631 30342 13640
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30392 13025 30420 13126
rect 30378 13016 30434 13025
rect 30196 12980 30248 12986
rect 30378 12951 30434 12960
rect 30196 12922 30248 12928
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 26948 12540 27256 12549
rect 26948 12538 26954 12540
rect 27010 12538 27034 12540
rect 27090 12538 27114 12540
rect 27170 12538 27194 12540
rect 27250 12538 27256 12540
rect 27010 12486 27012 12538
rect 27192 12486 27194 12538
rect 26948 12484 26954 12486
rect 27010 12484 27034 12486
rect 27090 12484 27114 12486
rect 27170 12484 27194 12486
rect 27250 12484 27256 12486
rect 26948 12475 27256 12484
rect 30300 12345 30328 12786
rect 30286 12336 30342 12345
rect 30286 12271 30342 12280
rect 27608 11996 27916 12005
rect 27608 11994 27614 11996
rect 27670 11994 27694 11996
rect 27750 11994 27774 11996
rect 27830 11994 27854 11996
rect 27910 11994 27916 11996
rect 27670 11942 27672 11994
rect 27852 11942 27854 11994
rect 27608 11940 27614 11942
rect 27670 11940 27694 11942
rect 27750 11940 27774 11942
rect 27830 11940 27854 11942
rect 27910 11940 27916 11942
rect 27608 11931 27916 11940
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25228 11280 25280 11286
rect 25228 11222 25280 11228
rect 25412 11280 25464 11286
rect 25412 11222 25464 11228
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 25148 10062 25176 10406
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 24952 9512 25004 9518
rect 25332 9489 25360 10066
rect 25424 10062 25452 11222
rect 25700 11218 25728 11494
rect 26948 11452 27256 11461
rect 26948 11450 26954 11452
rect 27010 11450 27034 11452
rect 27090 11450 27114 11452
rect 27170 11450 27194 11452
rect 27250 11450 27256 11452
rect 27010 11398 27012 11450
rect 27192 11398 27194 11450
rect 26948 11396 26954 11398
rect 27010 11396 27034 11398
rect 27090 11396 27114 11398
rect 27170 11396 27194 11398
rect 27250 11396 27256 11398
rect 26948 11387 27256 11396
rect 27632 11354 27660 11698
rect 30378 11656 30434 11665
rect 30378 11591 30380 11600
rect 30432 11591 30434 11600
rect 30380 11562 30432 11568
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 10810 26280 11018
rect 30300 10985 30328 11086
rect 30286 10976 30342 10985
rect 27608 10908 27916 10917
rect 30286 10911 30342 10920
rect 27608 10906 27614 10908
rect 27670 10906 27694 10908
rect 27750 10906 27774 10908
rect 27830 10906 27854 10908
rect 27910 10906 27916 10908
rect 27670 10854 27672 10906
rect 27852 10854 27854 10906
rect 27608 10852 27614 10854
rect 27670 10852 27694 10854
rect 27750 10852 27774 10854
rect 27830 10852 27854 10854
rect 27910 10852 27916 10854
rect 27608 10843 27916 10852
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 26948 10364 27256 10373
rect 26948 10362 26954 10364
rect 27010 10362 27034 10364
rect 27090 10362 27114 10364
rect 27170 10362 27194 10364
rect 27250 10362 27256 10364
rect 27010 10310 27012 10362
rect 27192 10310 27194 10362
rect 26948 10308 26954 10310
rect 27010 10308 27034 10310
rect 27090 10308 27114 10310
rect 27170 10308 27194 10310
rect 27250 10308 27256 10310
rect 26948 10299 27256 10308
rect 30944 10305 30972 10610
rect 30930 10296 30986 10305
rect 30930 10231 30986 10240
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 30288 10056 30340 10062
rect 30288 9998 30340 10004
rect 27608 9820 27916 9829
rect 27608 9818 27614 9820
rect 27670 9818 27694 9820
rect 27750 9818 27774 9820
rect 27830 9818 27854 9820
rect 27910 9818 27916 9820
rect 27670 9766 27672 9818
rect 27852 9766 27854 9818
rect 27608 9764 27614 9766
rect 27670 9764 27694 9766
rect 27750 9764 27774 9766
rect 27830 9764 27854 9766
rect 27910 9764 27916 9766
rect 27608 9755 27916 9764
rect 30300 9625 30328 9998
rect 30286 9616 30342 9625
rect 30286 9551 30342 9560
rect 25596 9512 25648 9518
rect 24952 9454 25004 9460
rect 25318 9480 25374 9489
rect 25596 9454 25648 9460
rect 25318 9415 25374 9424
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 9178 24992 9318
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 25608 8974 25636 9454
rect 26948 9276 27256 9285
rect 26948 9274 26954 9276
rect 27010 9274 27034 9276
rect 27090 9274 27114 9276
rect 27170 9274 27194 9276
rect 27250 9274 27256 9276
rect 27010 9222 27012 9274
rect 27192 9222 27194 9274
rect 26948 9220 26954 9222
rect 27010 9220 27034 9222
rect 27090 9220 27114 9222
rect 27170 9220 27194 9222
rect 27250 9220 27256 9222
rect 26948 9211 27256 9220
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 25596 8968 25648 8974
rect 30392 8945 30420 9114
rect 25596 8910 25648 8916
rect 30378 8936 30434 8945
rect 30378 8871 30434 8880
rect 27608 8732 27916 8741
rect 27608 8730 27614 8732
rect 27670 8730 27694 8732
rect 27750 8730 27774 8732
rect 27830 8730 27854 8732
rect 27910 8730 27916 8732
rect 27670 8678 27672 8730
rect 27852 8678 27854 8730
rect 27608 8676 27614 8678
rect 27670 8676 27694 8678
rect 27750 8676 27774 8678
rect 27830 8676 27854 8678
rect 27910 8676 27916 8678
rect 27608 8667 27916 8676
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23112 8084 23164 8090
rect 23112 8026 23164 8032
rect 23676 7886 23704 8434
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 30300 8265 30328 8298
rect 30286 8256 30342 8265
rect 26948 8188 27256 8197
rect 30286 8191 30342 8200
rect 26948 8186 26954 8188
rect 27010 8186 27034 8188
rect 27090 8186 27114 8188
rect 27170 8186 27194 8188
rect 27250 8186 27256 8188
rect 27010 8134 27012 8186
rect 27192 8134 27194 8186
rect 26948 8132 26954 8134
rect 27010 8132 27034 8134
rect 27090 8132 27114 8134
rect 27170 8132 27194 8134
rect 27250 8132 27256 8134
rect 26948 8123 27256 8132
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20180 6556 20488 6565
rect 20180 6554 20186 6556
rect 20242 6554 20266 6556
rect 20322 6554 20346 6556
rect 20402 6554 20426 6556
rect 20482 6554 20488 6556
rect 20242 6502 20244 6554
rect 20424 6502 20426 6554
rect 20180 6500 20186 6502
rect 20242 6500 20266 6502
rect 20322 6500 20346 6502
rect 20402 6500 20426 6502
rect 20482 6500 20488 6502
rect 20180 6491 20488 6500
rect 19520 6012 19828 6021
rect 19520 6010 19526 6012
rect 19582 6010 19606 6012
rect 19662 6010 19686 6012
rect 19742 6010 19766 6012
rect 19822 6010 19828 6012
rect 19582 5958 19584 6010
rect 19764 5958 19766 6010
rect 19520 5956 19526 5958
rect 19582 5956 19606 5958
rect 19662 5956 19686 5958
rect 19742 5956 19766 5958
rect 19822 5956 19828 5958
rect 19520 5947 19828 5956
rect 20180 5468 20488 5477
rect 20180 5466 20186 5468
rect 20242 5466 20266 5468
rect 20322 5466 20346 5468
rect 20402 5466 20426 5468
rect 20482 5466 20488 5468
rect 20242 5414 20244 5466
rect 20424 5414 20426 5466
rect 20180 5412 20186 5414
rect 20242 5412 20266 5414
rect 20322 5412 20346 5414
rect 20402 5412 20426 5414
rect 20482 5412 20488 5414
rect 20180 5403 20488 5412
rect 19520 4924 19828 4933
rect 19520 4922 19526 4924
rect 19582 4922 19606 4924
rect 19662 4922 19686 4924
rect 19742 4922 19766 4924
rect 19822 4922 19828 4924
rect 19582 4870 19584 4922
rect 19764 4870 19766 4922
rect 19520 4868 19526 4870
rect 19582 4868 19606 4870
rect 19662 4868 19686 4870
rect 19742 4868 19766 4870
rect 19822 4868 19828 4870
rect 19520 4859 19828 4868
rect 20180 4380 20488 4389
rect 20180 4378 20186 4380
rect 20242 4378 20266 4380
rect 20322 4378 20346 4380
rect 20402 4378 20426 4380
rect 20482 4378 20488 4380
rect 20242 4326 20244 4378
rect 20424 4326 20426 4378
rect 20180 4324 20186 4326
rect 20242 4324 20266 4326
rect 20322 4324 20346 4326
rect 20402 4324 20426 4326
rect 20482 4324 20488 4326
rect 20180 4315 20488 4324
rect 19520 3836 19828 3845
rect 19520 3834 19526 3836
rect 19582 3834 19606 3836
rect 19662 3834 19686 3836
rect 19742 3834 19766 3836
rect 19822 3834 19828 3836
rect 19582 3782 19584 3834
rect 19764 3782 19766 3834
rect 19520 3780 19526 3782
rect 19582 3780 19606 3782
rect 19662 3780 19686 3782
rect 19742 3780 19766 3782
rect 19822 3780 19828 3782
rect 19520 3771 19828 3780
rect 20180 3292 20488 3301
rect 20180 3290 20186 3292
rect 20242 3290 20266 3292
rect 20322 3290 20346 3292
rect 20402 3290 20426 3292
rect 20482 3290 20488 3292
rect 20242 3238 20244 3290
rect 20424 3238 20426 3290
rect 20180 3236 20186 3238
rect 20242 3236 20266 3238
rect 20322 3236 20346 3238
rect 20402 3236 20426 3238
rect 20482 3236 20488 3238
rect 20180 3227 20488 3236
rect 18892 2746 19012 2774
rect 18984 2650 19012 2746
rect 19520 2748 19828 2757
rect 19520 2746 19526 2748
rect 19582 2746 19606 2748
rect 19662 2746 19686 2748
rect 19742 2746 19766 2748
rect 19822 2746 19828 2748
rect 19582 2694 19584 2746
rect 19764 2694 19766 2746
rect 19520 2692 19526 2694
rect 19582 2692 19606 2694
rect 19662 2692 19686 2694
rect 19742 2692 19766 2694
rect 19822 2692 19828 2694
rect 19520 2683 19828 2692
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 21008 2446 21036 7142
rect 21376 2774 21404 7686
rect 22296 6798 22324 7686
rect 27608 7644 27916 7653
rect 27608 7642 27614 7644
rect 27670 7642 27694 7644
rect 27750 7642 27774 7644
rect 27830 7642 27854 7644
rect 27910 7642 27916 7644
rect 27670 7590 27672 7642
rect 27852 7590 27854 7642
rect 27608 7588 27614 7590
rect 27670 7588 27694 7590
rect 27750 7588 27774 7590
rect 27830 7588 27854 7590
rect 27910 7588 27916 7590
rect 27608 7579 27916 7588
rect 26948 7100 27256 7109
rect 26948 7098 26954 7100
rect 27010 7098 27034 7100
rect 27090 7098 27114 7100
rect 27170 7098 27194 7100
rect 27250 7098 27256 7100
rect 27010 7046 27012 7098
rect 27192 7046 27194 7098
rect 26948 7044 26954 7046
rect 27010 7044 27034 7046
rect 27090 7044 27114 7046
rect 27170 7044 27194 7046
rect 27250 7044 27256 7046
rect 26948 7035 27256 7044
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 27608 6556 27916 6565
rect 27608 6554 27614 6556
rect 27670 6554 27694 6556
rect 27750 6554 27774 6556
rect 27830 6554 27854 6556
rect 27910 6554 27916 6556
rect 27670 6502 27672 6554
rect 27852 6502 27854 6554
rect 27608 6500 27614 6502
rect 27670 6500 27694 6502
rect 27750 6500 27774 6502
rect 27830 6500 27854 6502
rect 27910 6500 27916 6502
rect 27608 6491 27916 6500
rect 26948 6012 27256 6021
rect 26948 6010 26954 6012
rect 27010 6010 27034 6012
rect 27090 6010 27114 6012
rect 27170 6010 27194 6012
rect 27250 6010 27256 6012
rect 27010 5958 27012 6010
rect 27192 5958 27194 6010
rect 26948 5956 26954 5958
rect 27010 5956 27034 5958
rect 27090 5956 27114 5958
rect 27170 5956 27194 5958
rect 27250 5956 27256 5958
rect 26948 5947 27256 5956
rect 27608 5468 27916 5477
rect 27608 5466 27614 5468
rect 27670 5466 27694 5468
rect 27750 5466 27774 5468
rect 27830 5466 27854 5468
rect 27910 5466 27916 5468
rect 27670 5414 27672 5466
rect 27852 5414 27854 5466
rect 27608 5412 27614 5414
rect 27670 5412 27694 5414
rect 27750 5412 27774 5414
rect 27830 5412 27854 5414
rect 27910 5412 27916 5414
rect 27608 5403 27916 5412
rect 26948 4924 27256 4933
rect 26948 4922 26954 4924
rect 27010 4922 27034 4924
rect 27090 4922 27114 4924
rect 27170 4922 27194 4924
rect 27250 4922 27256 4924
rect 27010 4870 27012 4922
rect 27192 4870 27194 4922
rect 26948 4868 26954 4870
rect 27010 4868 27034 4870
rect 27090 4868 27114 4870
rect 27170 4868 27194 4870
rect 27250 4868 27256 4870
rect 26948 4859 27256 4868
rect 27608 4380 27916 4389
rect 27608 4378 27614 4380
rect 27670 4378 27694 4380
rect 27750 4378 27774 4380
rect 27830 4378 27854 4380
rect 27910 4378 27916 4380
rect 27670 4326 27672 4378
rect 27852 4326 27854 4378
rect 27608 4324 27614 4326
rect 27670 4324 27694 4326
rect 27750 4324 27774 4326
rect 27830 4324 27854 4326
rect 27910 4324 27916 4326
rect 27608 4315 27916 4324
rect 26948 3836 27256 3845
rect 26948 3834 26954 3836
rect 27010 3834 27034 3836
rect 27090 3834 27114 3836
rect 27170 3834 27194 3836
rect 27250 3834 27256 3836
rect 27010 3782 27012 3834
rect 27192 3782 27194 3834
rect 26948 3780 26954 3782
rect 27010 3780 27034 3782
rect 27090 3780 27114 3782
rect 27170 3780 27194 3782
rect 27250 3780 27256 3782
rect 26948 3771 27256 3780
rect 27608 3292 27916 3301
rect 27608 3290 27614 3292
rect 27670 3290 27694 3292
rect 27750 3290 27774 3292
rect 27830 3290 27854 3292
rect 27910 3290 27916 3292
rect 27670 3238 27672 3290
rect 27852 3238 27854 3290
rect 27608 3236 27614 3238
rect 27670 3236 27694 3238
rect 27750 3236 27774 3238
rect 27830 3236 27854 3238
rect 27910 3236 27916 3238
rect 27608 3227 27916 3236
rect 21376 2746 21496 2774
rect 21468 2650 21496 2746
rect 26948 2748 27256 2757
rect 26948 2746 26954 2748
rect 27010 2746 27034 2748
rect 27090 2746 27114 2748
rect 27170 2746 27194 2748
rect 27250 2746 27256 2748
rect 27010 2694 27012 2746
rect 27192 2694 27194 2746
rect 26948 2692 26954 2694
rect 27010 2692 27034 2694
rect 27090 2692 27114 2694
rect 27170 2692 27194 2694
rect 27250 2692 27256 2694
rect 26948 2683 27256 2692
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 18420 2440 18472 2446
rect 18788 2440 18840 2446
rect 18420 2382 18472 2388
rect 18708 2400 18788 2428
rect 5324 2204 5632 2213
rect 5324 2202 5330 2204
rect 5386 2202 5410 2204
rect 5466 2202 5490 2204
rect 5546 2202 5570 2204
rect 5626 2202 5632 2204
rect 5386 2150 5388 2202
rect 5568 2150 5570 2202
rect 5324 2148 5330 2150
rect 5386 2148 5410 2150
rect 5466 2148 5490 2150
rect 5546 2148 5570 2150
rect 5626 2148 5632 2150
rect 5324 2139 5632 2148
rect 9140 1306 9168 2382
rect 9784 1306 9812 2382
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9048 1278 9168 1306
rect 9692 1278 9812 1306
rect 9048 800 9076 1278
rect 9692 800 9720 1278
rect 10336 800 10364 2246
rect 11716 1306 11744 2382
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 11624 1278 11744 1306
rect 11624 800 11652 1278
rect 12268 800 12296 2246
rect 12752 2204 13060 2213
rect 12752 2202 12758 2204
rect 12814 2202 12838 2204
rect 12894 2202 12918 2204
rect 12974 2202 12998 2204
rect 13054 2202 13060 2204
rect 12814 2150 12816 2202
rect 12996 2150 12998 2202
rect 12752 2148 12758 2150
rect 12814 2148 12838 2150
rect 12894 2148 12918 2150
rect 12974 2148 12998 2150
rect 13054 2148 13060 2150
rect 12752 2139 13060 2148
rect 13096 1170 13124 2246
rect 13648 1306 13676 2382
rect 15016 2372 15068 2378
rect 12912 1142 13124 1170
rect 13556 1278 13676 1306
rect 14844 2332 15016 2360
rect 12912 800 12940 1142
rect 13556 800 13584 1278
rect 14844 800 14872 2332
rect 15016 2314 15068 2320
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 15672 1170 15700 2246
rect 16316 1170 16344 2246
rect 16960 1170 16988 2314
rect 17604 1170 17632 2314
rect 18236 2304 18288 2310
rect 15488 1142 15700 1170
rect 16132 1142 16344 1170
rect 16776 1142 16988 1170
rect 17420 1142 17632 1170
rect 18064 2264 18236 2292
rect 15488 800 15516 1142
rect 16132 800 16160 1142
rect 16776 800 16804 1142
rect 17420 800 17448 1142
rect 18064 800 18092 2264
rect 18236 2246 18288 2252
rect 18708 800 18736 2400
rect 18788 2382 18840 2388
rect 20996 2440 21048 2446
rect 21364 2440 21416 2446
rect 20996 2382 21048 2388
rect 21284 2400 21364 2428
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20180 2204 20488 2213
rect 20180 2202 20186 2204
rect 20242 2202 20266 2204
rect 20322 2202 20346 2204
rect 20402 2202 20426 2204
rect 20482 2202 20488 2204
rect 20242 2150 20244 2202
rect 20424 2150 20426 2202
rect 20180 2148 20186 2150
rect 20242 2148 20266 2150
rect 20322 2148 20346 2150
rect 20402 2148 20426 2150
rect 20482 2148 20488 2150
rect 20180 2139 20488 2148
rect 20640 800 20668 2246
rect 21284 800 21312 2400
rect 21364 2382 21416 2388
rect 27608 2204 27916 2213
rect 27608 2202 27614 2204
rect 27670 2202 27694 2204
rect 27750 2202 27774 2204
rect 27830 2202 27854 2204
rect 27910 2202 27916 2204
rect 27670 2150 27672 2202
rect 27852 2150 27854 2202
rect 27608 2148 27614 2150
rect 27670 2148 27694 2150
rect 27750 2148 27774 2150
rect 27830 2148 27854 2150
rect 27910 2148 27916 2150
rect 27608 2139 27916 2148
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 21270 0 21326 800
<< via2 >>
rect 5330 29402 5386 29404
rect 5410 29402 5466 29404
rect 5490 29402 5546 29404
rect 5570 29402 5626 29404
rect 5330 29350 5376 29402
rect 5376 29350 5386 29402
rect 5410 29350 5440 29402
rect 5440 29350 5452 29402
rect 5452 29350 5466 29402
rect 5490 29350 5504 29402
rect 5504 29350 5516 29402
rect 5516 29350 5546 29402
rect 5570 29350 5580 29402
rect 5580 29350 5626 29402
rect 5330 29348 5386 29350
rect 5410 29348 5466 29350
rect 5490 29348 5546 29350
rect 5570 29348 5626 29350
rect 12758 29402 12814 29404
rect 12838 29402 12894 29404
rect 12918 29402 12974 29404
rect 12998 29402 13054 29404
rect 12758 29350 12804 29402
rect 12804 29350 12814 29402
rect 12838 29350 12868 29402
rect 12868 29350 12880 29402
rect 12880 29350 12894 29402
rect 12918 29350 12932 29402
rect 12932 29350 12944 29402
rect 12944 29350 12974 29402
rect 12998 29350 13008 29402
rect 13008 29350 13054 29402
rect 12758 29348 12814 29350
rect 12838 29348 12894 29350
rect 12918 29348 12974 29350
rect 12998 29348 13054 29350
rect 20186 29402 20242 29404
rect 20266 29402 20322 29404
rect 20346 29402 20402 29404
rect 20426 29402 20482 29404
rect 20186 29350 20232 29402
rect 20232 29350 20242 29402
rect 20266 29350 20296 29402
rect 20296 29350 20308 29402
rect 20308 29350 20322 29402
rect 20346 29350 20360 29402
rect 20360 29350 20372 29402
rect 20372 29350 20402 29402
rect 20426 29350 20436 29402
rect 20436 29350 20482 29402
rect 20186 29348 20242 29350
rect 20266 29348 20322 29350
rect 20346 29348 20402 29350
rect 20426 29348 20482 29350
rect 27614 29402 27670 29404
rect 27694 29402 27750 29404
rect 27774 29402 27830 29404
rect 27854 29402 27910 29404
rect 27614 29350 27660 29402
rect 27660 29350 27670 29402
rect 27694 29350 27724 29402
rect 27724 29350 27736 29402
rect 27736 29350 27750 29402
rect 27774 29350 27788 29402
rect 27788 29350 27800 29402
rect 27800 29350 27830 29402
rect 27854 29350 27864 29402
rect 27864 29350 27910 29402
rect 27614 29348 27670 29350
rect 27694 29348 27750 29350
rect 27774 29348 27830 29350
rect 27854 29348 27910 29350
rect 4670 28858 4726 28860
rect 4750 28858 4806 28860
rect 4830 28858 4886 28860
rect 4910 28858 4966 28860
rect 4670 28806 4716 28858
rect 4716 28806 4726 28858
rect 4750 28806 4780 28858
rect 4780 28806 4792 28858
rect 4792 28806 4806 28858
rect 4830 28806 4844 28858
rect 4844 28806 4856 28858
rect 4856 28806 4886 28858
rect 4910 28806 4920 28858
rect 4920 28806 4966 28858
rect 4670 28804 4726 28806
rect 4750 28804 4806 28806
rect 4830 28804 4886 28806
rect 4910 28804 4966 28806
rect 12098 28858 12154 28860
rect 12178 28858 12234 28860
rect 12258 28858 12314 28860
rect 12338 28858 12394 28860
rect 12098 28806 12144 28858
rect 12144 28806 12154 28858
rect 12178 28806 12208 28858
rect 12208 28806 12220 28858
rect 12220 28806 12234 28858
rect 12258 28806 12272 28858
rect 12272 28806 12284 28858
rect 12284 28806 12314 28858
rect 12338 28806 12348 28858
rect 12348 28806 12394 28858
rect 12098 28804 12154 28806
rect 12178 28804 12234 28806
rect 12258 28804 12314 28806
rect 12338 28804 12394 28806
rect 5330 28314 5386 28316
rect 5410 28314 5466 28316
rect 5490 28314 5546 28316
rect 5570 28314 5626 28316
rect 5330 28262 5376 28314
rect 5376 28262 5386 28314
rect 5410 28262 5440 28314
rect 5440 28262 5452 28314
rect 5452 28262 5466 28314
rect 5490 28262 5504 28314
rect 5504 28262 5516 28314
rect 5516 28262 5546 28314
rect 5570 28262 5580 28314
rect 5580 28262 5626 28314
rect 5330 28260 5386 28262
rect 5410 28260 5466 28262
rect 5490 28260 5546 28262
rect 5570 28260 5626 28262
rect 4670 27770 4726 27772
rect 4750 27770 4806 27772
rect 4830 27770 4886 27772
rect 4910 27770 4966 27772
rect 4670 27718 4716 27770
rect 4716 27718 4726 27770
rect 4750 27718 4780 27770
rect 4780 27718 4792 27770
rect 4792 27718 4806 27770
rect 4830 27718 4844 27770
rect 4844 27718 4856 27770
rect 4856 27718 4886 27770
rect 4910 27718 4920 27770
rect 4920 27718 4966 27770
rect 4670 27716 4726 27718
rect 4750 27716 4806 27718
rect 4830 27716 4886 27718
rect 4910 27716 4966 27718
rect 12098 27770 12154 27772
rect 12178 27770 12234 27772
rect 12258 27770 12314 27772
rect 12338 27770 12394 27772
rect 12098 27718 12144 27770
rect 12144 27718 12154 27770
rect 12178 27718 12208 27770
rect 12208 27718 12220 27770
rect 12220 27718 12234 27770
rect 12258 27718 12272 27770
rect 12272 27718 12284 27770
rect 12284 27718 12314 27770
rect 12338 27718 12348 27770
rect 12348 27718 12394 27770
rect 12098 27716 12154 27718
rect 12178 27716 12234 27718
rect 12258 27716 12314 27718
rect 12338 27716 12394 27718
rect 5330 27226 5386 27228
rect 5410 27226 5466 27228
rect 5490 27226 5546 27228
rect 5570 27226 5626 27228
rect 5330 27174 5376 27226
rect 5376 27174 5386 27226
rect 5410 27174 5440 27226
rect 5440 27174 5452 27226
rect 5452 27174 5466 27226
rect 5490 27174 5504 27226
rect 5504 27174 5516 27226
rect 5516 27174 5546 27226
rect 5570 27174 5580 27226
rect 5580 27174 5626 27226
rect 5330 27172 5386 27174
rect 5410 27172 5466 27174
rect 5490 27172 5546 27174
rect 5570 27172 5626 27174
rect 4670 26682 4726 26684
rect 4750 26682 4806 26684
rect 4830 26682 4886 26684
rect 4910 26682 4966 26684
rect 4670 26630 4716 26682
rect 4716 26630 4726 26682
rect 4750 26630 4780 26682
rect 4780 26630 4792 26682
rect 4792 26630 4806 26682
rect 4830 26630 4844 26682
rect 4844 26630 4856 26682
rect 4856 26630 4886 26682
rect 4910 26630 4920 26682
rect 4920 26630 4966 26682
rect 4670 26628 4726 26630
rect 4750 26628 4806 26630
rect 4830 26628 4886 26630
rect 4910 26628 4966 26630
rect 12098 26682 12154 26684
rect 12178 26682 12234 26684
rect 12258 26682 12314 26684
rect 12338 26682 12394 26684
rect 12098 26630 12144 26682
rect 12144 26630 12154 26682
rect 12178 26630 12208 26682
rect 12208 26630 12220 26682
rect 12220 26630 12234 26682
rect 12258 26630 12272 26682
rect 12272 26630 12284 26682
rect 12284 26630 12314 26682
rect 12338 26630 12348 26682
rect 12348 26630 12394 26682
rect 12098 26628 12154 26630
rect 12178 26628 12234 26630
rect 12258 26628 12314 26630
rect 12338 26628 12394 26630
rect 5330 26138 5386 26140
rect 5410 26138 5466 26140
rect 5490 26138 5546 26140
rect 5570 26138 5626 26140
rect 5330 26086 5376 26138
rect 5376 26086 5386 26138
rect 5410 26086 5440 26138
rect 5440 26086 5452 26138
rect 5452 26086 5466 26138
rect 5490 26086 5504 26138
rect 5504 26086 5516 26138
rect 5516 26086 5546 26138
rect 5570 26086 5580 26138
rect 5580 26086 5626 26138
rect 5330 26084 5386 26086
rect 5410 26084 5466 26086
rect 5490 26084 5546 26086
rect 5570 26084 5626 26086
rect 4670 25594 4726 25596
rect 4750 25594 4806 25596
rect 4830 25594 4886 25596
rect 4910 25594 4966 25596
rect 4670 25542 4716 25594
rect 4716 25542 4726 25594
rect 4750 25542 4780 25594
rect 4780 25542 4792 25594
rect 4792 25542 4806 25594
rect 4830 25542 4844 25594
rect 4844 25542 4856 25594
rect 4856 25542 4886 25594
rect 4910 25542 4920 25594
rect 4920 25542 4966 25594
rect 4670 25540 4726 25542
rect 4750 25540 4806 25542
rect 4830 25540 4886 25542
rect 4910 25540 4966 25542
rect 12098 25594 12154 25596
rect 12178 25594 12234 25596
rect 12258 25594 12314 25596
rect 12338 25594 12394 25596
rect 12098 25542 12144 25594
rect 12144 25542 12154 25594
rect 12178 25542 12208 25594
rect 12208 25542 12220 25594
rect 12220 25542 12234 25594
rect 12258 25542 12272 25594
rect 12272 25542 12284 25594
rect 12284 25542 12314 25594
rect 12338 25542 12348 25594
rect 12348 25542 12394 25594
rect 12098 25540 12154 25542
rect 12178 25540 12234 25542
rect 12258 25540 12314 25542
rect 12338 25540 12394 25542
rect 3422 25200 3478 25256
rect 1490 23432 1546 23488
rect 938 22500 994 22536
rect 938 22480 940 22500
rect 940 22480 992 22500
rect 992 22480 994 22500
rect 938 21836 940 21856
rect 940 21836 992 21856
rect 992 21836 994 21856
rect 938 21800 994 21836
rect 938 21120 994 21176
rect 1490 20576 1546 20632
rect 938 19780 994 19816
rect 938 19760 940 19780
rect 940 19760 992 19780
rect 992 19760 994 19780
rect 1398 19216 1454 19272
rect 938 18400 994 18456
rect 1490 17856 1546 17912
rect 938 17076 940 17096
rect 940 17076 992 17096
rect 992 17076 994 17096
rect 938 17040 994 17076
rect 5330 25050 5386 25052
rect 5410 25050 5466 25052
rect 5490 25050 5546 25052
rect 5570 25050 5626 25052
rect 5330 24998 5376 25050
rect 5376 24998 5386 25050
rect 5410 24998 5440 25050
rect 5440 24998 5452 25050
rect 5452 24998 5466 25050
rect 5490 24998 5504 25050
rect 5504 24998 5516 25050
rect 5516 24998 5546 25050
rect 5570 24998 5580 25050
rect 5580 24998 5626 25050
rect 5330 24996 5386 24998
rect 5410 24996 5466 24998
rect 5490 24996 5546 24998
rect 5570 24996 5626 24998
rect 4670 24506 4726 24508
rect 4750 24506 4806 24508
rect 4830 24506 4886 24508
rect 4910 24506 4966 24508
rect 4670 24454 4716 24506
rect 4716 24454 4726 24506
rect 4750 24454 4780 24506
rect 4780 24454 4792 24506
rect 4792 24454 4806 24506
rect 4830 24454 4844 24506
rect 4844 24454 4856 24506
rect 4856 24454 4886 24506
rect 4910 24454 4920 24506
rect 4920 24454 4966 24506
rect 4670 24452 4726 24454
rect 4750 24452 4806 24454
rect 4830 24452 4886 24454
rect 4910 24452 4966 24454
rect 12098 24506 12154 24508
rect 12178 24506 12234 24508
rect 12258 24506 12314 24508
rect 12338 24506 12394 24508
rect 12098 24454 12144 24506
rect 12144 24454 12154 24506
rect 12178 24454 12208 24506
rect 12208 24454 12220 24506
rect 12220 24454 12234 24506
rect 12258 24454 12272 24506
rect 12272 24454 12284 24506
rect 12284 24454 12314 24506
rect 12338 24454 12348 24506
rect 12348 24454 12394 24506
rect 12098 24452 12154 24454
rect 12178 24452 12234 24454
rect 12258 24452 12314 24454
rect 12338 24452 12394 24454
rect 5330 23962 5386 23964
rect 5410 23962 5466 23964
rect 5490 23962 5546 23964
rect 5570 23962 5626 23964
rect 5330 23910 5376 23962
rect 5376 23910 5386 23962
rect 5410 23910 5440 23962
rect 5440 23910 5452 23962
rect 5452 23910 5466 23962
rect 5490 23910 5504 23962
rect 5504 23910 5516 23962
rect 5516 23910 5546 23962
rect 5570 23910 5580 23962
rect 5580 23910 5626 23962
rect 5330 23908 5386 23910
rect 5410 23908 5466 23910
rect 5490 23908 5546 23910
rect 5570 23908 5626 23910
rect 4670 23418 4726 23420
rect 4750 23418 4806 23420
rect 4830 23418 4886 23420
rect 4910 23418 4966 23420
rect 4670 23366 4716 23418
rect 4716 23366 4726 23418
rect 4750 23366 4780 23418
rect 4780 23366 4792 23418
rect 4792 23366 4806 23418
rect 4830 23366 4844 23418
rect 4844 23366 4856 23418
rect 4856 23366 4886 23418
rect 4910 23366 4920 23418
rect 4920 23366 4966 23418
rect 4670 23364 4726 23366
rect 4750 23364 4806 23366
rect 4830 23364 4886 23366
rect 4910 23364 4966 23366
rect 5330 22874 5386 22876
rect 5410 22874 5466 22876
rect 5490 22874 5546 22876
rect 5570 22874 5626 22876
rect 5330 22822 5376 22874
rect 5376 22822 5386 22874
rect 5410 22822 5440 22874
rect 5440 22822 5452 22874
rect 5452 22822 5466 22874
rect 5490 22822 5504 22874
rect 5504 22822 5516 22874
rect 5516 22822 5546 22874
rect 5570 22822 5580 22874
rect 5580 22822 5626 22874
rect 5330 22820 5386 22822
rect 5410 22820 5466 22822
rect 5490 22820 5546 22822
rect 5570 22820 5626 22822
rect 4670 22330 4726 22332
rect 4750 22330 4806 22332
rect 4830 22330 4886 22332
rect 4910 22330 4966 22332
rect 4670 22278 4716 22330
rect 4716 22278 4726 22330
rect 4750 22278 4780 22330
rect 4780 22278 4792 22330
rect 4792 22278 4806 22330
rect 4830 22278 4844 22330
rect 4844 22278 4856 22330
rect 4856 22278 4886 22330
rect 4910 22278 4920 22330
rect 4920 22278 4966 22330
rect 4670 22276 4726 22278
rect 4750 22276 4806 22278
rect 4830 22276 4886 22278
rect 4910 22276 4966 22278
rect 4670 21242 4726 21244
rect 4750 21242 4806 21244
rect 4830 21242 4886 21244
rect 4910 21242 4966 21244
rect 4670 21190 4716 21242
rect 4716 21190 4726 21242
rect 4750 21190 4780 21242
rect 4780 21190 4792 21242
rect 4792 21190 4806 21242
rect 4830 21190 4844 21242
rect 4844 21190 4856 21242
rect 4856 21190 4886 21242
rect 4910 21190 4920 21242
rect 4920 21190 4966 21242
rect 4670 21188 4726 21190
rect 4750 21188 4806 21190
rect 4830 21188 4886 21190
rect 4910 21188 4966 21190
rect 5330 21786 5386 21788
rect 5410 21786 5466 21788
rect 5490 21786 5546 21788
rect 5570 21786 5626 21788
rect 5330 21734 5376 21786
rect 5376 21734 5386 21786
rect 5410 21734 5440 21786
rect 5440 21734 5452 21786
rect 5452 21734 5466 21786
rect 5490 21734 5504 21786
rect 5504 21734 5516 21786
rect 5516 21734 5546 21786
rect 5570 21734 5580 21786
rect 5580 21734 5626 21786
rect 5330 21732 5386 21734
rect 5410 21732 5466 21734
rect 5490 21732 5546 21734
rect 5570 21732 5626 21734
rect 5330 20698 5386 20700
rect 5410 20698 5466 20700
rect 5490 20698 5546 20700
rect 5570 20698 5626 20700
rect 5330 20646 5376 20698
rect 5376 20646 5386 20698
rect 5410 20646 5440 20698
rect 5440 20646 5452 20698
rect 5452 20646 5466 20698
rect 5490 20646 5504 20698
rect 5504 20646 5516 20698
rect 5516 20646 5546 20698
rect 5570 20646 5580 20698
rect 5580 20646 5626 20698
rect 5330 20644 5386 20646
rect 5410 20644 5466 20646
rect 5490 20644 5546 20646
rect 5570 20644 5626 20646
rect 4670 20154 4726 20156
rect 4750 20154 4806 20156
rect 4830 20154 4886 20156
rect 4910 20154 4966 20156
rect 4670 20102 4716 20154
rect 4716 20102 4726 20154
rect 4750 20102 4780 20154
rect 4780 20102 4792 20154
rect 4792 20102 4806 20154
rect 4830 20102 4844 20154
rect 4844 20102 4856 20154
rect 4856 20102 4886 20154
rect 4910 20102 4920 20154
rect 4920 20102 4966 20154
rect 4670 20100 4726 20102
rect 4750 20100 4806 20102
rect 4830 20100 4886 20102
rect 4910 20100 4966 20102
rect 5330 19610 5386 19612
rect 5410 19610 5466 19612
rect 5490 19610 5546 19612
rect 5570 19610 5626 19612
rect 5330 19558 5376 19610
rect 5376 19558 5386 19610
rect 5410 19558 5440 19610
rect 5440 19558 5452 19610
rect 5452 19558 5466 19610
rect 5490 19558 5504 19610
rect 5504 19558 5516 19610
rect 5516 19558 5546 19610
rect 5570 19558 5580 19610
rect 5580 19558 5626 19610
rect 5330 19556 5386 19558
rect 5410 19556 5466 19558
rect 5490 19556 5546 19558
rect 5570 19556 5626 19558
rect 938 16396 940 16416
rect 940 16396 992 16416
rect 992 16396 994 16416
rect 938 16360 994 16396
rect 938 15680 994 15736
rect 4670 19066 4726 19068
rect 4750 19066 4806 19068
rect 4830 19066 4886 19068
rect 4910 19066 4966 19068
rect 4670 19014 4716 19066
rect 4716 19014 4726 19066
rect 4750 19014 4780 19066
rect 4780 19014 4792 19066
rect 4792 19014 4806 19066
rect 4830 19014 4844 19066
rect 4844 19014 4856 19066
rect 4856 19014 4886 19066
rect 4910 19014 4920 19066
rect 4920 19014 4966 19066
rect 4670 19012 4726 19014
rect 4750 19012 4806 19014
rect 4830 19012 4886 19014
rect 4910 19012 4966 19014
rect 4670 17978 4726 17980
rect 4750 17978 4806 17980
rect 4830 17978 4886 17980
rect 4910 17978 4966 17980
rect 4670 17926 4716 17978
rect 4716 17926 4726 17978
rect 4750 17926 4780 17978
rect 4780 17926 4792 17978
rect 4792 17926 4806 17978
rect 4830 17926 4844 17978
rect 4844 17926 4856 17978
rect 4856 17926 4886 17978
rect 4910 17926 4920 17978
rect 4920 17926 4966 17978
rect 4670 17924 4726 17926
rect 4750 17924 4806 17926
rect 4830 17924 4886 17926
rect 4910 17924 4966 17926
rect 5330 18522 5386 18524
rect 5410 18522 5466 18524
rect 5490 18522 5546 18524
rect 5570 18522 5626 18524
rect 5330 18470 5376 18522
rect 5376 18470 5386 18522
rect 5410 18470 5440 18522
rect 5440 18470 5452 18522
rect 5452 18470 5466 18522
rect 5490 18470 5504 18522
rect 5504 18470 5516 18522
rect 5516 18470 5546 18522
rect 5570 18470 5580 18522
rect 5580 18470 5626 18522
rect 5330 18468 5386 18470
rect 5410 18468 5466 18470
rect 5490 18468 5546 18470
rect 5570 18468 5626 18470
rect 5330 17434 5386 17436
rect 5410 17434 5466 17436
rect 5490 17434 5546 17436
rect 5570 17434 5626 17436
rect 5330 17382 5376 17434
rect 5376 17382 5386 17434
rect 5410 17382 5440 17434
rect 5440 17382 5452 17434
rect 5452 17382 5466 17434
rect 5490 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5546 17434
rect 5570 17382 5580 17434
rect 5580 17382 5626 17434
rect 5330 17380 5386 17382
rect 5410 17380 5466 17382
rect 5490 17380 5546 17382
rect 5570 17380 5626 17382
rect 5722 17196 5778 17232
rect 5722 17176 5724 17196
rect 5724 17176 5776 17196
rect 5776 17176 5778 17196
rect 4670 16890 4726 16892
rect 4750 16890 4806 16892
rect 4830 16890 4886 16892
rect 4910 16890 4966 16892
rect 4670 16838 4716 16890
rect 4716 16838 4726 16890
rect 4750 16838 4780 16890
rect 4780 16838 4792 16890
rect 4792 16838 4806 16890
rect 4830 16838 4844 16890
rect 4844 16838 4856 16890
rect 4856 16838 4886 16890
rect 4910 16838 4920 16890
rect 4920 16838 4966 16890
rect 4670 16836 4726 16838
rect 4750 16836 4806 16838
rect 4830 16836 4886 16838
rect 4910 16836 4966 16838
rect 5330 16346 5386 16348
rect 5410 16346 5466 16348
rect 5490 16346 5546 16348
rect 5570 16346 5626 16348
rect 5330 16294 5376 16346
rect 5376 16294 5386 16346
rect 5410 16294 5440 16346
rect 5440 16294 5452 16346
rect 5452 16294 5466 16346
rect 5490 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5546 16346
rect 5570 16294 5580 16346
rect 5580 16294 5626 16346
rect 5330 16292 5386 16294
rect 5410 16292 5466 16294
rect 5490 16292 5546 16294
rect 5570 16292 5626 16294
rect 4670 15802 4726 15804
rect 4750 15802 4806 15804
rect 4830 15802 4886 15804
rect 4910 15802 4966 15804
rect 4670 15750 4716 15802
rect 4716 15750 4726 15802
rect 4750 15750 4780 15802
rect 4780 15750 4792 15802
rect 4792 15750 4806 15802
rect 4830 15750 4844 15802
rect 4844 15750 4856 15802
rect 4856 15750 4886 15802
rect 4910 15750 4920 15802
rect 4920 15750 4966 15802
rect 4670 15748 4726 15750
rect 4750 15748 4806 15750
rect 4830 15748 4886 15750
rect 4910 15748 4966 15750
rect 1398 15136 1454 15192
rect 938 14320 994 14376
rect 1398 13640 1454 13696
rect 938 12960 994 13016
rect 1490 12280 1546 12336
rect 938 11600 994 11656
rect 5330 15258 5386 15260
rect 5410 15258 5466 15260
rect 5490 15258 5546 15260
rect 5570 15258 5626 15260
rect 5330 15206 5376 15258
rect 5376 15206 5386 15258
rect 5410 15206 5440 15258
rect 5440 15206 5452 15258
rect 5452 15206 5466 15258
rect 5490 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5546 15258
rect 5570 15206 5580 15258
rect 5580 15206 5626 15258
rect 5330 15204 5386 15206
rect 5410 15204 5466 15206
rect 5490 15204 5546 15206
rect 5570 15204 5626 15206
rect 4670 14714 4726 14716
rect 4750 14714 4806 14716
rect 4830 14714 4886 14716
rect 4910 14714 4966 14716
rect 4670 14662 4716 14714
rect 4716 14662 4726 14714
rect 4750 14662 4780 14714
rect 4780 14662 4792 14714
rect 4792 14662 4806 14714
rect 4830 14662 4844 14714
rect 4844 14662 4856 14714
rect 4856 14662 4886 14714
rect 4910 14662 4920 14714
rect 4920 14662 4966 14714
rect 4670 14660 4726 14662
rect 4750 14660 4806 14662
rect 4830 14660 4886 14662
rect 4910 14660 4966 14662
rect 6274 17196 6330 17232
rect 6274 17176 6276 17196
rect 6276 17176 6328 17196
rect 6328 17176 6330 17196
rect 12098 23418 12154 23420
rect 12178 23418 12234 23420
rect 12258 23418 12314 23420
rect 12338 23418 12394 23420
rect 12098 23366 12144 23418
rect 12144 23366 12154 23418
rect 12178 23366 12208 23418
rect 12208 23366 12220 23418
rect 12220 23366 12234 23418
rect 12258 23366 12272 23418
rect 12272 23366 12284 23418
rect 12284 23366 12314 23418
rect 12338 23366 12348 23418
rect 12348 23366 12394 23418
rect 12098 23364 12154 23366
rect 12178 23364 12234 23366
rect 12258 23364 12314 23366
rect 12338 23364 12394 23366
rect 12098 22330 12154 22332
rect 12178 22330 12234 22332
rect 12258 22330 12314 22332
rect 12338 22330 12394 22332
rect 12098 22278 12144 22330
rect 12144 22278 12154 22330
rect 12178 22278 12208 22330
rect 12208 22278 12220 22330
rect 12220 22278 12234 22330
rect 12258 22278 12272 22330
rect 12272 22278 12284 22330
rect 12284 22278 12314 22330
rect 12338 22278 12348 22330
rect 12348 22278 12394 22330
rect 12098 22276 12154 22278
rect 12178 22276 12234 22278
rect 12258 22276 12314 22278
rect 12338 22276 12394 22278
rect 5330 14170 5386 14172
rect 5410 14170 5466 14172
rect 5490 14170 5546 14172
rect 5570 14170 5626 14172
rect 5330 14118 5376 14170
rect 5376 14118 5386 14170
rect 5410 14118 5440 14170
rect 5440 14118 5452 14170
rect 5452 14118 5466 14170
rect 5490 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5546 14170
rect 5570 14118 5580 14170
rect 5580 14118 5626 14170
rect 5330 14116 5386 14118
rect 5410 14116 5466 14118
rect 5490 14116 5546 14118
rect 5570 14116 5626 14118
rect 4670 13626 4726 13628
rect 4750 13626 4806 13628
rect 4830 13626 4886 13628
rect 4910 13626 4966 13628
rect 4670 13574 4716 13626
rect 4716 13574 4726 13626
rect 4750 13574 4780 13626
rect 4780 13574 4792 13626
rect 4792 13574 4806 13626
rect 4830 13574 4844 13626
rect 4844 13574 4856 13626
rect 4856 13574 4886 13626
rect 4910 13574 4920 13626
rect 4920 13574 4966 13626
rect 4670 13572 4726 13574
rect 4750 13572 4806 13574
rect 4830 13572 4886 13574
rect 4910 13572 4966 13574
rect 5330 13082 5386 13084
rect 5410 13082 5466 13084
rect 5490 13082 5546 13084
rect 5570 13082 5626 13084
rect 5330 13030 5376 13082
rect 5376 13030 5386 13082
rect 5410 13030 5440 13082
rect 5440 13030 5452 13082
rect 5452 13030 5466 13082
rect 5490 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5546 13082
rect 5570 13030 5580 13082
rect 5580 13030 5626 13082
rect 5330 13028 5386 13030
rect 5410 13028 5466 13030
rect 5490 13028 5546 13030
rect 5570 13028 5626 13030
rect 4670 12538 4726 12540
rect 4750 12538 4806 12540
rect 4830 12538 4886 12540
rect 4910 12538 4966 12540
rect 4670 12486 4716 12538
rect 4716 12486 4726 12538
rect 4750 12486 4780 12538
rect 4780 12486 4792 12538
rect 4792 12486 4806 12538
rect 4830 12486 4844 12538
rect 4844 12486 4856 12538
rect 4856 12486 4886 12538
rect 4910 12486 4920 12538
rect 4920 12486 4966 12538
rect 4670 12484 4726 12486
rect 4750 12484 4806 12486
rect 4830 12484 4886 12486
rect 4910 12484 4966 12486
rect 5330 11994 5386 11996
rect 5410 11994 5466 11996
rect 5490 11994 5546 11996
rect 5570 11994 5626 11996
rect 5330 11942 5376 11994
rect 5376 11942 5386 11994
rect 5410 11942 5440 11994
rect 5440 11942 5452 11994
rect 5452 11942 5466 11994
rect 5490 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5546 11994
rect 5570 11942 5580 11994
rect 5580 11942 5626 11994
rect 5330 11940 5386 11942
rect 5410 11940 5466 11942
rect 5490 11940 5546 11942
rect 5570 11940 5626 11942
rect 4670 11450 4726 11452
rect 4750 11450 4806 11452
rect 4830 11450 4886 11452
rect 4910 11450 4966 11452
rect 4670 11398 4716 11450
rect 4716 11398 4726 11450
rect 4750 11398 4780 11450
rect 4780 11398 4792 11450
rect 4792 11398 4806 11450
rect 4830 11398 4844 11450
rect 4844 11398 4856 11450
rect 4856 11398 4886 11450
rect 4910 11398 4920 11450
rect 4920 11398 4966 11450
rect 4670 11396 4726 11398
rect 4750 11396 4806 11398
rect 4830 11396 4886 11398
rect 4910 11396 4966 11398
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 938 10240 994 10296
rect 1490 9560 1546 9616
rect 5330 10906 5386 10908
rect 5410 10906 5466 10908
rect 5490 10906 5546 10908
rect 5570 10906 5626 10908
rect 5330 10854 5376 10906
rect 5376 10854 5386 10906
rect 5410 10854 5440 10906
rect 5440 10854 5452 10906
rect 5452 10854 5466 10906
rect 5490 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5546 10906
rect 5570 10854 5580 10906
rect 5580 10854 5626 10906
rect 5330 10852 5386 10854
rect 5410 10852 5466 10854
rect 5490 10852 5546 10854
rect 5570 10852 5626 10854
rect 4670 10362 4726 10364
rect 4750 10362 4806 10364
rect 4830 10362 4886 10364
rect 4910 10362 4966 10364
rect 4670 10310 4716 10362
rect 4716 10310 4726 10362
rect 4750 10310 4780 10362
rect 4780 10310 4792 10362
rect 4792 10310 4806 10362
rect 4830 10310 4844 10362
rect 4844 10310 4856 10362
rect 4856 10310 4886 10362
rect 4910 10310 4920 10362
rect 4920 10310 4966 10362
rect 4670 10308 4726 10310
rect 4750 10308 4806 10310
rect 4830 10308 4886 10310
rect 4910 10308 4966 10310
rect 5330 9818 5386 9820
rect 5410 9818 5466 9820
rect 5490 9818 5546 9820
rect 5570 9818 5626 9820
rect 5330 9766 5376 9818
rect 5376 9766 5386 9818
rect 5410 9766 5440 9818
rect 5440 9766 5452 9818
rect 5452 9766 5466 9818
rect 5490 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5546 9818
rect 5570 9766 5580 9818
rect 5580 9766 5626 9818
rect 5330 9764 5386 9766
rect 5410 9764 5466 9766
rect 5490 9764 5546 9766
rect 5570 9764 5626 9766
rect 4670 9274 4726 9276
rect 4750 9274 4806 9276
rect 4830 9274 4886 9276
rect 4910 9274 4966 9276
rect 4670 9222 4716 9274
rect 4716 9222 4726 9274
rect 4750 9222 4780 9274
rect 4780 9222 4792 9274
rect 4792 9222 4806 9274
rect 4830 9222 4844 9274
rect 4844 9222 4856 9274
rect 4856 9222 4886 9274
rect 4910 9222 4920 9274
rect 4920 9222 4966 9274
rect 4670 9220 4726 9222
rect 4750 9220 4806 9222
rect 4830 9220 4886 9222
rect 4910 9220 4966 9222
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 1398 8200 1454 8256
rect 4670 8186 4726 8188
rect 4750 8186 4806 8188
rect 4830 8186 4886 8188
rect 4910 8186 4966 8188
rect 4670 8134 4716 8186
rect 4716 8134 4726 8186
rect 4750 8134 4780 8186
rect 4780 8134 4792 8186
rect 4792 8134 4806 8186
rect 4830 8134 4844 8186
rect 4844 8134 4856 8186
rect 4856 8134 4886 8186
rect 4910 8134 4920 8186
rect 4920 8134 4966 8186
rect 4670 8132 4726 8134
rect 4750 8132 4806 8134
rect 4830 8132 4886 8134
rect 4910 8132 4966 8134
rect 938 7520 994 7576
rect 5330 8730 5386 8732
rect 5410 8730 5466 8732
rect 5490 8730 5546 8732
rect 5570 8730 5626 8732
rect 5330 8678 5376 8730
rect 5376 8678 5386 8730
rect 5410 8678 5440 8730
rect 5440 8678 5452 8730
rect 5452 8678 5466 8730
rect 5490 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5546 8730
rect 5570 8678 5580 8730
rect 5580 8678 5626 8730
rect 5330 8676 5386 8678
rect 5410 8676 5466 8678
rect 5490 8676 5546 8678
rect 5570 8676 5626 8678
rect 5998 8744 6054 8800
rect 10506 16532 10508 16552
rect 10508 16532 10560 16552
rect 10560 16532 10562 16552
rect 10506 16496 10562 16532
rect 12098 21242 12154 21244
rect 12178 21242 12234 21244
rect 12258 21242 12314 21244
rect 12338 21242 12394 21244
rect 12098 21190 12144 21242
rect 12144 21190 12154 21242
rect 12178 21190 12208 21242
rect 12208 21190 12220 21242
rect 12220 21190 12234 21242
rect 12258 21190 12272 21242
rect 12272 21190 12284 21242
rect 12284 21190 12314 21242
rect 12338 21190 12348 21242
rect 12348 21190 12394 21242
rect 12098 21188 12154 21190
rect 12178 21188 12234 21190
rect 12258 21188 12314 21190
rect 12338 21188 12394 21190
rect 12758 28314 12814 28316
rect 12838 28314 12894 28316
rect 12918 28314 12974 28316
rect 12998 28314 13054 28316
rect 12758 28262 12804 28314
rect 12804 28262 12814 28314
rect 12838 28262 12868 28314
rect 12868 28262 12880 28314
rect 12880 28262 12894 28314
rect 12918 28262 12932 28314
rect 12932 28262 12944 28314
rect 12944 28262 12974 28314
rect 12998 28262 13008 28314
rect 13008 28262 13054 28314
rect 12758 28260 12814 28262
rect 12838 28260 12894 28262
rect 12918 28260 12974 28262
rect 12998 28260 13054 28262
rect 12758 27226 12814 27228
rect 12838 27226 12894 27228
rect 12918 27226 12974 27228
rect 12998 27226 13054 27228
rect 12758 27174 12804 27226
rect 12804 27174 12814 27226
rect 12838 27174 12868 27226
rect 12868 27174 12880 27226
rect 12880 27174 12894 27226
rect 12918 27174 12932 27226
rect 12932 27174 12944 27226
rect 12944 27174 12974 27226
rect 12998 27174 13008 27226
rect 13008 27174 13054 27226
rect 12758 27172 12814 27174
rect 12838 27172 12894 27174
rect 12918 27172 12974 27174
rect 12998 27172 13054 27174
rect 12758 26138 12814 26140
rect 12838 26138 12894 26140
rect 12918 26138 12974 26140
rect 12998 26138 13054 26140
rect 12758 26086 12804 26138
rect 12804 26086 12814 26138
rect 12838 26086 12868 26138
rect 12868 26086 12880 26138
rect 12880 26086 12894 26138
rect 12918 26086 12932 26138
rect 12932 26086 12944 26138
rect 12944 26086 12974 26138
rect 12998 26086 13008 26138
rect 13008 26086 13054 26138
rect 12758 26084 12814 26086
rect 12838 26084 12894 26086
rect 12918 26084 12974 26086
rect 12998 26084 13054 26086
rect 12758 25050 12814 25052
rect 12838 25050 12894 25052
rect 12918 25050 12974 25052
rect 12998 25050 13054 25052
rect 12758 24998 12804 25050
rect 12804 24998 12814 25050
rect 12838 24998 12868 25050
rect 12868 24998 12880 25050
rect 12880 24998 12894 25050
rect 12918 24998 12932 25050
rect 12932 24998 12944 25050
rect 12944 24998 12974 25050
rect 12998 24998 13008 25050
rect 13008 24998 13054 25050
rect 12758 24996 12814 24998
rect 12838 24996 12894 24998
rect 12918 24996 12974 24998
rect 12998 24996 13054 24998
rect 12758 23962 12814 23964
rect 12838 23962 12894 23964
rect 12918 23962 12974 23964
rect 12998 23962 13054 23964
rect 12758 23910 12804 23962
rect 12804 23910 12814 23962
rect 12838 23910 12868 23962
rect 12868 23910 12880 23962
rect 12880 23910 12894 23962
rect 12918 23910 12932 23962
rect 12932 23910 12944 23962
rect 12944 23910 12974 23962
rect 12998 23910 13008 23962
rect 13008 23910 13054 23962
rect 12758 23908 12814 23910
rect 12838 23908 12894 23910
rect 12918 23908 12974 23910
rect 12998 23908 13054 23910
rect 12758 22874 12814 22876
rect 12838 22874 12894 22876
rect 12918 22874 12974 22876
rect 12998 22874 13054 22876
rect 12758 22822 12804 22874
rect 12804 22822 12814 22874
rect 12838 22822 12868 22874
rect 12868 22822 12880 22874
rect 12880 22822 12894 22874
rect 12918 22822 12932 22874
rect 12932 22822 12944 22874
rect 12944 22822 12974 22874
rect 12998 22822 13008 22874
rect 13008 22822 13054 22874
rect 12758 22820 12814 22822
rect 12838 22820 12894 22822
rect 12918 22820 12974 22822
rect 12998 22820 13054 22822
rect 12758 21786 12814 21788
rect 12838 21786 12894 21788
rect 12918 21786 12974 21788
rect 12998 21786 13054 21788
rect 12758 21734 12804 21786
rect 12804 21734 12814 21786
rect 12838 21734 12868 21786
rect 12868 21734 12880 21786
rect 12880 21734 12894 21786
rect 12918 21734 12932 21786
rect 12932 21734 12944 21786
rect 12944 21734 12974 21786
rect 12998 21734 13008 21786
rect 13008 21734 13054 21786
rect 12758 21732 12814 21734
rect 12838 21732 12894 21734
rect 12918 21732 12974 21734
rect 12998 21732 13054 21734
rect 12758 20698 12814 20700
rect 12838 20698 12894 20700
rect 12918 20698 12974 20700
rect 12998 20698 13054 20700
rect 12758 20646 12804 20698
rect 12804 20646 12814 20698
rect 12838 20646 12868 20698
rect 12868 20646 12880 20698
rect 12880 20646 12894 20698
rect 12918 20646 12932 20698
rect 12932 20646 12944 20698
rect 12944 20646 12974 20698
rect 12998 20646 13008 20698
rect 13008 20646 13054 20698
rect 12758 20644 12814 20646
rect 12838 20644 12894 20646
rect 12918 20644 12974 20646
rect 12998 20644 13054 20646
rect 12098 20154 12154 20156
rect 12178 20154 12234 20156
rect 12258 20154 12314 20156
rect 12338 20154 12394 20156
rect 12098 20102 12144 20154
rect 12144 20102 12154 20154
rect 12178 20102 12208 20154
rect 12208 20102 12220 20154
rect 12220 20102 12234 20154
rect 12258 20102 12272 20154
rect 12272 20102 12284 20154
rect 12284 20102 12314 20154
rect 12338 20102 12348 20154
rect 12348 20102 12394 20154
rect 12098 20100 12154 20102
rect 12178 20100 12234 20102
rect 12258 20100 12314 20102
rect 12338 20100 12394 20102
rect 12758 19610 12814 19612
rect 12838 19610 12894 19612
rect 12918 19610 12974 19612
rect 12998 19610 13054 19612
rect 12758 19558 12804 19610
rect 12804 19558 12814 19610
rect 12838 19558 12868 19610
rect 12868 19558 12880 19610
rect 12880 19558 12894 19610
rect 12918 19558 12932 19610
rect 12932 19558 12944 19610
rect 12944 19558 12974 19610
rect 12998 19558 13008 19610
rect 13008 19558 13054 19610
rect 12758 19556 12814 19558
rect 12838 19556 12894 19558
rect 12918 19556 12974 19558
rect 12998 19556 13054 19558
rect 12098 19066 12154 19068
rect 12178 19066 12234 19068
rect 12258 19066 12314 19068
rect 12338 19066 12394 19068
rect 12098 19014 12144 19066
rect 12144 19014 12154 19066
rect 12178 19014 12208 19066
rect 12208 19014 12220 19066
rect 12220 19014 12234 19066
rect 12258 19014 12272 19066
rect 12272 19014 12284 19066
rect 12284 19014 12314 19066
rect 12338 19014 12348 19066
rect 12348 19014 12394 19066
rect 12098 19012 12154 19014
rect 12178 19012 12234 19014
rect 12258 19012 12314 19014
rect 12338 19012 12394 19014
rect 11978 18264 12034 18320
rect 12098 17978 12154 17980
rect 12178 17978 12234 17980
rect 12258 17978 12314 17980
rect 12338 17978 12394 17980
rect 12098 17926 12144 17978
rect 12144 17926 12154 17978
rect 12178 17926 12208 17978
rect 12208 17926 12220 17978
rect 12220 17926 12234 17978
rect 12258 17926 12272 17978
rect 12272 17926 12284 17978
rect 12284 17926 12314 17978
rect 12338 17926 12348 17978
rect 12348 17926 12394 17978
rect 12098 17924 12154 17926
rect 12178 17924 12234 17926
rect 12258 17924 12314 17926
rect 12338 17924 12394 17926
rect 12758 18522 12814 18524
rect 12838 18522 12894 18524
rect 12918 18522 12974 18524
rect 12998 18522 13054 18524
rect 12758 18470 12804 18522
rect 12804 18470 12814 18522
rect 12838 18470 12868 18522
rect 12868 18470 12880 18522
rect 12880 18470 12894 18522
rect 12918 18470 12932 18522
rect 12932 18470 12944 18522
rect 12944 18470 12974 18522
rect 12998 18470 13008 18522
rect 13008 18470 13054 18522
rect 12758 18468 12814 18470
rect 12838 18468 12894 18470
rect 12918 18468 12974 18470
rect 12998 18468 13054 18470
rect 12758 17434 12814 17436
rect 12838 17434 12894 17436
rect 12918 17434 12974 17436
rect 12998 17434 13054 17436
rect 12758 17382 12804 17434
rect 12804 17382 12814 17434
rect 12838 17382 12868 17434
rect 12868 17382 12880 17434
rect 12880 17382 12894 17434
rect 12918 17382 12932 17434
rect 12932 17382 12944 17434
rect 12944 17382 12974 17434
rect 12998 17382 13008 17434
rect 13008 17382 13054 17434
rect 12758 17380 12814 17382
rect 12838 17380 12894 17382
rect 12918 17380 12974 17382
rect 12998 17380 13054 17382
rect 12098 16890 12154 16892
rect 12178 16890 12234 16892
rect 12258 16890 12314 16892
rect 12338 16890 12394 16892
rect 12098 16838 12144 16890
rect 12144 16838 12154 16890
rect 12178 16838 12208 16890
rect 12208 16838 12220 16890
rect 12220 16838 12234 16890
rect 12258 16838 12272 16890
rect 12272 16838 12284 16890
rect 12284 16838 12314 16890
rect 12338 16838 12348 16890
rect 12348 16838 12394 16890
rect 12098 16836 12154 16838
rect 12178 16836 12234 16838
rect 12258 16836 12314 16838
rect 12338 16836 12394 16838
rect 12758 16346 12814 16348
rect 12838 16346 12894 16348
rect 12918 16346 12974 16348
rect 12998 16346 13054 16348
rect 12758 16294 12804 16346
rect 12804 16294 12814 16346
rect 12838 16294 12868 16346
rect 12868 16294 12880 16346
rect 12880 16294 12894 16346
rect 12918 16294 12932 16346
rect 12932 16294 12944 16346
rect 12944 16294 12974 16346
rect 12998 16294 13008 16346
rect 13008 16294 13054 16346
rect 12758 16292 12814 16294
rect 12838 16292 12894 16294
rect 12918 16292 12974 16294
rect 12998 16292 13054 16294
rect 12098 15802 12154 15804
rect 12178 15802 12234 15804
rect 12258 15802 12314 15804
rect 12338 15802 12394 15804
rect 12098 15750 12144 15802
rect 12144 15750 12154 15802
rect 12178 15750 12208 15802
rect 12208 15750 12220 15802
rect 12220 15750 12234 15802
rect 12258 15750 12272 15802
rect 12272 15750 12284 15802
rect 12284 15750 12314 15802
rect 12338 15750 12348 15802
rect 12348 15750 12394 15802
rect 12098 15748 12154 15750
rect 12178 15748 12234 15750
rect 12258 15748 12314 15750
rect 12338 15748 12394 15750
rect 12758 15258 12814 15260
rect 12838 15258 12894 15260
rect 12918 15258 12974 15260
rect 12998 15258 13054 15260
rect 12758 15206 12804 15258
rect 12804 15206 12814 15258
rect 12838 15206 12868 15258
rect 12868 15206 12880 15258
rect 12880 15206 12894 15258
rect 12918 15206 12932 15258
rect 12932 15206 12944 15258
rect 12944 15206 12974 15258
rect 12998 15206 13008 15258
rect 13008 15206 13054 15258
rect 12758 15204 12814 15206
rect 12838 15204 12894 15206
rect 12918 15204 12974 15206
rect 12998 15204 13054 15206
rect 12098 14714 12154 14716
rect 12178 14714 12234 14716
rect 12258 14714 12314 14716
rect 12338 14714 12394 14716
rect 12098 14662 12144 14714
rect 12144 14662 12154 14714
rect 12178 14662 12208 14714
rect 12208 14662 12220 14714
rect 12220 14662 12234 14714
rect 12258 14662 12272 14714
rect 12272 14662 12284 14714
rect 12284 14662 12314 14714
rect 12338 14662 12348 14714
rect 12348 14662 12394 14714
rect 12098 14660 12154 14662
rect 12178 14660 12234 14662
rect 12258 14660 12314 14662
rect 12338 14660 12394 14662
rect 11058 12688 11114 12744
rect 5330 7642 5386 7644
rect 5410 7642 5466 7644
rect 5490 7642 5546 7644
rect 5570 7642 5626 7644
rect 5330 7590 5376 7642
rect 5376 7590 5386 7642
rect 5410 7590 5440 7642
rect 5440 7590 5452 7642
rect 5452 7590 5466 7642
rect 5490 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5546 7642
rect 5570 7590 5580 7642
rect 5580 7590 5626 7642
rect 5330 7588 5386 7590
rect 5410 7588 5466 7590
rect 5490 7588 5546 7590
rect 5570 7588 5626 7590
rect 4670 7098 4726 7100
rect 4750 7098 4806 7100
rect 4830 7098 4886 7100
rect 4910 7098 4966 7100
rect 4670 7046 4716 7098
rect 4716 7046 4726 7098
rect 4750 7046 4780 7098
rect 4780 7046 4792 7098
rect 4792 7046 4806 7098
rect 4830 7046 4844 7098
rect 4844 7046 4856 7098
rect 4856 7046 4886 7098
rect 4910 7046 4920 7098
rect 4920 7046 4966 7098
rect 4670 7044 4726 7046
rect 4750 7044 4806 7046
rect 4830 7044 4886 7046
rect 4910 7044 4966 7046
rect 1398 6840 1454 6896
rect 9494 8744 9550 8800
rect 5330 6554 5386 6556
rect 5410 6554 5466 6556
rect 5490 6554 5546 6556
rect 5570 6554 5626 6556
rect 5330 6502 5376 6554
rect 5376 6502 5386 6554
rect 5410 6502 5440 6554
rect 5440 6502 5452 6554
rect 5452 6502 5466 6554
rect 5490 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5546 6554
rect 5570 6502 5580 6554
rect 5580 6502 5626 6554
rect 5330 6500 5386 6502
rect 5410 6500 5466 6502
rect 5490 6500 5546 6502
rect 5570 6500 5626 6502
rect 4670 6010 4726 6012
rect 4750 6010 4806 6012
rect 4830 6010 4886 6012
rect 4910 6010 4966 6012
rect 4670 5958 4716 6010
rect 4716 5958 4726 6010
rect 4750 5958 4780 6010
rect 4780 5958 4792 6010
rect 4792 5958 4806 6010
rect 4830 5958 4844 6010
rect 4844 5958 4856 6010
rect 4856 5958 4886 6010
rect 4910 5958 4920 6010
rect 4920 5958 4966 6010
rect 4670 5956 4726 5958
rect 4750 5956 4806 5958
rect 4830 5956 4886 5958
rect 4910 5956 4966 5958
rect 5330 5466 5386 5468
rect 5410 5466 5466 5468
rect 5490 5466 5546 5468
rect 5570 5466 5626 5468
rect 5330 5414 5376 5466
rect 5376 5414 5386 5466
rect 5410 5414 5440 5466
rect 5440 5414 5452 5466
rect 5452 5414 5466 5466
rect 5490 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5546 5466
rect 5570 5414 5580 5466
rect 5580 5414 5626 5466
rect 5330 5412 5386 5414
rect 5410 5412 5466 5414
rect 5490 5412 5546 5414
rect 5570 5412 5626 5414
rect 4670 4922 4726 4924
rect 4750 4922 4806 4924
rect 4830 4922 4886 4924
rect 4910 4922 4966 4924
rect 4670 4870 4716 4922
rect 4716 4870 4726 4922
rect 4750 4870 4780 4922
rect 4780 4870 4792 4922
rect 4792 4870 4806 4922
rect 4830 4870 4844 4922
rect 4844 4870 4856 4922
rect 4856 4870 4886 4922
rect 4910 4870 4920 4922
rect 4920 4870 4966 4922
rect 4670 4868 4726 4870
rect 4750 4868 4806 4870
rect 4830 4868 4886 4870
rect 4910 4868 4966 4870
rect 5330 4378 5386 4380
rect 5410 4378 5466 4380
rect 5490 4378 5546 4380
rect 5570 4378 5626 4380
rect 5330 4326 5376 4378
rect 5376 4326 5386 4378
rect 5410 4326 5440 4378
rect 5440 4326 5452 4378
rect 5452 4326 5466 4378
rect 5490 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5546 4378
rect 5570 4326 5580 4378
rect 5580 4326 5626 4378
rect 5330 4324 5386 4326
rect 5410 4324 5466 4326
rect 5490 4324 5546 4326
rect 5570 4324 5626 4326
rect 4670 3834 4726 3836
rect 4750 3834 4806 3836
rect 4830 3834 4886 3836
rect 4910 3834 4966 3836
rect 4670 3782 4716 3834
rect 4716 3782 4726 3834
rect 4750 3782 4780 3834
rect 4780 3782 4792 3834
rect 4792 3782 4806 3834
rect 4830 3782 4844 3834
rect 4844 3782 4856 3834
rect 4856 3782 4886 3834
rect 4910 3782 4920 3834
rect 4920 3782 4966 3834
rect 4670 3780 4726 3782
rect 4750 3780 4806 3782
rect 4830 3780 4886 3782
rect 4910 3780 4966 3782
rect 5330 3290 5386 3292
rect 5410 3290 5466 3292
rect 5490 3290 5546 3292
rect 5570 3290 5626 3292
rect 5330 3238 5376 3290
rect 5376 3238 5386 3290
rect 5410 3238 5440 3290
rect 5440 3238 5452 3290
rect 5452 3238 5466 3290
rect 5490 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5546 3290
rect 5570 3238 5580 3290
rect 5580 3238 5626 3290
rect 5330 3236 5386 3238
rect 5410 3236 5466 3238
rect 5490 3236 5546 3238
rect 5570 3236 5626 3238
rect 4670 2746 4726 2748
rect 4750 2746 4806 2748
rect 4830 2746 4886 2748
rect 4910 2746 4966 2748
rect 4670 2694 4716 2746
rect 4716 2694 4726 2746
rect 4750 2694 4780 2746
rect 4780 2694 4792 2746
rect 4792 2694 4806 2746
rect 4830 2694 4844 2746
rect 4844 2694 4856 2746
rect 4856 2694 4886 2746
rect 4910 2694 4920 2746
rect 4920 2694 4966 2746
rect 4670 2692 4726 2694
rect 4750 2692 4806 2694
rect 4830 2692 4886 2694
rect 4910 2692 4966 2694
rect 12098 13626 12154 13628
rect 12178 13626 12234 13628
rect 12258 13626 12314 13628
rect 12338 13626 12394 13628
rect 12098 13574 12144 13626
rect 12144 13574 12154 13626
rect 12178 13574 12208 13626
rect 12208 13574 12220 13626
rect 12220 13574 12234 13626
rect 12258 13574 12272 13626
rect 12272 13574 12284 13626
rect 12284 13574 12314 13626
rect 12338 13574 12348 13626
rect 12348 13574 12394 13626
rect 12098 13572 12154 13574
rect 12178 13572 12234 13574
rect 12258 13572 12314 13574
rect 12338 13572 12394 13574
rect 12098 12538 12154 12540
rect 12178 12538 12234 12540
rect 12258 12538 12314 12540
rect 12338 12538 12394 12540
rect 12098 12486 12144 12538
rect 12144 12486 12154 12538
rect 12178 12486 12208 12538
rect 12208 12486 12220 12538
rect 12220 12486 12234 12538
rect 12258 12486 12272 12538
rect 12272 12486 12284 12538
rect 12284 12486 12314 12538
rect 12338 12486 12348 12538
rect 12348 12486 12394 12538
rect 12098 12484 12154 12486
rect 12178 12484 12234 12486
rect 12258 12484 12314 12486
rect 12338 12484 12394 12486
rect 12758 14170 12814 14172
rect 12838 14170 12894 14172
rect 12918 14170 12974 14172
rect 12998 14170 13054 14172
rect 12758 14118 12804 14170
rect 12804 14118 12814 14170
rect 12838 14118 12868 14170
rect 12868 14118 12880 14170
rect 12880 14118 12894 14170
rect 12918 14118 12932 14170
rect 12932 14118 12944 14170
rect 12944 14118 12974 14170
rect 12998 14118 13008 14170
rect 13008 14118 13054 14170
rect 12758 14116 12814 14118
rect 12838 14116 12894 14118
rect 12918 14116 12974 14118
rect 12998 14116 13054 14118
rect 12758 13082 12814 13084
rect 12838 13082 12894 13084
rect 12918 13082 12974 13084
rect 12998 13082 13054 13084
rect 12758 13030 12804 13082
rect 12804 13030 12814 13082
rect 12838 13030 12868 13082
rect 12868 13030 12880 13082
rect 12880 13030 12894 13082
rect 12918 13030 12932 13082
rect 12932 13030 12944 13082
rect 12944 13030 12974 13082
rect 12998 13030 13008 13082
rect 13008 13030 13054 13082
rect 12758 13028 12814 13030
rect 12838 13028 12894 13030
rect 12918 13028 12974 13030
rect 12998 13028 13054 13030
rect 12098 11450 12154 11452
rect 12178 11450 12234 11452
rect 12258 11450 12314 11452
rect 12338 11450 12394 11452
rect 12098 11398 12144 11450
rect 12144 11398 12154 11450
rect 12178 11398 12208 11450
rect 12208 11398 12220 11450
rect 12220 11398 12234 11450
rect 12258 11398 12272 11450
rect 12272 11398 12284 11450
rect 12284 11398 12314 11450
rect 12338 11398 12348 11450
rect 12348 11398 12394 11450
rect 12098 11396 12154 11398
rect 12178 11396 12234 11398
rect 12258 11396 12314 11398
rect 12338 11396 12394 11398
rect 12098 10362 12154 10364
rect 12178 10362 12234 10364
rect 12258 10362 12314 10364
rect 12338 10362 12394 10364
rect 12098 10310 12144 10362
rect 12144 10310 12154 10362
rect 12178 10310 12208 10362
rect 12208 10310 12220 10362
rect 12220 10310 12234 10362
rect 12258 10310 12272 10362
rect 12272 10310 12284 10362
rect 12284 10310 12314 10362
rect 12338 10310 12348 10362
rect 12348 10310 12394 10362
rect 12098 10308 12154 10310
rect 12178 10308 12234 10310
rect 12258 10308 12314 10310
rect 12338 10308 12394 10310
rect 12098 9274 12154 9276
rect 12178 9274 12234 9276
rect 12258 9274 12314 9276
rect 12338 9274 12394 9276
rect 12098 9222 12144 9274
rect 12144 9222 12154 9274
rect 12178 9222 12208 9274
rect 12208 9222 12220 9274
rect 12220 9222 12234 9274
rect 12258 9222 12272 9274
rect 12272 9222 12284 9274
rect 12284 9222 12314 9274
rect 12338 9222 12348 9274
rect 12348 9222 12394 9274
rect 12098 9220 12154 9222
rect 12178 9220 12234 9222
rect 12258 9220 12314 9222
rect 12338 9220 12394 9222
rect 12098 8186 12154 8188
rect 12178 8186 12234 8188
rect 12258 8186 12314 8188
rect 12338 8186 12394 8188
rect 12098 8134 12144 8186
rect 12144 8134 12154 8186
rect 12178 8134 12208 8186
rect 12208 8134 12220 8186
rect 12220 8134 12234 8186
rect 12258 8134 12272 8186
rect 12272 8134 12284 8186
rect 12284 8134 12314 8186
rect 12338 8134 12348 8186
rect 12348 8134 12394 8186
rect 12098 8132 12154 8134
rect 12178 8132 12234 8134
rect 12258 8132 12314 8134
rect 12338 8132 12394 8134
rect 12758 11994 12814 11996
rect 12838 11994 12894 11996
rect 12918 11994 12974 11996
rect 12998 11994 13054 11996
rect 12758 11942 12804 11994
rect 12804 11942 12814 11994
rect 12838 11942 12868 11994
rect 12868 11942 12880 11994
rect 12880 11942 12894 11994
rect 12918 11942 12932 11994
rect 12932 11942 12944 11994
rect 12944 11942 12974 11994
rect 12998 11942 13008 11994
rect 13008 11942 13054 11994
rect 12758 11940 12814 11942
rect 12838 11940 12894 11942
rect 12918 11940 12974 11942
rect 12998 11940 13054 11942
rect 14278 16516 14334 16552
rect 14278 16496 14280 16516
rect 14280 16496 14332 16516
rect 14332 16496 14334 16516
rect 12758 10906 12814 10908
rect 12838 10906 12894 10908
rect 12918 10906 12974 10908
rect 12998 10906 13054 10908
rect 12758 10854 12804 10906
rect 12804 10854 12814 10906
rect 12838 10854 12868 10906
rect 12868 10854 12880 10906
rect 12880 10854 12894 10906
rect 12918 10854 12932 10906
rect 12932 10854 12944 10906
rect 12944 10854 12974 10906
rect 12998 10854 13008 10906
rect 13008 10854 13054 10906
rect 12758 10852 12814 10854
rect 12838 10852 12894 10854
rect 12918 10852 12974 10854
rect 12998 10852 13054 10854
rect 12758 9818 12814 9820
rect 12838 9818 12894 9820
rect 12918 9818 12974 9820
rect 12998 9818 13054 9820
rect 12758 9766 12804 9818
rect 12804 9766 12814 9818
rect 12838 9766 12868 9818
rect 12868 9766 12880 9818
rect 12880 9766 12894 9818
rect 12918 9766 12932 9818
rect 12932 9766 12944 9818
rect 12944 9766 12974 9818
rect 12998 9766 13008 9818
rect 13008 9766 13054 9818
rect 12758 9764 12814 9766
rect 12838 9764 12894 9766
rect 12918 9764 12974 9766
rect 12998 9764 13054 9766
rect 12758 8730 12814 8732
rect 12838 8730 12894 8732
rect 12918 8730 12974 8732
rect 12998 8730 13054 8732
rect 12758 8678 12804 8730
rect 12804 8678 12814 8730
rect 12838 8678 12868 8730
rect 12868 8678 12880 8730
rect 12880 8678 12894 8730
rect 12918 8678 12932 8730
rect 12932 8678 12944 8730
rect 12944 8678 12974 8730
rect 12998 8678 13008 8730
rect 13008 8678 13054 8730
rect 12758 8676 12814 8678
rect 12838 8676 12894 8678
rect 12918 8676 12974 8678
rect 12998 8676 13054 8678
rect 12758 7642 12814 7644
rect 12838 7642 12894 7644
rect 12918 7642 12974 7644
rect 12998 7642 13054 7644
rect 12758 7590 12804 7642
rect 12804 7590 12814 7642
rect 12838 7590 12868 7642
rect 12868 7590 12880 7642
rect 12880 7590 12894 7642
rect 12918 7590 12932 7642
rect 12932 7590 12944 7642
rect 12944 7590 12974 7642
rect 12998 7590 13008 7642
rect 13008 7590 13054 7642
rect 12758 7588 12814 7590
rect 12838 7588 12894 7590
rect 12918 7588 12974 7590
rect 12998 7588 13054 7590
rect 12098 7098 12154 7100
rect 12178 7098 12234 7100
rect 12258 7098 12314 7100
rect 12338 7098 12394 7100
rect 12098 7046 12144 7098
rect 12144 7046 12154 7098
rect 12178 7046 12208 7098
rect 12208 7046 12220 7098
rect 12220 7046 12234 7098
rect 12258 7046 12272 7098
rect 12272 7046 12284 7098
rect 12284 7046 12314 7098
rect 12338 7046 12348 7098
rect 12348 7046 12394 7098
rect 12098 7044 12154 7046
rect 12178 7044 12234 7046
rect 12258 7044 12314 7046
rect 12338 7044 12394 7046
rect 12098 6010 12154 6012
rect 12178 6010 12234 6012
rect 12258 6010 12314 6012
rect 12338 6010 12394 6012
rect 12098 5958 12144 6010
rect 12144 5958 12154 6010
rect 12178 5958 12208 6010
rect 12208 5958 12220 6010
rect 12220 5958 12234 6010
rect 12258 5958 12272 6010
rect 12272 5958 12284 6010
rect 12284 5958 12314 6010
rect 12338 5958 12348 6010
rect 12348 5958 12394 6010
rect 12098 5956 12154 5958
rect 12178 5956 12234 5958
rect 12258 5956 12314 5958
rect 12338 5956 12394 5958
rect 12098 4922 12154 4924
rect 12178 4922 12234 4924
rect 12258 4922 12314 4924
rect 12338 4922 12394 4924
rect 12098 4870 12144 4922
rect 12144 4870 12154 4922
rect 12178 4870 12208 4922
rect 12208 4870 12220 4922
rect 12220 4870 12234 4922
rect 12258 4870 12272 4922
rect 12272 4870 12284 4922
rect 12284 4870 12314 4922
rect 12338 4870 12348 4922
rect 12348 4870 12394 4922
rect 12098 4868 12154 4870
rect 12178 4868 12234 4870
rect 12258 4868 12314 4870
rect 12338 4868 12394 4870
rect 12098 3834 12154 3836
rect 12178 3834 12234 3836
rect 12258 3834 12314 3836
rect 12338 3834 12394 3836
rect 12098 3782 12144 3834
rect 12144 3782 12154 3834
rect 12178 3782 12208 3834
rect 12208 3782 12220 3834
rect 12220 3782 12234 3834
rect 12258 3782 12272 3834
rect 12272 3782 12284 3834
rect 12284 3782 12314 3834
rect 12338 3782 12348 3834
rect 12348 3782 12394 3834
rect 12098 3780 12154 3782
rect 12178 3780 12234 3782
rect 12258 3780 12314 3782
rect 12338 3780 12394 3782
rect 12098 2746 12154 2748
rect 12178 2746 12234 2748
rect 12258 2746 12314 2748
rect 12338 2746 12394 2748
rect 12098 2694 12144 2746
rect 12144 2694 12154 2746
rect 12178 2694 12208 2746
rect 12208 2694 12220 2746
rect 12220 2694 12234 2746
rect 12258 2694 12272 2746
rect 12272 2694 12284 2746
rect 12284 2694 12314 2746
rect 12338 2694 12348 2746
rect 12348 2694 12394 2746
rect 12098 2692 12154 2694
rect 12178 2692 12234 2694
rect 12258 2692 12314 2694
rect 12338 2692 12394 2694
rect 12758 6554 12814 6556
rect 12838 6554 12894 6556
rect 12918 6554 12974 6556
rect 12998 6554 13054 6556
rect 12758 6502 12804 6554
rect 12804 6502 12814 6554
rect 12838 6502 12868 6554
rect 12868 6502 12880 6554
rect 12880 6502 12894 6554
rect 12918 6502 12932 6554
rect 12932 6502 12944 6554
rect 12944 6502 12974 6554
rect 12998 6502 13008 6554
rect 13008 6502 13054 6554
rect 12758 6500 12814 6502
rect 12838 6500 12894 6502
rect 12918 6500 12974 6502
rect 12998 6500 13054 6502
rect 12758 5466 12814 5468
rect 12838 5466 12894 5468
rect 12918 5466 12974 5468
rect 12998 5466 13054 5468
rect 12758 5414 12804 5466
rect 12804 5414 12814 5466
rect 12838 5414 12868 5466
rect 12868 5414 12880 5466
rect 12880 5414 12894 5466
rect 12918 5414 12932 5466
rect 12932 5414 12944 5466
rect 12944 5414 12974 5466
rect 12998 5414 13008 5466
rect 13008 5414 13054 5466
rect 12758 5412 12814 5414
rect 12838 5412 12894 5414
rect 12918 5412 12974 5414
rect 12998 5412 13054 5414
rect 12758 4378 12814 4380
rect 12838 4378 12894 4380
rect 12918 4378 12974 4380
rect 12998 4378 13054 4380
rect 12758 4326 12804 4378
rect 12804 4326 12814 4378
rect 12838 4326 12868 4378
rect 12868 4326 12880 4378
rect 12880 4326 12894 4378
rect 12918 4326 12932 4378
rect 12932 4326 12944 4378
rect 12944 4326 12974 4378
rect 12998 4326 13008 4378
rect 13008 4326 13054 4378
rect 12758 4324 12814 4326
rect 12838 4324 12894 4326
rect 12918 4324 12974 4326
rect 12998 4324 13054 4326
rect 12758 3290 12814 3292
rect 12838 3290 12894 3292
rect 12918 3290 12974 3292
rect 12998 3290 13054 3292
rect 12758 3238 12804 3290
rect 12804 3238 12814 3290
rect 12838 3238 12868 3290
rect 12868 3238 12880 3290
rect 12880 3238 12894 3290
rect 12918 3238 12932 3290
rect 12932 3238 12944 3290
rect 12944 3238 12974 3290
rect 12998 3238 13008 3290
rect 13008 3238 13054 3290
rect 12758 3236 12814 3238
rect 12838 3236 12894 3238
rect 12918 3236 12974 3238
rect 12998 3236 13054 3238
rect 14922 12280 14978 12336
rect 17590 18264 17646 18320
rect 19526 28858 19582 28860
rect 19606 28858 19662 28860
rect 19686 28858 19742 28860
rect 19766 28858 19822 28860
rect 19526 28806 19572 28858
rect 19572 28806 19582 28858
rect 19606 28806 19636 28858
rect 19636 28806 19648 28858
rect 19648 28806 19662 28858
rect 19686 28806 19700 28858
rect 19700 28806 19712 28858
rect 19712 28806 19742 28858
rect 19766 28806 19776 28858
rect 19776 28806 19822 28858
rect 19526 28804 19582 28806
rect 19606 28804 19662 28806
rect 19686 28804 19742 28806
rect 19766 28804 19822 28806
rect 19526 27770 19582 27772
rect 19606 27770 19662 27772
rect 19686 27770 19742 27772
rect 19766 27770 19822 27772
rect 19526 27718 19572 27770
rect 19572 27718 19582 27770
rect 19606 27718 19636 27770
rect 19636 27718 19648 27770
rect 19648 27718 19662 27770
rect 19686 27718 19700 27770
rect 19700 27718 19712 27770
rect 19712 27718 19742 27770
rect 19766 27718 19776 27770
rect 19776 27718 19822 27770
rect 19526 27716 19582 27718
rect 19606 27716 19662 27718
rect 19686 27716 19742 27718
rect 19766 27716 19822 27718
rect 19526 26682 19582 26684
rect 19606 26682 19662 26684
rect 19686 26682 19742 26684
rect 19766 26682 19822 26684
rect 19526 26630 19572 26682
rect 19572 26630 19582 26682
rect 19606 26630 19636 26682
rect 19636 26630 19648 26682
rect 19648 26630 19662 26682
rect 19686 26630 19700 26682
rect 19700 26630 19712 26682
rect 19712 26630 19742 26682
rect 19766 26630 19776 26682
rect 19776 26630 19822 26682
rect 19526 26628 19582 26630
rect 19606 26628 19662 26630
rect 19686 26628 19742 26630
rect 19766 26628 19822 26630
rect 19526 25594 19582 25596
rect 19606 25594 19662 25596
rect 19686 25594 19742 25596
rect 19766 25594 19822 25596
rect 19526 25542 19572 25594
rect 19572 25542 19582 25594
rect 19606 25542 19636 25594
rect 19636 25542 19648 25594
rect 19648 25542 19662 25594
rect 19686 25542 19700 25594
rect 19700 25542 19712 25594
rect 19712 25542 19742 25594
rect 19766 25542 19776 25594
rect 19776 25542 19822 25594
rect 19526 25540 19582 25542
rect 19606 25540 19662 25542
rect 19686 25540 19742 25542
rect 19766 25540 19822 25542
rect 19526 24506 19582 24508
rect 19606 24506 19662 24508
rect 19686 24506 19742 24508
rect 19766 24506 19822 24508
rect 19526 24454 19572 24506
rect 19572 24454 19582 24506
rect 19606 24454 19636 24506
rect 19636 24454 19648 24506
rect 19648 24454 19662 24506
rect 19686 24454 19700 24506
rect 19700 24454 19712 24506
rect 19712 24454 19742 24506
rect 19766 24454 19776 24506
rect 19776 24454 19822 24506
rect 19526 24452 19582 24454
rect 19606 24452 19662 24454
rect 19686 24452 19742 24454
rect 19766 24452 19822 24454
rect 19526 23418 19582 23420
rect 19606 23418 19662 23420
rect 19686 23418 19742 23420
rect 19766 23418 19822 23420
rect 19526 23366 19572 23418
rect 19572 23366 19582 23418
rect 19606 23366 19636 23418
rect 19636 23366 19648 23418
rect 19648 23366 19662 23418
rect 19686 23366 19700 23418
rect 19700 23366 19712 23418
rect 19712 23366 19742 23418
rect 19766 23366 19776 23418
rect 19776 23366 19822 23418
rect 19526 23364 19582 23366
rect 19606 23364 19662 23366
rect 19686 23364 19742 23366
rect 19766 23364 19822 23366
rect 19526 22330 19582 22332
rect 19606 22330 19662 22332
rect 19686 22330 19742 22332
rect 19766 22330 19822 22332
rect 19526 22278 19572 22330
rect 19572 22278 19582 22330
rect 19606 22278 19636 22330
rect 19636 22278 19648 22330
rect 19648 22278 19662 22330
rect 19686 22278 19700 22330
rect 19700 22278 19712 22330
rect 19712 22278 19742 22330
rect 19766 22278 19776 22330
rect 19776 22278 19822 22330
rect 19526 22276 19582 22278
rect 19606 22276 19662 22278
rect 19686 22276 19742 22278
rect 19766 22276 19822 22278
rect 20186 28314 20242 28316
rect 20266 28314 20322 28316
rect 20346 28314 20402 28316
rect 20426 28314 20482 28316
rect 20186 28262 20232 28314
rect 20232 28262 20242 28314
rect 20266 28262 20296 28314
rect 20296 28262 20308 28314
rect 20308 28262 20322 28314
rect 20346 28262 20360 28314
rect 20360 28262 20372 28314
rect 20372 28262 20402 28314
rect 20426 28262 20436 28314
rect 20436 28262 20482 28314
rect 20186 28260 20242 28262
rect 20266 28260 20322 28262
rect 20346 28260 20402 28262
rect 20426 28260 20482 28262
rect 20186 27226 20242 27228
rect 20266 27226 20322 27228
rect 20346 27226 20402 27228
rect 20426 27226 20482 27228
rect 20186 27174 20232 27226
rect 20232 27174 20242 27226
rect 20266 27174 20296 27226
rect 20296 27174 20308 27226
rect 20308 27174 20322 27226
rect 20346 27174 20360 27226
rect 20360 27174 20372 27226
rect 20372 27174 20402 27226
rect 20426 27174 20436 27226
rect 20436 27174 20482 27226
rect 20186 27172 20242 27174
rect 20266 27172 20322 27174
rect 20346 27172 20402 27174
rect 20426 27172 20482 27174
rect 20186 26138 20242 26140
rect 20266 26138 20322 26140
rect 20346 26138 20402 26140
rect 20426 26138 20482 26140
rect 20186 26086 20232 26138
rect 20232 26086 20242 26138
rect 20266 26086 20296 26138
rect 20296 26086 20308 26138
rect 20308 26086 20322 26138
rect 20346 26086 20360 26138
rect 20360 26086 20372 26138
rect 20372 26086 20402 26138
rect 20426 26086 20436 26138
rect 20436 26086 20482 26138
rect 20186 26084 20242 26086
rect 20266 26084 20322 26086
rect 20346 26084 20402 26086
rect 20426 26084 20482 26086
rect 20186 25050 20242 25052
rect 20266 25050 20322 25052
rect 20346 25050 20402 25052
rect 20426 25050 20482 25052
rect 20186 24998 20232 25050
rect 20232 24998 20242 25050
rect 20266 24998 20296 25050
rect 20296 24998 20308 25050
rect 20308 24998 20322 25050
rect 20346 24998 20360 25050
rect 20360 24998 20372 25050
rect 20372 24998 20402 25050
rect 20426 24998 20436 25050
rect 20436 24998 20482 25050
rect 20186 24996 20242 24998
rect 20266 24996 20322 24998
rect 20346 24996 20402 24998
rect 20426 24996 20482 24998
rect 20186 23962 20242 23964
rect 20266 23962 20322 23964
rect 20346 23962 20402 23964
rect 20426 23962 20482 23964
rect 20186 23910 20232 23962
rect 20232 23910 20242 23962
rect 20266 23910 20296 23962
rect 20296 23910 20308 23962
rect 20308 23910 20322 23962
rect 20346 23910 20360 23962
rect 20360 23910 20372 23962
rect 20372 23910 20402 23962
rect 20426 23910 20436 23962
rect 20436 23910 20482 23962
rect 20186 23908 20242 23910
rect 20266 23908 20322 23910
rect 20346 23908 20402 23910
rect 20426 23908 20482 23910
rect 20186 22874 20242 22876
rect 20266 22874 20322 22876
rect 20346 22874 20402 22876
rect 20426 22874 20482 22876
rect 20186 22822 20232 22874
rect 20232 22822 20242 22874
rect 20266 22822 20296 22874
rect 20296 22822 20308 22874
rect 20308 22822 20322 22874
rect 20346 22822 20360 22874
rect 20360 22822 20372 22874
rect 20372 22822 20402 22874
rect 20426 22822 20436 22874
rect 20436 22822 20482 22874
rect 20186 22820 20242 22822
rect 20266 22820 20322 22822
rect 20346 22820 20402 22822
rect 20426 22820 20482 22822
rect 20186 21786 20242 21788
rect 20266 21786 20322 21788
rect 20346 21786 20402 21788
rect 20426 21786 20482 21788
rect 20186 21734 20232 21786
rect 20232 21734 20242 21786
rect 20266 21734 20296 21786
rect 20296 21734 20308 21786
rect 20308 21734 20322 21786
rect 20346 21734 20360 21786
rect 20360 21734 20372 21786
rect 20372 21734 20402 21786
rect 20426 21734 20436 21786
rect 20436 21734 20482 21786
rect 20186 21732 20242 21734
rect 20266 21732 20322 21734
rect 20346 21732 20402 21734
rect 20426 21732 20482 21734
rect 19526 21242 19582 21244
rect 19606 21242 19662 21244
rect 19686 21242 19742 21244
rect 19766 21242 19822 21244
rect 19526 21190 19572 21242
rect 19572 21190 19582 21242
rect 19606 21190 19636 21242
rect 19636 21190 19648 21242
rect 19648 21190 19662 21242
rect 19686 21190 19700 21242
rect 19700 21190 19712 21242
rect 19712 21190 19742 21242
rect 19766 21190 19776 21242
rect 19776 21190 19822 21242
rect 19526 21188 19582 21190
rect 19606 21188 19662 21190
rect 19686 21188 19742 21190
rect 19766 21188 19822 21190
rect 19526 20154 19582 20156
rect 19606 20154 19662 20156
rect 19686 20154 19742 20156
rect 19766 20154 19822 20156
rect 19526 20102 19572 20154
rect 19572 20102 19582 20154
rect 19606 20102 19636 20154
rect 19636 20102 19648 20154
rect 19648 20102 19662 20154
rect 19686 20102 19700 20154
rect 19700 20102 19712 20154
rect 19712 20102 19742 20154
rect 19766 20102 19776 20154
rect 19776 20102 19822 20154
rect 19526 20100 19582 20102
rect 19606 20100 19662 20102
rect 19686 20100 19742 20102
rect 19766 20100 19822 20102
rect 19526 19066 19582 19068
rect 19606 19066 19662 19068
rect 19686 19066 19742 19068
rect 19766 19066 19822 19068
rect 19526 19014 19572 19066
rect 19572 19014 19582 19066
rect 19606 19014 19636 19066
rect 19636 19014 19648 19066
rect 19648 19014 19662 19066
rect 19686 19014 19700 19066
rect 19700 19014 19712 19066
rect 19712 19014 19742 19066
rect 19766 19014 19776 19066
rect 19776 19014 19822 19066
rect 19526 19012 19582 19014
rect 19606 19012 19662 19014
rect 19686 19012 19742 19014
rect 19766 19012 19822 19014
rect 20186 20698 20242 20700
rect 20266 20698 20322 20700
rect 20346 20698 20402 20700
rect 20426 20698 20482 20700
rect 20186 20646 20232 20698
rect 20232 20646 20242 20698
rect 20266 20646 20296 20698
rect 20296 20646 20308 20698
rect 20308 20646 20322 20698
rect 20346 20646 20360 20698
rect 20360 20646 20372 20698
rect 20372 20646 20402 20698
rect 20426 20646 20436 20698
rect 20436 20646 20482 20698
rect 20186 20644 20242 20646
rect 20266 20644 20322 20646
rect 20346 20644 20402 20646
rect 20426 20644 20482 20646
rect 20994 22636 21050 22672
rect 20994 22616 20996 22636
rect 20996 22616 21048 22636
rect 21048 22616 21050 22636
rect 26954 28858 27010 28860
rect 27034 28858 27090 28860
rect 27114 28858 27170 28860
rect 27194 28858 27250 28860
rect 26954 28806 27000 28858
rect 27000 28806 27010 28858
rect 27034 28806 27064 28858
rect 27064 28806 27076 28858
rect 27076 28806 27090 28858
rect 27114 28806 27128 28858
rect 27128 28806 27140 28858
rect 27140 28806 27170 28858
rect 27194 28806 27204 28858
rect 27204 28806 27250 28858
rect 26954 28804 27010 28806
rect 27034 28804 27090 28806
rect 27114 28804 27170 28806
rect 27194 28804 27250 28806
rect 27614 28314 27670 28316
rect 27694 28314 27750 28316
rect 27774 28314 27830 28316
rect 27854 28314 27910 28316
rect 27614 28262 27660 28314
rect 27660 28262 27670 28314
rect 27694 28262 27724 28314
rect 27724 28262 27736 28314
rect 27736 28262 27750 28314
rect 27774 28262 27788 28314
rect 27788 28262 27800 28314
rect 27800 28262 27830 28314
rect 27854 28262 27864 28314
rect 27864 28262 27910 28314
rect 27614 28260 27670 28262
rect 27694 28260 27750 28262
rect 27774 28260 27830 28262
rect 27854 28260 27910 28262
rect 26954 27770 27010 27772
rect 27034 27770 27090 27772
rect 27114 27770 27170 27772
rect 27194 27770 27250 27772
rect 26954 27718 27000 27770
rect 27000 27718 27010 27770
rect 27034 27718 27064 27770
rect 27064 27718 27076 27770
rect 27076 27718 27090 27770
rect 27114 27718 27128 27770
rect 27128 27718 27140 27770
rect 27140 27718 27170 27770
rect 27194 27718 27204 27770
rect 27204 27718 27250 27770
rect 26954 27716 27010 27718
rect 27034 27716 27090 27718
rect 27114 27716 27170 27718
rect 27194 27716 27250 27718
rect 27614 27226 27670 27228
rect 27694 27226 27750 27228
rect 27774 27226 27830 27228
rect 27854 27226 27910 27228
rect 27614 27174 27660 27226
rect 27660 27174 27670 27226
rect 27694 27174 27724 27226
rect 27724 27174 27736 27226
rect 27736 27174 27750 27226
rect 27774 27174 27788 27226
rect 27788 27174 27800 27226
rect 27800 27174 27830 27226
rect 27854 27174 27864 27226
rect 27864 27174 27910 27226
rect 27614 27172 27670 27174
rect 27694 27172 27750 27174
rect 27774 27172 27830 27174
rect 27854 27172 27910 27174
rect 26954 26682 27010 26684
rect 27034 26682 27090 26684
rect 27114 26682 27170 26684
rect 27194 26682 27250 26684
rect 26954 26630 27000 26682
rect 27000 26630 27010 26682
rect 27034 26630 27064 26682
rect 27064 26630 27076 26682
rect 27076 26630 27090 26682
rect 27114 26630 27128 26682
rect 27128 26630 27140 26682
rect 27140 26630 27170 26682
rect 27194 26630 27204 26682
rect 27204 26630 27250 26682
rect 26954 26628 27010 26630
rect 27034 26628 27090 26630
rect 27114 26628 27170 26630
rect 27194 26628 27250 26630
rect 27614 26138 27670 26140
rect 27694 26138 27750 26140
rect 27774 26138 27830 26140
rect 27854 26138 27910 26140
rect 27614 26086 27660 26138
rect 27660 26086 27670 26138
rect 27694 26086 27724 26138
rect 27724 26086 27736 26138
rect 27736 26086 27750 26138
rect 27774 26086 27788 26138
rect 27788 26086 27800 26138
rect 27800 26086 27830 26138
rect 27854 26086 27864 26138
rect 27864 26086 27910 26138
rect 27614 26084 27670 26086
rect 27694 26084 27750 26086
rect 27774 26084 27830 26086
rect 27854 26084 27910 26086
rect 26954 25594 27010 25596
rect 27034 25594 27090 25596
rect 27114 25594 27170 25596
rect 27194 25594 27250 25596
rect 26954 25542 27000 25594
rect 27000 25542 27010 25594
rect 27034 25542 27064 25594
rect 27064 25542 27076 25594
rect 27076 25542 27090 25594
rect 27114 25542 27128 25594
rect 27128 25542 27140 25594
rect 27140 25542 27170 25594
rect 27194 25542 27204 25594
rect 27204 25542 27250 25594
rect 26954 25540 27010 25542
rect 27034 25540 27090 25542
rect 27114 25540 27170 25542
rect 27194 25540 27250 25542
rect 22006 22516 22008 22536
rect 22008 22516 22060 22536
rect 22060 22516 22062 22536
rect 22006 22480 22062 22516
rect 22558 22636 22614 22672
rect 22558 22616 22560 22636
rect 22560 22616 22612 22636
rect 22612 22616 22614 22636
rect 20186 19610 20242 19612
rect 20266 19610 20322 19612
rect 20346 19610 20402 19612
rect 20426 19610 20482 19612
rect 20186 19558 20232 19610
rect 20232 19558 20242 19610
rect 20266 19558 20296 19610
rect 20296 19558 20308 19610
rect 20308 19558 20322 19610
rect 20346 19558 20360 19610
rect 20360 19558 20372 19610
rect 20372 19558 20402 19610
rect 20426 19558 20436 19610
rect 20436 19558 20482 19610
rect 20186 19556 20242 19558
rect 20266 19556 20322 19558
rect 20346 19556 20402 19558
rect 20426 19556 20482 19558
rect 20186 18522 20242 18524
rect 20266 18522 20322 18524
rect 20346 18522 20402 18524
rect 20426 18522 20482 18524
rect 20186 18470 20232 18522
rect 20232 18470 20242 18522
rect 20266 18470 20296 18522
rect 20296 18470 20308 18522
rect 20308 18470 20322 18522
rect 20346 18470 20360 18522
rect 20360 18470 20372 18522
rect 20372 18470 20402 18522
rect 20426 18470 20436 18522
rect 20436 18470 20482 18522
rect 20186 18468 20242 18470
rect 20266 18468 20322 18470
rect 20346 18468 20402 18470
rect 20426 18468 20482 18470
rect 19526 17978 19582 17980
rect 19606 17978 19662 17980
rect 19686 17978 19742 17980
rect 19766 17978 19822 17980
rect 19526 17926 19572 17978
rect 19572 17926 19582 17978
rect 19606 17926 19636 17978
rect 19636 17926 19648 17978
rect 19648 17926 19662 17978
rect 19686 17926 19700 17978
rect 19700 17926 19712 17978
rect 19712 17926 19742 17978
rect 19766 17926 19776 17978
rect 19776 17926 19822 17978
rect 19526 17924 19582 17926
rect 19606 17924 19662 17926
rect 19686 17924 19742 17926
rect 19766 17924 19822 17926
rect 16486 14320 16542 14376
rect 16302 12688 16358 12744
rect 19526 16890 19582 16892
rect 19606 16890 19662 16892
rect 19686 16890 19742 16892
rect 19766 16890 19822 16892
rect 19526 16838 19572 16890
rect 19572 16838 19582 16890
rect 19606 16838 19636 16890
rect 19636 16838 19648 16890
rect 19648 16838 19662 16890
rect 19686 16838 19700 16890
rect 19700 16838 19712 16890
rect 19712 16838 19742 16890
rect 19766 16838 19776 16890
rect 19776 16838 19822 16890
rect 19526 16836 19582 16838
rect 19606 16836 19662 16838
rect 19686 16836 19742 16838
rect 19766 16836 19822 16838
rect 20186 17434 20242 17436
rect 20266 17434 20322 17436
rect 20346 17434 20402 17436
rect 20426 17434 20482 17436
rect 20186 17382 20232 17434
rect 20232 17382 20242 17434
rect 20266 17382 20296 17434
rect 20296 17382 20308 17434
rect 20308 17382 20322 17434
rect 20346 17382 20360 17434
rect 20360 17382 20372 17434
rect 20372 17382 20402 17434
rect 20426 17382 20436 17434
rect 20436 17382 20482 17434
rect 20186 17380 20242 17382
rect 20266 17380 20322 17382
rect 20346 17380 20402 17382
rect 20426 17380 20482 17382
rect 20186 16346 20242 16348
rect 20266 16346 20322 16348
rect 20346 16346 20402 16348
rect 20426 16346 20482 16348
rect 20186 16294 20232 16346
rect 20232 16294 20242 16346
rect 20266 16294 20296 16346
rect 20296 16294 20308 16346
rect 20308 16294 20322 16346
rect 20346 16294 20360 16346
rect 20360 16294 20372 16346
rect 20372 16294 20402 16346
rect 20426 16294 20436 16346
rect 20436 16294 20482 16346
rect 20186 16292 20242 16294
rect 20266 16292 20322 16294
rect 20346 16292 20402 16294
rect 20426 16292 20482 16294
rect 27614 25050 27670 25052
rect 27694 25050 27750 25052
rect 27774 25050 27830 25052
rect 27854 25050 27910 25052
rect 27614 24998 27660 25050
rect 27660 24998 27670 25050
rect 27694 24998 27724 25050
rect 27724 24998 27736 25050
rect 27736 24998 27750 25050
rect 27774 24998 27788 25050
rect 27788 24998 27800 25050
rect 27800 24998 27830 25050
rect 27854 24998 27864 25050
rect 27864 24998 27910 25050
rect 27614 24996 27670 24998
rect 27694 24996 27750 24998
rect 27774 24996 27830 24998
rect 27854 24996 27910 24998
rect 24030 22480 24086 22536
rect 26954 24506 27010 24508
rect 27034 24506 27090 24508
rect 27114 24506 27170 24508
rect 27194 24506 27250 24508
rect 26954 24454 27000 24506
rect 27000 24454 27010 24506
rect 27034 24454 27064 24506
rect 27064 24454 27076 24506
rect 27076 24454 27090 24506
rect 27114 24454 27128 24506
rect 27128 24454 27140 24506
rect 27140 24454 27170 24506
rect 27194 24454 27204 24506
rect 27204 24454 27250 24506
rect 26954 24452 27010 24454
rect 27034 24452 27090 24454
rect 27114 24452 27170 24454
rect 27194 24452 27250 24454
rect 27614 23962 27670 23964
rect 27694 23962 27750 23964
rect 27774 23962 27830 23964
rect 27854 23962 27910 23964
rect 27614 23910 27660 23962
rect 27660 23910 27670 23962
rect 27694 23910 27724 23962
rect 27724 23910 27736 23962
rect 27736 23910 27750 23962
rect 27774 23910 27788 23962
rect 27788 23910 27800 23962
rect 27800 23910 27830 23962
rect 27854 23910 27864 23962
rect 27864 23910 27910 23962
rect 27614 23908 27670 23910
rect 27694 23908 27750 23910
rect 27774 23908 27830 23910
rect 27854 23908 27910 23910
rect 20810 16532 20812 16552
rect 20812 16532 20864 16552
rect 20864 16532 20866 16552
rect 20810 16496 20866 16532
rect 19526 15802 19582 15804
rect 19606 15802 19662 15804
rect 19686 15802 19742 15804
rect 19766 15802 19822 15804
rect 19526 15750 19572 15802
rect 19572 15750 19582 15802
rect 19606 15750 19636 15802
rect 19636 15750 19648 15802
rect 19648 15750 19662 15802
rect 19686 15750 19700 15802
rect 19700 15750 19712 15802
rect 19712 15750 19742 15802
rect 19766 15750 19776 15802
rect 19776 15750 19822 15802
rect 19526 15748 19582 15750
rect 19606 15748 19662 15750
rect 19686 15748 19742 15750
rect 19766 15748 19822 15750
rect 20186 15258 20242 15260
rect 20266 15258 20322 15260
rect 20346 15258 20402 15260
rect 20426 15258 20482 15260
rect 20186 15206 20232 15258
rect 20232 15206 20242 15258
rect 20266 15206 20296 15258
rect 20296 15206 20308 15258
rect 20308 15206 20322 15258
rect 20346 15206 20360 15258
rect 20360 15206 20372 15258
rect 20372 15206 20402 15258
rect 20426 15206 20436 15258
rect 20436 15206 20482 15258
rect 20186 15204 20242 15206
rect 20266 15204 20322 15206
rect 20346 15204 20402 15206
rect 20426 15204 20482 15206
rect 19526 14714 19582 14716
rect 19606 14714 19662 14716
rect 19686 14714 19742 14716
rect 19766 14714 19822 14716
rect 19526 14662 19572 14714
rect 19572 14662 19582 14714
rect 19606 14662 19636 14714
rect 19636 14662 19648 14714
rect 19648 14662 19662 14714
rect 19686 14662 19700 14714
rect 19700 14662 19712 14714
rect 19712 14662 19742 14714
rect 19766 14662 19776 14714
rect 19776 14662 19822 14714
rect 19526 14660 19582 14662
rect 19606 14660 19662 14662
rect 19686 14660 19742 14662
rect 19766 14660 19822 14662
rect 18234 12280 18290 12336
rect 20186 14170 20242 14172
rect 20266 14170 20322 14172
rect 20346 14170 20402 14172
rect 20426 14170 20482 14172
rect 20186 14118 20232 14170
rect 20232 14118 20242 14170
rect 20266 14118 20296 14170
rect 20296 14118 20308 14170
rect 20308 14118 20322 14170
rect 20346 14118 20360 14170
rect 20360 14118 20372 14170
rect 20372 14118 20402 14170
rect 20426 14118 20436 14170
rect 20436 14118 20482 14170
rect 20186 14116 20242 14118
rect 20266 14116 20322 14118
rect 20346 14116 20402 14118
rect 20426 14116 20482 14118
rect 19526 13626 19582 13628
rect 19606 13626 19662 13628
rect 19686 13626 19742 13628
rect 19766 13626 19822 13628
rect 19526 13574 19572 13626
rect 19572 13574 19582 13626
rect 19606 13574 19636 13626
rect 19636 13574 19648 13626
rect 19648 13574 19662 13626
rect 19686 13574 19700 13626
rect 19700 13574 19712 13626
rect 19712 13574 19742 13626
rect 19766 13574 19776 13626
rect 19776 13574 19822 13626
rect 19526 13572 19582 13574
rect 19606 13572 19662 13574
rect 19686 13572 19742 13574
rect 19766 13572 19822 13574
rect 20186 13082 20242 13084
rect 20266 13082 20322 13084
rect 20346 13082 20402 13084
rect 20426 13082 20482 13084
rect 20186 13030 20232 13082
rect 20232 13030 20242 13082
rect 20266 13030 20296 13082
rect 20296 13030 20308 13082
rect 20308 13030 20322 13082
rect 20346 13030 20360 13082
rect 20360 13030 20372 13082
rect 20372 13030 20402 13082
rect 20426 13030 20436 13082
rect 20436 13030 20482 13082
rect 20186 13028 20242 13030
rect 20266 13028 20322 13030
rect 20346 13028 20402 13030
rect 20426 13028 20482 13030
rect 19526 12538 19582 12540
rect 19606 12538 19662 12540
rect 19686 12538 19742 12540
rect 19766 12538 19822 12540
rect 19526 12486 19572 12538
rect 19572 12486 19582 12538
rect 19606 12486 19636 12538
rect 19636 12486 19648 12538
rect 19648 12486 19662 12538
rect 19686 12486 19700 12538
rect 19700 12486 19712 12538
rect 19712 12486 19742 12538
rect 19766 12486 19776 12538
rect 19776 12486 19822 12538
rect 19526 12484 19582 12486
rect 19606 12484 19662 12486
rect 19686 12484 19742 12486
rect 19766 12484 19822 12486
rect 19526 11450 19582 11452
rect 19606 11450 19662 11452
rect 19686 11450 19742 11452
rect 19766 11450 19822 11452
rect 19526 11398 19572 11450
rect 19572 11398 19582 11450
rect 19606 11398 19636 11450
rect 19636 11398 19648 11450
rect 19648 11398 19662 11450
rect 19686 11398 19700 11450
rect 19700 11398 19712 11450
rect 19712 11398 19742 11450
rect 19766 11398 19776 11450
rect 19776 11398 19822 11450
rect 19526 11396 19582 11398
rect 19606 11396 19662 11398
rect 19686 11396 19742 11398
rect 19766 11396 19822 11398
rect 19526 10362 19582 10364
rect 19606 10362 19662 10364
rect 19686 10362 19742 10364
rect 19766 10362 19822 10364
rect 19526 10310 19572 10362
rect 19572 10310 19582 10362
rect 19606 10310 19636 10362
rect 19636 10310 19648 10362
rect 19648 10310 19662 10362
rect 19686 10310 19700 10362
rect 19700 10310 19712 10362
rect 19712 10310 19742 10362
rect 19766 10310 19776 10362
rect 19776 10310 19822 10362
rect 19526 10308 19582 10310
rect 19606 10308 19662 10310
rect 19686 10308 19742 10310
rect 19766 10308 19822 10310
rect 19798 10124 19854 10160
rect 19798 10104 19800 10124
rect 19800 10104 19852 10124
rect 19852 10104 19854 10124
rect 20442 12164 20498 12200
rect 20442 12144 20444 12164
rect 20444 12144 20496 12164
rect 20496 12144 20498 12164
rect 20186 11994 20242 11996
rect 20266 11994 20322 11996
rect 20346 11994 20402 11996
rect 20426 11994 20482 11996
rect 20186 11942 20232 11994
rect 20232 11942 20242 11994
rect 20266 11942 20296 11994
rect 20296 11942 20308 11994
rect 20308 11942 20322 11994
rect 20346 11942 20360 11994
rect 20360 11942 20372 11994
rect 20372 11942 20402 11994
rect 20426 11942 20436 11994
rect 20436 11942 20482 11994
rect 20186 11940 20242 11942
rect 20266 11940 20322 11942
rect 20346 11940 20402 11942
rect 20426 11940 20482 11942
rect 19526 9274 19582 9276
rect 19606 9274 19662 9276
rect 19686 9274 19742 9276
rect 19766 9274 19822 9276
rect 19526 9222 19572 9274
rect 19572 9222 19582 9274
rect 19606 9222 19636 9274
rect 19636 9222 19648 9274
rect 19648 9222 19662 9274
rect 19686 9222 19700 9274
rect 19700 9222 19712 9274
rect 19712 9222 19742 9274
rect 19766 9222 19776 9274
rect 19776 9222 19822 9274
rect 19526 9220 19582 9222
rect 19606 9220 19662 9222
rect 19686 9220 19742 9222
rect 19766 9220 19822 9222
rect 20186 10906 20242 10908
rect 20266 10906 20322 10908
rect 20346 10906 20402 10908
rect 20426 10906 20482 10908
rect 20186 10854 20232 10906
rect 20232 10854 20242 10906
rect 20266 10854 20296 10906
rect 20296 10854 20308 10906
rect 20308 10854 20322 10906
rect 20346 10854 20360 10906
rect 20360 10854 20372 10906
rect 20372 10854 20402 10906
rect 20426 10854 20436 10906
rect 20436 10854 20482 10906
rect 20186 10852 20242 10854
rect 20266 10852 20322 10854
rect 20346 10852 20402 10854
rect 20426 10852 20482 10854
rect 20166 10140 20168 10160
rect 20168 10140 20220 10160
rect 20220 10140 20222 10160
rect 20166 10104 20222 10140
rect 21454 14340 21510 14376
rect 21454 14320 21456 14340
rect 21456 14320 21508 14340
rect 21508 14320 21510 14340
rect 21270 12180 21272 12200
rect 21272 12180 21324 12200
rect 21324 12180 21326 12200
rect 21270 12144 21326 12180
rect 20186 9818 20242 9820
rect 20266 9818 20322 9820
rect 20346 9818 20402 9820
rect 20426 9818 20482 9820
rect 20186 9766 20232 9818
rect 20232 9766 20242 9818
rect 20266 9766 20296 9818
rect 20296 9766 20308 9818
rect 20308 9766 20322 9818
rect 20346 9766 20360 9818
rect 20360 9766 20372 9818
rect 20372 9766 20402 9818
rect 20426 9766 20436 9818
rect 20436 9766 20482 9818
rect 20186 9764 20242 9766
rect 20266 9764 20322 9766
rect 20346 9764 20402 9766
rect 20426 9764 20482 9766
rect 20534 9424 20590 9480
rect 20186 8730 20242 8732
rect 20266 8730 20322 8732
rect 20346 8730 20402 8732
rect 20426 8730 20482 8732
rect 20186 8678 20232 8730
rect 20232 8678 20242 8730
rect 20266 8678 20296 8730
rect 20296 8678 20308 8730
rect 20308 8678 20322 8730
rect 20346 8678 20360 8730
rect 20360 8678 20372 8730
rect 20372 8678 20402 8730
rect 20426 8678 20436 8730
rect 20436 8678 20482 8730
rect 20186 8676 20242 8678
rect 20266 8676 20322 8678
rect 20346 8676 20402 8678
rect 20426 8676 20482 8678
rect 19526 8186 19582 8188
rect 19606 8186 19662 8188
rect 19686 8186 19742 8188
rect 19766 8186 19822 8188
rect 19526 8134 19572 8186
rect 19572 8134 19582 8186
rect 19606 8134 19636 8186
rect 19636 8134 19648 8186
rect 19648 8134 19662 8186
rect 19686 8134 19700 8186
rect 19700 8134 19712 8186
rect 19712 8134 19742 8186
rect 19766 8134 19776 8186
rect 19776 8134 19822 8186
rect 19526 8132 19582 8134
rect 19606 8132 19662 8134
rect 19686 8132 19742 8134
rect 19766 8132 19822 8134
rect 20186 7642 20242 7644
rect 20266 7642 20322 7644
rect 20346 7642 20402 7644
rect 20426 7642 20482 7644
rect 20186 7590 20232 7642
rect 20232 7590 20242 7642
rect 20266 7590 20296 7642
rect 20296 7590 20308 7642
rect 20308 7590 20322 7642
rect 20346 7590 20360 7642
rect 20360 7590 20372 7642
rect 20372 7590 20402 7642
rect 20426 7590 20436 7642
rect 20436 7590 20482 7642
rect 20186 7588 20242 7590
rect 20266 7588 20322 7590
rect 20346 7588 20402 7590
rect 20426 7588 20482 7590
rect 19526 7098 19582 7100
rect 19606 7098 19662 7100
rect 19686 7098 19742 7100
rect 19766 7098 19822 7100
rect 19526 7046 19572 7098
rect 19572 7046 19582 7098
rect 19606 7046 19636 7098
rect 19636 7046 19648 7098
rect 19648 7046 19662 7098
rect 19686 7046 19700 7098
rect 19700 7046 19712 7098
rect 19712 7046 19742 7098
rect 19766 7046 19776 7098
rect 19776 7046 19822 7098
rect 19526 7044 19582 7046
rect 19606 7044 19662 7046
rect 19686 7044 19742 7046
rect 19766 7044 19822 7046
rect 23662 16532 23664 16552
rect 23664 16532 23716 16552
rect 23716 16532 23718 16552
rect 23662 16496 23718 16532
rect 26954 23418 27010 23420
rect 27034 23418 27090 23420
rect 27114 23418 27170 23420
rect 27194 23418 27250 23420
rect 26954 23366 27000 23418
rect 27000 23366 27010 23418
rect 27034 23366 27064 23418
rect 27064 23366 27076 23418
rect 27076 23366 27090 23418
rect 27114 23366 27128 23418
rect 27128 23366 27140 23418
rect 27140 23366 27170 23418
rect 27194 23366 27204 23418
rect 27204 23366 27250 23418
rect 26954 23364 27010 23366
rect 27034 23364 27090 23366
rect 27114 23364 27170 23366
rect 27194 23364 27250 23366
rect 30286 23160 30342 23216
rect 27614 22874 27670 22876
rect 27694 22874 27750 22876
rect 27774 22874 27830 22876
rect 27854 22874 27910 22876
rect 27614 22822 27660 22874
rect 27660 22822 27670 22874
rect 27694 22822 27724 22874
rect 27724 22822 27736 22874
rect 27736 22822 27750 22874
rect 27774 22822 27788 22874
rect 27788 22822 27800 22874
rect 27800 22822 27830 22874
rect 27854 22822 27864 22874
rect 27864 22822 27910 22874
rect 27614 22820 27670 22822
rect 27694 22820 27750 22822
rect 27774 22820 27830 22822
rect 27854 22820 27910 22822
rect 30930 22480 30986 22536
rect 26954 22330 27010 22332
rect 27034 22330 27090 22332
rect 27114 22330 27170 22332
rect 27194 22330 27250 22332
rect 26954 22278 27000 22330
rect 27000 22278 27010 22330
rect 27034 22278 27064 22330
rect 27064 22278 27076 22330
rect 27076 22278 27090 22330
rect 27114 22278 27128 22330
rect 27128 22278 27140 22330
rect 27140 22278 27170 22330
rect 27194 22278 27204 22330
rect 27204 22278 27250 22330
rect 26954 22276 27010 22278
rect 27034 22276 27090 22278
rect 27114 22276 27170 22278
rect 27194 22276 27250 22278
rect 27614 21786 27670 21788
rect 27694 21786 27750 21788
rect 27774 21786 27830 21788
rect 27854 21786 27910 21788
rect 27614 21734 27660 21786
rect 27660 21734 27670 21786
rect 27694 21734 27724 21786
rect 27724 21734 27736 21786
rect 27736 21734 27750 21786
rect 27774 21734 27788 21786
rect 27788 21734 27800 21786
rect 27800 21734 27830 21786
rect 27854 21734 27864 21786
rect 27864 21734 27910 21786
rect 27614 21732 27670 21734
rect 27694 21732 27750 21734
rect 27774 21732 27830 21734
rect 27854 21732 27910 21734
rect 26954 21242 27010 21244
rect 27034 21242 27090 21244
rect 27114 21242 27170 21244
rect 27194 21242 27250 21244
rect 26954 21190 27000 21242
rect 27000 21190 27010 21242
rect 27034 21190 27064 21242
rect 27064 21190 27076 21242
rect 27076 21190 27090 21242
rect 27114 21190 27128 21242
rect 27128 21190 27140 21242
rect 27140 21190 27170 21242
rect 27194 21190 27204 21242
rect 27204 21190 27250 21242
rect 26954 21188 27010 21190
rect 27034 21188 27090 21190
rect 27114 21188 27170 21190
rect 27194 21188 27250 21190
rect 30470 21800 30526 21856
rect 30378 21120 30434 21176
rect 27614 20698 27670 20700
rect 27694 20698 27750 20700
rect 27774 20698 27830 20700
rect 27854 20698 27910 20700
rect 27614 20646 27660 20698
rect 27660 20646 27670 20698
rect 27694 20646 27724 20698
rect 27724 20646 27736 20698
rect 27736 20646 27750 20698
rect 27774 20646 27788 20698
rect 27788 20646 27800 20698
rect 27800 20646 27830 20698
rect 27854 20646 27864 20698
rect 27864 20646 27910 20698
rect 27614 20644 27670 20646
rect 27694 20644 27750 20646
rect 27774 20644 27830 20646
rect 27854 20644 27910 20646
rect 30286 20440 30342 20496
rect 26954 20154 27010 20156
rect 27034 20154 27090 20156
rect 27114 20154 27170 20156
rect 27194 20154 27250 20156
rect 26954 20102 27000 20154
rect 27000 20102 27010 20154
rect 27034 20102 27064 20154
rect 27064 20102 27076 20154
rect 27076 20102 27090 20154
rect 27114 20102 27128 20154
rect 27128 20102 27140 20154
rect 27140 20102 27170 20154
rect 27194 20102 27204 20154
rect 27204 20102 27250 20154
rect 26954 20100 27010 20102
rect 27034 20100 27090 20102
rect 27114 20100 27170 20102
rect 27194 20100 27250 20102
rect 30378 19760 30434 19816
rect 27614 19610 27670 19612
rect 27694 19610 27750 19612
rect 27774 19610 27830 19612
rect 27854 19610 27910 19612
rect 27614 19558 27660 19610
rect 27660 19558 27670 19610
rect 27694 19558 27724 19610
rect 27724 19558 27736 19610
rect 27736 19558 27750 19610
rect 27774 19558 27788 19610
rect 27788 19558 27800 19610
rect 27800 19558 27830 19610
rect 27854 19558 27864 19610
rect 27864 19558 27910 19610
rect 27614 19556 27670 19558
rect 27694 19556 27750 19558
rect 27774 19556 27830 19558
rect 27854 19556 27910 19558
rect 30286 19080 30342 19136
rect 26954 19066 27010 19068
rect 27034 19066 27090 19068
rect 27114 19066 27170 19068
rect 27194 19066 27250 19068
rect 26954 19014 27000 19066
rect 27000 19014 27010 19066
rect 27034 19014 27064 19066
rect 27064 19014 27076 19066
rect 27076 19014 27090 19066
rect 27114 19014 27128 19066
rect 27128 19014 27140 19066
rect 27140 19014 27170 19066
rect 27194 19014 27204 19066
rect 27204 19014 27250 19066
rect 26954 19012 27010 19014
rect 27034 19012 27090 19014
rect 27114 19012 27170 19014
rect 27194 19012 27250 19014
rect 27614 18522 27670 18524
rect 27694 18522 27750 18524
rect 27774 18522 27830 18524
rect 27854 18522 27910 18524
rect 27614 18470 27660 18522
rect 27660 18470 27670 18522
rect 27694 18470 27724 18522
rect 27724 18470 27736 18522
rect 27736 18470 27750 18522
rect 27774 18470 27788 18522
rect 27788 18470 27800 18522
rect 27800 18470 27830 18522
rect 27854 18470 27864 18522
rect 27864 18470 27910 18522
rect 27614 18468 27670 18470
rect 27694 18468 27750 18470
rect 27774 18468 27830 18470
rect 27854 18468 27910 18470
rect 30378 18400 30434 18456
rect 26954 17978 27010 17980
rect 27034 17978 27090 17980
rect 27114 17978 27170 17980
rect 27194 17978 27250 17980
rect 26954 17926 27000 17978
rect 27000 17926 27010 17978
rect 27034 17926 27064 17978
rect 27064 17926 27076 17978
rect 27076 17926 27090 17978
rect 27114 17926 27128 17978
rect 27128 17926 27140 17978
rect 27140 17926 27170 17978
rect 27194 17926 27204 17978
rect 27204 17926 27250 17978
rect 26954 17924 27010 17926
rect 27034 17924 27090 17926
rect 27114 17924 27170 17926
rect 27194 17924 27250 17926
rect 30286 17720 30342 17776
rect 27614 17434 27670 17436
rect 27694 17434 27750 17436
rect 27774 17434 27830 17436
rect 27854 17434 27910 17436
rect 27614 17382 27660 17434
rect 27660 17382 27670 17434
rect 27694 17382 27724 17434
rect 27724 17382 27736 17434
rect 27736 17382 27750 17434
rect 27774 17382 27788 17434
rect 27788 17382 27800 17434
rect 27800 17382 27830 17434
rect 27854 17382 27864 17434
rect 27864 17382 27910 17434
rect 27614 17380 27670 17382
rect 27694 17380 27750 17382
rect 27774 17380 27830 17382
rect 27854 17380 27910 17382
rect 26954 16890 27010 16892
rect 27034 16890 27090 16892
rect 27114 16890 27170 16892
rect 27194 16890 27250 16892
rect 26954 16838 27000 16890
rect 27000 16838 27010 16890
rect 27034 16838 27064 16890
rect 27064 16838 27076 16890
rect 27076 16838 27090 16890
rect 27114 16838 27128 16890
rect 27128 16838 27140 16890
rect 27140 16838 27170 16890
rect 27194 16838 27204 16890
rect 27204 16838 27250 16890
rect 26954 16836 27010 16838
rect 27034 16836 27090 16838
rect 27114 16836 27170 16838
rect 27194 16836 27250 16838
rect 30378 17060 30434 17096
rect 30378 17040 30380 17060
rect 30380 17040 30432 17060
rect 30432 17040 30434 17060
rect 30930 16360 30986 16416
rect 27614 16346 27670 16348
rect 27694 16346 27750 16348
rect 27774 16346 27830 16348
rect 27854 16346 27910 16348
rect 27614 16294 27660 16346
rect 27660 16294 27670 16346
rect 27694 16294 27724 16346
rect 27724 16294 27736 16346
rect 27736 16294 27750 16346
rect 27774 16294 27788 16346
rect 27788 16294 27800 16346
rect 27800 16294 27830 16346
rect 27854 16294 27864 16346
rect 27864 16294 27910 16346
rect 27614 16292 27670 16294
rect 27694 16292 27750 16294
rect 27774 16292 27830 16294
rect 27854 16292 27910 16294
rect 26954 15802 27010 15804
rect 27034 15802 27090 15804
rect 27114 15802 27170 15804
rect 27194 15802 27250 15804
rect 26954 15750 27000 15802
rect 27000 15750 27010 15802
rect 27034 15750 27064 15802
rect 27064 15750 27076 15802
rect 27076 15750 27090 15802
rect 27114 15750 27128 15802
rect 27128 15750 27140 15802
rect 27140 15750 27170 15802
rect 27194 15750 27204 15802
rect 27204 15750 27250 15802
rect 26954 15748 27010 15750
rect 27034 15748 27090 15750
rect 27114 15748 27170 15750
rect 27194 15748 27250 15750
rect 30378 15680 30434 15736
rect 27614 15258 27670 15260
rect 27694 15258 27750 15260
rect 27774 15258 27830 15260
rect 27854 15258 27910 15260
rect 27614 15206 27660 15258
rect 27660 15206 27670 15258
rect 27694 15206 27724 15258
rect 27724 15206 27736 15258
rect 27736 15206 27750 15258
rect 27774 15206 27788 15258
rect 27788 15206 27800 15258
rect 27800 15206 27830 15258
rect 27854 15206 27864 15258
rect 27864 15206 27910 15258
rect 27614 15204 27670 15206
rect 27694 15204 27750 15206
rect 27774 15204 27830 15206
rect 27854 15204 27910 15206
rect 30286 15000 30342 15056
rect 26954 14714 27010 14716
rect 27034 14714 27090 14716
rect 27114 14714 27170 14716
rect 27194 14714 27250 14716
rect 26954 14662 27000 14714
rect 27000 14662 27010 14714
rect 27034 14662 27064 14714
rect 27064 14662 27076 14714
rect 27076 14662 27090 14714
rect 27114 14662 27128 14714
rect 27128 14662 27140 14714
rect 27140 14662 27170 14714
rect 27194 14662 27204 14714
rect 27204 14662 27250 14714
rect 26954 14660 27010 14662
rect 27034 14660 27090 14662
rect 27114 14660 27170 14662
rect 27194 14660 27250 14662
rect 30378 14320 30434 14376
rect 27614 14170 27670 14172
rect 27694 14170 27750 14172
rect 27774 14170 27830 14172
rect 27854 14170 27910 14172
rect 27614 14118 27660 14170
rect 27660 14118 27670 14170
rect 27694 14118 27724 14170
rect 27724 14118 27736 14170
rect 27736 14118 27750 14170
rect 27774 14118 27788 14170
rect 27788 14118 27800 14170
rect 27800 14118 27830 14170
rect 27854 14118 27864 14170
rect 27864 14118 27910 14170
rect 27614 14116 27670 14118
rect 27694 14116 27750 14118
rect 27774 14116 27830 14118
rect 27854 14116 27910 14118
rect 26954 13626 27010 13628
rect 27034 13626 27090 13628
rect 27114 13626 27170 13628
rect 27194 13626 27250 13628
rect 26954 13574 27000 13626
rect 27000 13574 27010 13626
rect 27034 13574 27064 13626
rect 27064 13574 27076 13626
rect 27076 13574 27090 13626
rect 27114 13574 27128 13626
rect 27128 13574 27140 13626
rect 27140 13574 27170 13626
rect 27194 13574 27204 13626
rect 27204 13574 27250 13626
rect 26954 13572 27010 13574
rect 27034 13572 27090 13574
rect 27114 13572 27170 13574
rect 27194 13572 27250 13574
rect 27614 13082 27670 13084
rect 27694 13082 27750 13084
rect 27774 13082 27830 13084
rect 27854 13082 27910 13084
rect 27614 13030 27660 13082
rect 27660 13030 27670 13082
rect 27694 13030 27724 13082
rect 27724 13030 27736 13082
rect 27736 13030 27750 13082
rect 27774 13030 27788 13082
rect 27788 13030 27800 13082
rect 27800 13030 27830 13082
rect 27854 13030 27864 13082
rect 27864 13030 27910 13082
rect 27614 13028 27670 13030
rect 27694 13028 27750 13030
rect 27774 13028 27830 13030
rect 27854 13028 27910 13030
rect 30286 13640 30342 13696
rect 30378 12960 30434 13016
rect 26954 12538 27010 12540
rect 27034 12538 27090 12540
rect 27114 12538 27170 12540
rect 27194 12538 27250 12540
rect 26954 12486 27000 12538
rect 27000 12486 27010 12538
rect 27034 12486 27064 12538
rect 27064 12486 27076 12538
rect 27076 12486 27090 12538
rect 27114 12486 27128 12538
rect 27128 12486 27140 12538
rect 27140 12486 27170 12538
rect 27194 12486 27204 12538
rect 27204 12486 27250 12538
rect 26954 12484 27010 12486
rect 27034 12484 27090 12486
rect 27114 12484 27170 12486
rect 27194 12484 27250 12486
rect 30286 12280 30342 12336
rect 27614 11994 27670 11996
rect 27694 11994 27750 11996
rect 27774 11994 27830 11996
rect 27854 11994 27910 11996
rect 27614 11942 27660 11994
rect 27660 11942 27670 11994
rect 27694 11942 27724 11994
rect 27724 11942 27736 11994
rect 27736 11942 27750 11994
rect 27774 11942 27788 11994
rect 27788 11942 27800 11994
rect 27800 11942 27830 11994
rect 27854 11942 27864 11994
rect 27864 11942 27910 11994
rect 27614 11940 27670 11942
rect 27694 11940 27750 11942
rect 27774 11940 27830 11942
rect 27854 11940 27910 11942
rect 26954 11450 27010 11452
rect 27034 11450 27090 11452
rect 27114 11450 27170 11452
rect 27194 11450 27250 11452
rect 26954 11398 27000 11450
rect 27000 11398 27010 11450
rect 27034 11398 27064 11450
rect 27064 11398 27076 11450
rect 27076 11398 27090 11450
rect 27114 11398 27128 11450
rect 27128 11398 27140 11450
rect 27140 11398 27170 11450
rect 27194 11398 27204 11450
rect 27204 11398 27250 11450
rect 26954 11396 27010 11398
rect 27034 11396 27090 11398
rect 27114 11396 27170 11398
rect 27194 11396 27250 11398
rect 30378 11620 30434 11656
rect 30378 11600 30380 11620
rect 30380 11600 30432 11620
rect 30432 11600 30434 11620
rect 30286 10920 30342 10976
rect 27614 10906 27670 10908
rect 27694 10906 27750 10908
rect 27774 10906 27830 10908
rect 27854 10906 27910 10908
rect 27614 10854 27660 10906
rect 27660 10854 27670 10906
rect 27694 10854 27724 10906
rect 27724 10854 27736 10906
rect 27736 10854 27750 10906
rect 27774 10854 27788 10906
rect 27788 10854 27800 10906
rect 27800 10854 27830 10906
rect 27854 10854 27864 10906
rect 27864 10854 27910 10906
rect 27614 10852 27670 10854
rect 27694 10852 27750 10854
rect 27774 10852 27830 10854
rect 27854 10852 27910 10854
rect 26954 10362 27010 10364
rect 27034 10362 27090 10364
rect 27114 10362 27170 10364
rect 27194 10362 27250 10364
rect 26954 10310 27000 10362
rect 27000 10310 27010 10362
rect 27034 10310 27064 10362
rect 27064 10310 27076 10362
rect 27076 10310 27090 10362
rect 27114 10310 27128 10362
rect 27128 10310 27140 10362
rect 27140 10310 27170 10362
rect 27194 10310 27204 10362
rect 27204 10310 27250 10362
rect 26954 10308 27010 10310
rect 27034 10308 27090 10310
rect 27114 10308 27170 10310
rect 27194 10308 27250 10310
rect 30930 10240 30986 10296
rect 27614 9818 27670 9820
rect 27694 9818 27750 9820
rect 27774 9818 27830 9820
rect 27854 9818 27910 9820
rect 27614 9766 27660 9818
rect 27660 9766 27670 9818
rect 27694 9766 27724 9818
rect 27724 9766 27736 9818
rect 27736 9766 27750 9818
rect 27774 9766 27788 9818
rect 27788 9766 27800 9818
rect 27800 9766 27830 9818
rect 27854 9766 27864 9818
rect 27864 9766 27910 9818
rect 27614 9764 27670 9766
rect 27694 9764 27750 9766
rect 27774 9764 27830 9766
rect 27854 9764 27910 9766
rect 30286 9560 30342 9616
rect 25318 9424 25374 9480
rect 26954 9274 27010 9276
rect 27034 9274 27090 9276
rect 27114 9274 27170 9276
rect 27194 9274 27250 9276
rect 26954 9222 27000 9274
rect 27000 9222 27010 9274
rect 27034 9222 27064 9274
rect 27064 9222 27076 9274
rect 27076 9222 27090 9274
rect 27114 9222 27128 9274
rect 27128 9222 27140 9274
rect 27140 9222 27170 9274
rect 27194 9222 27204 9274
rect 27204 9222 27250 9274
rect 26954 9220 27010 9222
rect 27034 9220 27090 9222
rect 27114 9220 27170 9222
rect 27194 9220 27250 9222
rect 30378 8880 30434 8936
rect 27614 8730 27670 8732
rect 27694 8730 27750 8732
rect 27774 8730 27830 8732
rect 27854 8730 27910 8732
rect 27614 8678 27660 8730
rect 27660 8678 27670 8730
rect 27694 8678 27724 8730
rect 27724 8678 27736 8730
rect 27736 8678 27750 8730
rect 27774 8678 27788 8730
rect 27788 8678 27800 8730
rect 27800 8678 27830 8730
rect 27854 8678 27864 8730
rect 27864 8678 27910 8730
rect 27614 8676 27670 8678
rect 27694 8676 27750 8678
rect 27774 8676 27830 8678
rect 27854 8676 27910 8678
rect 30286 8200 30342 8256
rect 26954 8186 27010 8188
rect 27034 8186 27090 8188
rect 27114 8186 27170 8188
rect 27194 8186 27250 8188
rect 26954 8134 27000 8186
rect 27000 8134 27010 8186
rect 27034 8134 27064 8186
rect 27064 8134 27076 8186
rect 27076 8134 27090 8186
rect 27114 8134 27128 8186
rect 27128 8134 27140 8186
rect 27140 8134 27170 8186
rect 27194 8134 27204 8186
rect 27204 8134 27250 8186
rect 26954 8132 27010 8134
rect 27034 8132 27090 8134
rect 27114 8132 27170 8134
rect 27194 8132 27250 8134
rect 20186 6554 20242 6556
rect 20266 6554 20322 6556
rect 20346 6554 20402 6556
rect 20426 6554 20482 6556
rect 20186 6502 20232 6554
rect 20232 6502 20242 6554
rect 20266 6502 20296 6554
rect 20296 6502 20308 6554
rect 20308 6502 20322 6554
rect 20346 6502 20360 6554
rect 20360 6502 20372 6554
rect 20372 6502 20402 6554
rect 20426 6502 20436 6554
rect 20436 6502 20482 6554
rect 20186 6500 20242 6502
rect 20266 6500 20322 6502
rect 20346 6500 20402 6502
rect 20426 6500 20482 6502
rect 19526 6010 19582 6012
rect 19606 6010 19662 6012
rect 19686 6010 19742 6012
rect 19766 6010 19822 6012
rect 19526 5958 19572 6010
rect 19572 5958 19582 6010
rect 19606 5958 19636 6010
rect 19636 5958 19648 6010
rect 19648 5958 19662 6010
rect 19686 5958 19700 6010
rect 19700 5958 19712 6010
rect 19712 5958 19742 6010
rect 19766 5958 19776 6010
rect 19776 5958 19822 6010
rect 19526 5956 19582 5958
rect 19606 5956 19662 5958
rect 19686 5956 19742 5958
rect 19766 5956 19822 5958
rect 20186 5466 20242 5468
rect 20266 5466 20322 5468
rect 20346 5466 20402 5468
rect 20426 5466 20482 5468
rect 20186 5414 20232 5466
rect 20232 5414 20242 5466
rect 20266 5414 20296 5466
rect 20296 5414 20308 5466
rect 20308 5414 20322 5466
rect 20346 5414 20360 5466
rect 20360 5414 20372 5466
rect 20372 5414 20402 5466
rect 20426 5414 20436 5466
rect 20436 5414 20482 5466
rect 20186 5412 20242 5414
rect 20266 5412 20322 5414
rect 20346 5412 20402 5414
rect 20426 5412 20482 5414
rect 19526 4922 19582 4924
rect 19606 4922 19662 4924
rect 19686 4922 19742 4924
rect 19766 4922 19822 4924
rect 19526 4870 19572 4922
rect 19572 4870 19582 4922
rect 19606 4870 19636 4922
rect 19636 4870 19648 4922
rect 19648 4870 19662 4922
rect 19686 4870 19700 4922
rect 19700 4870 19712 4922
rect 19712 4870 19742 4922
rect 19766 4870 19776 4922
rect 19776 4870 19822 4922
rect 19526 4868 19582 4870
rect 19606 4868 19662 4870
rect 19686 4868 19742 4870
rect 19766 4868 19822 4870
rect 20186 4378 20242 4380
rect 20266 4378 20322 4380
rect 20346 4378 20402 4380
rect 20426 4378 20482 4380
rect 20186 4326 20232 4378
rect 20232 4326 20242 4378
rect 20266 4326 20296 4378
rect 20296 4326 20308 4378
rect 20308 4326 20322 4378
rect 20346 4326 20360 4378
rect 20360 4326 20372 4378
rect 20372 4326 20402 4378
rect 20426 4326 20436 4378
rect 20436 4326 20482 4378
rect 20186 4324 20242 4326
rect 20266 4324 20322 4326
rect 20346 4324 20402 4326
rect 20426 4324 20482 4326
rect 19526 3834 19582 3836
rect 19606 3834 19662 3836
rect 19686 3834 19742 3836
rect 19766 3834 19822 3836
rect 19526 3782 19572 3834
rect 19572 3782 19582 3834
rect 19606 3782 19636 3834
rect 19636 3782 19648 3834
rect 19648 3782 19662 3834
rect 19686 3782 19700 3834
rect 19700 3782 19712 3834
rect 19712 3782 19742 3834
rect 19766 3782 19776 3834
rect 19776 3782 19822 3834
rect 19526 3780 19582 3782
rect 19606 3780 19662 3782
rect 19686 3780 19742 3782
rect 19766 3780 19822 3782
rect 20186 3290 20242 3292
rect 20266 3290 20322 3292
rect 20346 3290 20402 3292
rect 20426 3290 20482 3292
rect 20186 3238 20232 3290
rect 20232 3238 20242 3290
rect 20266 3238 20296 3290
rect 20296 3238 20308 3290
rect 20308 3238 20322 3290
rect 20346 3238 20360 3290
rect 20360 3238 20372 3290
rect 20372 3238 20402 3290
rect 20426 3238 20436 3290
rect 20436 3238 20482 3290
rect 20186 3236 20242 3238
rect 20266 3236 20322 3238
rect 20346 3236 20402 3238
rect 20426 3236 20482 3238
rect 19526 2746 19582 2748
rect 19606 2746 19662 2748
rect 19686 2746 19742 2748
rect 19766 2746 19822 2748
rect 19526 2694 19572 2746
rect 19572 2694 19582 2746
rect 19606 2694 19636 2746
rect 19636 2694 19648 2746
rect 19648 2694 19662 2746
rect 19686 2694 19700 2746
rect 19700 2694 19712 2746
rect 19712 2694 19742 2746
rect 19766 2694 19776 2746
rect 19776 2694 19822 2746
rect 19526 2692 19582 2694
rect 19606 2692 19662 2694
rect 19686 2692 19742 2694
rect 19766 2692 19822 2694
rect 27614 7642 27670 7644
rect 27694 7642 27750 7644
rect 27774 7642 27830 7644
rect 27854 7642 27910 7644
rect 27614 7590 27660 7642
rect 27660 7590 27670 7642
rect 27694 7590 27724 7642
rect 27724 7590 27736 7642
rect 27736 7590 27750 7642
rect 27774 7590 27788 7642
rect 27788 7590 27800 7642
rect 27800 7590 27830 7642
rect 27854 7590 27864 7642
rect 27864 7590 27910 7642
rect 27614 7588 27670 7590
rect 27694 7588 27750 7590
rect 27774 7588 27830 7590
rect 27854 7588 27910 7590
rect 26954 7098 27010 7100
rect 27034 7098 27090 7100
rect 27114 7098 27170 7100
rect 27194 7098 27250 7100
rect 26954 7046 27000 7098
rect 27000 7046 27010 7098
rect 27034 7046 27064 7098
rect 27064 7046 27076 7098
rect 27076 7046 27090 7098
rect 27114 7046 27128 7098
rect 27128 7046 27140 7098
rect 27140 7046 27170 7098
rect 27194 7046 27204 7098
rect 27204 7046 27250 7098
rect 26954 7044 27010 7046
rect 27034 7044 27090 7046
rect 27114 7044 27170 7046
rect 27194 7044 27250 7046
rect 27614 6554 27670 6556
rect 27694 6554 27750 6556
rect 27774 6554 27830 6556
rect 27854 6554 27910 6556
rect 27614 6502 27660 6554
rect 27660 6502 27670 6554
rect 27694 6502 27724 6554
rect 27724 6502 27736 6554
rect 27736 6502 27750 6554
rect 27774 6502 27788 6554
rect 27788 6502 27800 6554
rect 27800 6502 27830 6554
rect 27854 6502 27864 6554
rect 27864 6502 27910 6554
rect 27614 6500 27670 6502
rect 27694 6500 27750 6502
rect 27774 6500 27830 6502
rect 27854 6500 27910 6502
rect 26954 6010 27010 6012
rect 27034 6010 27090 6012
rect 27114 6010 27170 6012
rect 27194 6010 27250 6012
rect 26954 5958 27000 6010
rect 27000 5958 27010 6010
rect 27034 5958 27064 6010
rect 27064 5958 27076 6010
rect 27076 5958 27090 6010
rect 27114 5958 27128 6010
rect 27128 5958 27140 6010
rect 27140 5958 27170 6010
rect 27194 5958 27204 6010
rect 27204 5958 27250 6010
rect 26954 5956 27010 5958
rect 27034 5956 27090 5958
rect 27114 5956 27170 5958
rect 27194 5956 27250 5958
rect 27614 5466 27670 5468
rect 27694 5466 27750 5468
rect 27774 5466 27830 5468
rect 27854 5466 27910 5468
rect 27614 5414 27660 5466
rect 27660 5414 27670 5466
rect 27694 5414 27724 5466
rect 27724 5414 27736 5466
rect 27736 5414 27750 5466
rect 27774 5414 27788 5466
rect 27788 5414 27800 5466
rect 27800 5414 27830 5466
rect 27854 5414 27864 5466
rect 27864 5414 27910 5466
rect 27614 5412 27670 5414
rect 27694 5412 27750 5414
rect 27774 5412 27830 5414
rect 27854 5412 27910 5414
rect 26954 4922 27010 4924
rect 27034 4922 27090 4924
rect 27114 4922 27170 4924
rect 27194 4922 27250 4924
rect 26954 4870 27000 4922
rect 27000 4870 27010 4922
rect 27034 4870 27064 4922
rect 27064 4870 27076 4922
rect 27076 4870 27090 4922
rect 27114 4870 27128 4922
rect 27128 4870 27140 4922
rect 27140 4870 27170 4922
rect 27194 4870 27204 4922
rect 27204 4870 27250 4922
rect 26954 4868 27010 4870
rect 27034 4868 27090 4870
rect 27114 4868 27170 4870
rect 27194 4868 27250 4870
rect 27614 4378 27670 4380
rect 27694 4378 27750 4380
rect 27774 4378 27830 4380
rect 27854 4378 27910 4380
rect 27614 4326 27660 4378
rect 27660 4326 27670 4378
rect 27694 4326 27724 4378
rect 27724 4326 27736 4378
rect 27736 4326 27750 4378
rect 27774 4326 27788 4378
rect 27788 4326 27800 4378
rect 27800 4326 27830 4378
rect 27854 4326 27864 4378
rect 27864 4326 27910 4378
rect 27614 4324 27670 4326
rect 27694 4324 27750 4326
rect 27774 4324 27830 4326
rect 27854 4324 27910 4326
rect 26954 3834 27010 3836
rect 27034 3834 27090 3836
rect 27114 3834 27170 3836
rect 27194 3834 27250 3836
rect 26954 3782 27000 3834
rect 27000 3782 27010 3834
rect 27034 3782 27064 3834
rect 27064 3782 27076 3834
rect 27076 3782 27090 3834
rect 27114 3782 27128 3834
rect 27128 3782 27140 3834
rect 27140 3782 27170 3834
rect 27194 3782 27204 3834
rect 27204 3782 27250 3834
rect 26954 3780 27010 3782
rect 27034 3780 27090 3782
rect 27114 3780 27170 3782
rect 27194 3780 27250 3782
rect 27614 3290 27670 3292
rect 27694 3290 27750 3292
rect 27774 3290 27830 3292
rect 27854 3290 27910 3292
rect 27614 3238 27660 3290
rect 27660 3238 27670 3290
rect 27694 3238 27724 3290
rect 27724 3238 27736 3290
rect 27736 3238 27750 3290
rect 27774 3238 27788 3290
rect 27788 3238 27800 3290
rect 27800 3238 27830 3290
rect 27854 3238 27864 3290
rect 27864 3238 27910 3290
rect 27614 3236 27670 3238
rect 27694 3236 27750 3238
rect 27774 3236 27830 3238
rect 27854 3236 27910 3238
rect 26954 2746 27010 2748
rect 27034 2746 27090 2748
rect 27114 2746 27170 2748
rect 27194 2746 27250 2748
rect 26954 2694 27000 2746
rect 27000 2694 27010 2746
rect 27034 2694 27064 2746
rect 27064 2694 27076 2746
rect 27076 2694 27090 2746
rect 27114 2694 27128 2746
rect 27128 2694 27140 2746
rect 27140 2694 27170 2746
rect 27194 2694 27204 2746
rect 27204 2694 27250 2746
rect 26954 2692 27010 2694
rect 27034 2692 27090 2694
rect 27114 2692 27170 2694
rect 27194 2692 27250 2694
rect 5330 2202 5386 2204
rect 5410 2202 5466 2204
rect 5490 2202 5546 2204
rect 5570 2202 5626 2204
rect 5330 2150 5376 2202
rect 5376 2150 5386 2202
rect 5410 2150 5440 2202
rect 5440 2150 5452 2202
rect 5452 2150 5466 2202
rect 5490 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5546 2202
rect 5570 2150 5580 2202
rect 5580 2150 5626 2202
rect 5330 2148 5386 2150
rect 5410 2148 5466 2150
rect 5490 2148 5546 2150
rect 5570 2148 5626 2150
rect 12758 2202 12814 2204
rect 12838 2202 12894 2204
rect 12918 2202 12974 2204
rect 12998 2202 13054 2204
rect 12758 2150 12804 2202
rect 12804 2150 12814 2202
rect 12838 2150 12868 2202
rect 12868 2150 12880 2202
rect 12880 2150 12894 2202
rect 12918 2150 12932 2202
rect 12932 2150 12944 2202
rect 12944 2150 12974 2202
rect 12998 2150 13008 2202
rect 13008 2150 13054 2202
rect 12758 2148 12814 2150
rect 12838 2148 12894 2150
rect 12918 2148 12974 2150
rect 12998 2148 13054 2150
rect 20186 2202 20242 2204
rect 20266 2202 20322 2204
rect 20346 2202 20402 2204
rect 20426 2202 20482 2204
rect 20186 2150 20232 2202
rect 20232 2150 20242 2202
rect 20266 2150 20296 2202
rect 20296 2150 20308 2202
rect 20308 2150 20322 2202
rect 20346 2150 20360 2202
rect 20360 2150 20372 2202
rect 20372 2150 20402 2202
rect 20426 2150 20436 2202
rect 20436 2150 20482 2202
rect 20186 2148 20242 2150
rect 20266 2148 20322 2150
rect 20346 2148 20402 2150
rect 20426 2148 20482 2150
rect 27614 2202 27670 2204
rect 27694 2202 27750 2204
rect 27774 2202 27830 2204
rect 27854 2202 27910 2204
rect 27614 2150 27660 2202
rect 27660 2150 27670 2202
rect 27694 2150 27724 2202
rect 27724 2150 27736 2202
rect 27736 2150 27750 2202
rect 27774 2150 27788 2202
rect 27788 2150 27800 2202
rect 27800 2150 27830 2202
rect 27854 2150 27864 2202
rect 27864 2150 27910 2202
rect 27614 2148 27670 2150
rect 27694 2148 27750 2150
rect 27774 2148 27830 2150
rect 27854 2148 27910 2150
<< metal3 >>
rect 5320 29408 5636 29409
rect 5320 29344 5326 29408
rect 5390 29344 5406 29408
rect 5470 29344 5486 29408
rect 5550 29344 5566 29408
rect 5630 29344 5636 29408
rect 5320 29343 5636 29344
rect 12748 29408 13064 29409
rect 12748 29344 12754 29408
rect 12818 29344 12834 29408
rect 12898 29344 12914 29408
rect 12978 29344 12994 29408
rect 13058 29344 13064 29408
rect 12748 29343 13064 29344
rect 20176 29408 20492 29409
rect 20176 29344 20182 29408
rect 20246 29344 20262 29408
rect 20326 29344 20342 29408
rect 20406 29344 20422 29408
rect 20486 29344 20492 29408
rect 20176 29343 20492 29344
rect 27604 29408 27920 29409
rect 27604 29344 27610 29408
rect 27674 29344 27690 29408
rect 27754 29344 27770 29408
rect 27834 29344 27850 29408
rect 27914 29344 27920 29408
rect 27604 29343 27920 29344
rect 4660 28864 4976 28865
rect 4660 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4976 28864
rect 4660 28799 4976 28800
rect 12088 28864 12404 28865
rect 12088 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12404 28864
rect 12088 28799 12404 28800
rect 19516 28864 19832 28865
rect 19516 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19832 28864
rect 19516 28799 19832 28800
rect 26944 28864 27260 28865
rect 26944 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27260 28864
rect 26944 28799 27260 28800
rect 5320 28320 5636 28321
rect 5320 28256 5326 28320
rect 5390 28256 5406 28320
rect 5470 28256 5486 28320
rect 5550 28256 5566 28320
rect 5630 28256 5636 28320
rect 5320 28255 5636 28256
rect 12748 28320 13064 28321
rect 12748 28256 12754 28320
rect 12818 28256 12834 28320
rect 12898 28256 12914 28320
rect 12978 28256 12994 28320
rect 13058 28256 13064 28320
rect 12748 28255 13064 28256
rect 20176 28320 20492 28321
rect 20176 28256 20182 28320
rect 20246 28256 20262 28320
rect 20326 28256 20342 28320
rect 20406 28256 20422 28320
rect 20486 28256 20492 28320
rect 20176 28255 20492 28256
rect 27604 28320 27920 28321
rect 27604 28256 27610 28320
rect 27674 28256 27690 28320
rect 27754 28256 27770 28320
rect 27834 28256 27850 28320
rect 27914 28256 27920 28320
rect 27604 28255 27920 28256
rect 4660 27776 4976 27777
rect 4660 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4976 27776
rect 4660 27711 4976 27712
rect 12088 27776 12404 27777
rect 12088 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12404 27776
rect 12088 27711 12404 27712
rect 19516 27776 19832 27777
rect 19516 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19832 27776
rect 19516 27711 19832 27712
rect 26944 27776 27260 27777
rect 26944 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27260 27776
rect 26944 27711 27260 27712
rect 5320 27232 5636 27233
rect 5320 27168 5326 27232
rect 5390 27168 5406 27232
rect 5470 27168 5486 27232
rect 5550 27168 5566 27232
rect 5630 27168 5636 27232
rect 5320 27167 5636 27168
rect 12748 27232 13064 27233
rect 12748 27168 12754 27232
rect 12818 27168 12834 27232
rect 12898 27168 12914 27232
rect 12978 27168 12994 27232
rect 13058 27168 13064 27232
rect 12748 27167 13064 27168
rect 20176 27232 20492 27233
rect 20176 27168 20182 27232
rect 20246 27168 20262 27232
rect 20326 27168 20342 27232
rect 20406 27168 20422 27232
rect 20486 27168 20492 27232
rect 20176 27167 20492 27168
rect 27604 27232 27920 27233
rect 27604 27168 27610 27232
rect 27674 27168 27690 27232
rect 27754 27168 27770 27232
rect 27834 27168 27850 27232
rect 27914 27168 27920 27232
rect 27604 27167 27920 27168
rect 4660 26688 4976 26689
rect 4660 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4976 26688
rect 4660 26623 4976 26624
rect 12088 26688 12404 26689
rect 12088 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12404 26688
rect 12088 26623 12404 26624
rect 19516 26688 19832 26689
rect 19516 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19832 26688
rect 19516 26623 19832 26624
rect 26944 26688 27260 26689
rect 26944 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27260 26688
rect 26944 26623 27260 26624
rect 5320 26144 5636 26145
rect 5320 26080 5326 26144
rect 5390 26080 5406 26144
rect 5470 26080 5486 26144
rect 5550 26080 5566 26144
rect 5630 26080 5636 26144
rect 5320 26079 5636 26080
rect 12748 26144 13064 26145
rect 12748 26080 12754 26144
rect 12818 26080 12834 26144
rect 12898 26080 12914 26144
rect 12978 26080 12994 26144
rect 13058 26080 13064 26144
rect 12748 26079 13064 26080
rect 20176 26144 20492 26145
rect 20176 26080 20182 26144
rect 20246 26080 20262 26144
rect 20326 26080 20342 26144
rect 20406 26080 20422 26144
rect 20486 26080 20492 26144
rect 20176 26079 20492 26080
rect 27604 26144 27920 26145
rect 27604 26080 27610 26144
rect 27674 26080 27690 26144
rect 27754 26080 27770 26144
rect 27834 26080 27850 26144
rect 27914 26080 27920 26144
rect 27604 26079 27920 26080
rect 4660 25600 4976 25601
rect 4660 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4976 25600
rect 4660 25535 4976 25536
rect 12088 25600 12404 25601
rect 12088 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12404 25600
rect 12088 25535 12404 25536
rect 19516 25600 19832 25601
rect 19516 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19832 25600
rect 19516 25535 19832 25536
rect 26944 25600 27260 25601
rect 26944 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27260 25600
rect 26944 25535 27260 25536
rect 0 25258 800 25288
rect 3417 25258 3483 25261
rect 0 25256 3483 25258
rect 0 25200 3422 25256
rect 3478 25200 3483 25256
rect 0 25198 3483 25200
rect 0 25168 800 25198
rect 3417 25195 3483 25198
rect 5320 25056 5636 25057
rect 5320 24992 5326 25056
rect 5390 24992 5406 25056
rect 5470 24992 5486 25056
rect 5550 24992 5566 25056
rect 5630 24992 5636 25056
rect 5320 24991 5636 24992
rect 12748 25056 13064 25057
rect 12748 24992 12754 25056
rect 12818 24992 12834 25056
rect 12898 24992 12914 25056
rect 12978 24992 12994 25056
rect 13058 24992 13064 25056
rect 12748 24991 13064 24992
rect 20176 25056 20492 25057
rect 20176 24992 20182 25056
rect 20246 24992 20262 25056
rect 20326 24992 20342 25056
rect 20406 24992 20422 25056
rect 20486 24992 20492 25056
rect 20176 24991 20492 24992
rect 27604 25056 27920 25057
rect 27604 24992 27610 25056
rect 27674 24992 27690 25056
rect 27754 24992 27770 25056
rect 27834 24992 27850 25056
rect 27914 24992 27920 25056
rect 27604 24991 27920 24992
rect 4660 24512 4976 24513
rect 4660 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4976 24512
rect 4660 24447 4976 24448
rect 12088 24512 12404 24513
rect 12088 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12404 24512
rect 12088 24447 12404 24448
rect 19516 24512 19832 24513
rect 19516 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19832 24512
rect 19516 24447 19832 24448
rect 26944 24512 27260 24513
rect 26944 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27260 24512
rect 26944 24447 27260 24448
rect 5320 23968 5636 23969
rect 5320 23904 5326 23968
rect 5390 23904 5406 23968
rect 5470 23904 5486 23968
rect 5550 23904 5566 23968
rect 5630 23904 5636 23968
rect 5320 23903 5636 23904
rect 12748 23968 13064 23969
rect 12748 23904 12754 23968
rect 12818 23904 12834 23968
rect 12898 23904 12914 23968
rect 12978 23904 12994 23968
rect 13058 23904 13064 23968
rect 12748 23903 13064 23904
rect 20176 23968 20492 23969
rect 20176 23904 20182 23968
rect 20246 23904 20262 23968
rect 20326 23904 20342 23968
rect 20406 23904 20422 23968
rect 20486 23904 20492 23968
rect 20176 23903 20492 23904
rect 27604 23968 27920 23969
rect 27604 23904 27610 23968
rect 27674 23904 27690 23968
rect 27754 23904 27770 23968
rect 27834 23904 27850 23968
rect 27914 23904 27920 23968
rect 27604 23903 27920 23904
rect 1485 23490 1551 23493
rect 798 23488 1551 23490
rect 798 23432 1490 23488
rect 1546 23432 1551 23488
rect 798 23430 1551 23432
rect 798 23248 858 23430
rect 1485 23427 1551 23430
rect 4660 23424 4976 23425
rect 4660 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4976 23424
rect 4660 23359 4976 23360
rect 12088 23424 12404 23425
rect 12088 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12404 23424
rect 12088 23359 12404 23360
rect 19516 23424 19832 23425
rect 19516 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19832 23424
rect 19516 23359 19832 23360
rect 26944 23424 27260 23425
rect 26944 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27260 23424
rect 26944 23359 27260 23360
rect 0 23158 858 23248
rect 30281 23218 30347 23221
rect 31200 23218 32000 23248
rect 30281 23216 32000 23218
rect 30281 23160 30286 23216
rect 30342 23160 32000 23216
rect 30281 23158 32000 23160
rect 0 23128 800 23158
rect 30281 23155 30347 23158
rect 31200 23128 32000 23158
rect 5320 22880 5636 22881
rect 5320 22816 5326 22880
rect 5390 22816 5406 22880
rect 5470 22816 5486 22880
rect 5550 22816 5566 22880
rect 5630 22816 5636 22880
rect 5320 22815 5636 22816
rect 12748 22880 13064 22881
rect 12748 22816 12754 22880
rect 12818 22816 12834 22880
rect 12898 22816 12914 22880
rect 12978 22816 12994 22880
rect 13058 22816 13064 22880
rect 12748 22815 13064 22816
rect 20176 22880 20492 22881
rect 20176 22816 20182 22880
rect 20246 22816 20262 22880
rect 20326 22816 20342 22880
rect 20406 22816 20422 22880
rect 20486 22816 20492 22880
rect 20176 22815 20492 22816
rect 27604 22880 27920 22881
rect 27604 22816 27610 22880
rect 27674 22816 27690 22880
rect 27754 22816 27770 22880
rect 27834 22816 27850 22880
rect 27914 22816 27920 22880
rect 27604 22815 27920 22816
rect 20989 22674 21055 22677
rect 22553 22674 22619 22677
rect 20989 22672 22619 22674
rect 20989 22616 20994 22672
rect 21050 22616 22558 22672
rect 22614 22616 22619 22672
rect 20989 22614 22619 22616
rect 20989 22611 21055 22614
rect 22553 22611 22619 22614
rect 0 22538 800 22568
rect 933 22538 999 22541
rect 0 22536 999 22538
rect 0 22480 938 22536
rect 994 22480 999 22536
rect 0 22478 999 22480
rect 0 22448 800 22478
rect 933 22475 999 22478
rect 22001 22538 22067 22541
rect 24025 22538 24091 22541
rect 22001 22536 24091 22538
rect 22001 22480 22006 22536
rect 22062 22480 24030 22536
rect 24086 22480 24091 22536
rect 22001 22478 24091 22480
rect 22001 22475 22067 22478
rect 24025 22475 24091 22478
rect 30925 22538 30991 22541
rect 31200 22538 32000 22568
rect 30925 22536 32000 22538
rect 30925 22480 30930 22536
rect 30986 22480 32000 22536
rect 30925 22478 32000 22480
rect 30925 22475 30991 22478
rect 31200 22448 32000 22478
rect 4660 22336 4976 22337
rect 4660 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4976 22336
rect 4660 22271 4976 22272
rect 12088 22336 12404 22337
rect 12088 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12404 22336
rect 12088 22271 12404 22272
rect 19516 22336 19832 22337
rect 19516 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19832 22336
rect 19516 22271 19832 22272
rect 26944 22336 27260 22337
rect 26944 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27260 22336
rect 26944 22271 27260 22272
rect 0 21858 800 21888
rect 933 21858 999 21861
rect 0 21856 999 21858
rect 0 21800 938 21856
rect 994 21800 999 21856
rect 0 21798 999 21800
rect 0 21768 800 21798
rect 933 21795 999 21798
rect 30465 21858 30531 21861
rect 31200 21858 32000 21888
rect 30465 21856 32000 21858
rect 30465 21800 30470 21856
rect 30526 21800 32000 21856
rect 30465 21798 32000 21800
rect 30465 21795 30531 21798
rect 5320 21792 5636 21793
rect 5320 21728 5326 21792
rect 5390 21728 5406 21792
rect 5470 21728 5486 21792
rect 5550 21728 5566 21792
rect 5630 21728 5636 21792
rect 5320 21727 5636 21728
rect 12748 21792 13064 21793
rect 12748 21728 12754 21792
rect 12818 21728 12834 21792
rect 12898 21728 12914 21792
rect 12978 21728 12994 21792
rect 13058 21728 13064 21792
rect 12748 21727 13064 21728
rect 20176 21792 20492 21793
rect 20176 21728 20182 21792
rect 20246 21728 20262 21792
rect 20326 21728 20342 21792
rect 20406 21728 20422 21792
rect 20486 21728 20492 21792
rect 20176 21727 20492 21728
rect 27604 21792 27920 21793
rect 27604 21728 27610 21792
rect 27674 21728 27690 21792
rect 27754 21728 27770 21792
rect 27834 21728 27850 21792
rect 27914 21728 27920 21792
rect 31200 21768 32000 21798
rect 27604 21727 27920 21728
rect 4660 21248 4976 21249
rect 0 21178 800 21208
rect 4660 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4976 21248
rect 4660 21183 4976 21184
rect 12088 21248 12404 21249
rect 12088 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12404 21248
rect 12088 21183 12404 21184
rect 19516 21248 19832 21249
rect 19516 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19832 21248
rect 19516 21183 19832 21184
rect 26944 21248 27260 21249
rect 26944 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27260 21248
rect 26944 21183 27260 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 30373 21178 30439 21181
rect 31200 21178 32000 21208
rect 30373 21176 32000 21178
rect 30373 21120 30378 21176
rect 30434 21120 32000 21176
rect 30373 21118 32000 21120
rect 30373 21115 30439 21118
rect 31200 21088 32000 21118
rect 5320 20704 5636 20705
rect 5320 20640 5326 20704
rect 5390 20640 5406 20704
rect 5470 20640 5486 20704
rect 5550 20640 5566 20704
rect 5630 20640 5636 20704
rect 5320 20639 5636 20640
rect 12748 20704 13064 20705
rect 12748 20640 12754 20704
rect 12818 20640 12834 20704
rect 12898 20640 12914 20704
rect 12978 20640 12994 20704
rect 13058 20640 13064 20704
rect 12748 20639 13064 20640
rect 20176 20704 20492 20705
rect 20176 20640 20182 20704
rect 20246 20640 20262 20704
rect 20326 20640 20342 20704
rect 20406 20640 20422 20704
rect 20486 20640 20492 20704
rect 20176 20639 20492 20640
rect 27604 20704 27920 20705
rect 27604 20640 27610 20704
rect 27674 20640 27690 20704
rect 27754 20640 27770 20704
rect 27834 20640 27850 20704
rect 27914 20640 27920 20704
rect 27604 20639 27920 20640
rect 1485 20634 1551 20637
rect 798 20632 1551 20634
rect 798 20576 1490 20632
rect 1546 20576 1551 20632
rect 798 20574 1551 20576
rect 798 20528 858 20574
rect 1485 20571 1551 20574
rect 0 20438 858 20528
rect 30281 20498 30347 20501
rect 31200 20498 32000 20528
rect 30281 20496 32000 20498
rect 30281 20440 30286 20496
rect 30342 20440 32000 20496
rect 30281 20438 32000 20440
rect 0 20408 800 20438
rect 30281 20435 30347 20438
rect 31200 20408 32000 20438
rect 4660 20160 4976 20161
rect 4660 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4976 20160
rect 4660 20095 4976 20096
rect 12088 20160 12404 20161
rect 12088 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12404 20160
rect 12088 20095 12404 20096
rect 19516 20160 19832 20161
rect 19516 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19832 20160
rect 19516 20095 19832 20096
rect 26944 20160 27260 20161
rect 26944 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27260 20160
rect 26944 20095 27260 20096
rect 0 19818 800 19848
rect 933 19818 999 19821
rect 0 19816 999 19818
rect 0 19760 938 19816
rect 994 19760 999 19816
rect 0 19758 999 19760
rect 0 19728 800 19758
rect 933 19755 999 19758
rect 30373 19818 30439 19821
rect 31200 19818 32000 19848
rect 30373 19816 32000 19818
rect 30373 19760 30378 19816
rect 30434 19760 32000 19816
rect 30373 19758 32000 19760
rect 30373 19755 30439 19758
rect 31200 19728 32000 19758
rect 5320 19616 5636 19617
rect 5320 19552 5326 19616
rect 5390 19552 5406 19616
rect 5470 19552 5486 19616
rect 5550 19552 5566 19616
rect 5630 19552 5636 19616
rect 5320 19551 5636 19552
rect 12748 19616 13064 19617
rect 12748 19552 12754 19616
rect 12818 19552 12834 19616
rect 12898 19552 12914 19616
rect 12978 19552 12994 19616
rect 13058 19552 13064 19616
rect 12748 19551 13064 19552
rect 20176 19616 20492 19617
rect 20176 19552 20182 19616
rect 20246 19552 20262 19616
rect 20326 19552 20342 19616
rect 20406 19552 20422 19616
rect 20486 19552 20492 19616
rect 20176 19551 20492 19552
rect 27604 19616 27920 19617
rect 27604 19552 27610 19616
rect 27674 19552 27690 19616
rect 27754 19552 27770 19616
rect 27834 19552 27850 19616
rect 27914 19552 27920 19616
rect 27604 19551 27920 19552
rect 1393 19274 1459 19277
rect 798 19272 1459 19274
rect 798 19216 1398 19272
rect 1454 19216 1459 19272
rect 798 19214 1459 19216
rect 798 19168 858 19214
rect 1393 19211 1459 19214
rect 0 19078 858 19168
rect 30281 19138 30347 19141
rect 31200 19138 32000 19168
rect 30281 19136 32000 19138
rect 30281 19080 30286 19136
rect 30342 19080 32000 19136
rect 30281 19078 32000 19080
rect 0 19048 800 19078
rect 30281 19075 30347 19078
rect 4660 19072 4976 19073
rect 4660 19008 4666 19072
rect 4730 19008 4746 19072
rect 4810 19008 4826 19072
rect 4890 19008 4906 19072
rect 4970 19008 4976 19072
rect 4660 19007 4976 19008
rect 12088 19072 12404 19073
rect 12088 19008 12094 19072
rect 12158 19008 12174 19072
rect 12238 19008 12254 19072
rect 12318 19008 12334 19072
rect 12398 19008 12404 19072
rect 12088 19007 12404 19008
rect 19516 19072 19832 19073
rect 19516 19008 19522 19072
rect 19586 19008 19602 19072
rect 19666 19008 19682 19072
rect 19746 19008 19762 19072
rect 19826 19008 19832 19072
rect 19516 19007 19832 19008
rect 26944 19072 27260 19073
rect 26944 19008 26950 19072
rect 27014 19008 27030 19072
rect 27094 19008 27110 19072
rect 27174 19008 27190 19072
rect 27254 19008 27260 19072
rect 31200 19048 32000 19078
rect 26944 19007 27260 19008
rect 5320 18528 5636 18529
rect 0 18458 800 18488
rect 5320 18464 5326 18528
rect 5390 18464 5406 18528
rect 5470 18464 5486 18528
rect 5550 18464 5566 18528
rect 5630 18464 5636 18528
rect 5320 18463 5636 18464
rect 12748 18528 13064 18529
rect 12748 18464 12754 18528
rect 12818 18464 12834 18528
rect 12898 18464 12914 18528
rect 12978 18464 12994 18528
rect 13058 18464 13064 18528
rect 12748 18463 13064 18464
rect 20176 18528 20492 18529
rect 20176 18464 20182 18528
rect 20246 18464 20262 18528
rect 20326 18464 20342 18528
rect 20406 18464 20422 18528
rect 20486 18464 20492 18528
rect 20176 18463 20492 18464
rect 27604 18528 27920 18529
rect 27604 18464 27610 18528
rect 27674 18464 27690 18528
rect 27754 18464 27770 18528
rect 27834 18464 27850 18528
rect 27914 18464 27920 18528
rect 27604 18463 27920 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 30373 18458 30439 18461
rect 31200 18458 32000 18488
rect 30373 18456 32000 18458
rect 30373 18400 30378 18456
rect 30434 18400 32000 18456
rect 30373 18398 32000 18400
rect 30373 18395 30439 18398
rect 31200 18368 32000 18398
rect 11973 18322 12039 18325
rect 17585 18322 17651 18325
rect 11973 18320 17651 18322
rect 11973 18264 11978 18320
rect 12034 18264 17590 18320
rect 17646 18264 17651 18320
rect 11973 18262 17651 18264
rect 11973 18259 12039 18262
rect 17585 18259 17651 18262
rect 4660 17984 4976 17985
rect 4660 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4976 17984
rect 4660 17919 4976 17920
rect 12088 17984 12404 17985
rect 12088 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12404 17984
rect 12088 17919 12404 17920
rect 19516 17984 19832 17985
rect 19516 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19832 17984
rect 19516 17919 19832 17920
rect 26944 17984 27260 17985
rect 26944 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27260 17984
rect 26944 17919 27260 17920
rect 1485 17914 1551 17917
rect 798 17912 1551 17914
rect 798 17856 1490 17912
rect 1546 17856 1551 17912
rect 798 17854 1551 17856
rect 798 17808 858 17854
rect 1485 17851 1551 17854
rect 0 17718 858 17808
rect 30281 17778 30347 17781
rect 31200 17778 32000 17808
rect 30281 17776 32000 17778
rect 30281 17720 30286 17776
rect 30342 17720 32000 17776
rect 30281 17718 32000 17720
rect 0 17688 800 17718
rect 30281 17715 30347 17718
rect 31200 17688 32000 17718
rect 5320 17440 5636 17441
rect 5320 17376 5326 17440
rect 5390 17376 5406 17440
rect 5470 17376 5486 17440
rect 5550 17376 5566 17440
rect 5630 17376 5636 17440
rect 5320 17375 5636 17376
rect 12748 17440 13064 17441
rect 12748 17376 12754 17440
rect 12818 17376 12834 17440
rect 12898 17376 12914 17440
rect 12978 17376 12994 17440
rect 13058 17376 13064 17440
rect 12748 17375 13064 17376
rect 20176 17440 20492 17441
rect 20176 17376 20182 17440
rect 20246 17376 20262 17440
rect 20326 17376 20342 17440
rect 20406 17376 20422 17440
rect 20486 17376 20492 17440
rect 20176 17375 20492 17376
rect 27604 17440 27920 17441
rect 27604 17376 27610 17440
rect 27674 17376 27690 17440
rect 27754 17376 27770 17440
rect 27834 17376 27850 17440
rect 27914 17376 27920 17440
rect 27604 17375 27920 17376
rect 5717 17234 5783 17237
rect 6269 17234 6335 17237
rect 5717 17232 6335 17234
rect 5717 17176 5722 17232
rect 5778 17176 6274 17232
rect 6330 17176 6335 17232
rect 5717 17174 6335 17176
rect 5717 17171 5783 17174
rect 6269 17171 6335 17174
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 30373 17098 30439 17101
rect 31200 17098 32000 17128
rect 30373 17096 32000 17098
rect 30373 17040 30378 17096
rect 30434 17040 32000 17096
rect 30373 17038 32000 17040
rect 30373 17035 30439 17038
rect 31200 17008 32000 17038
rect 4660 16896 4976 16897
rect 4660 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4976 16896
rect 4660 16831 4976 16832
rect 12088 16896 12404 16897
rect 12088 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12404 16896
rect 12088 16831 12404 16832
rect 19516 16896 19832 16897
rect 19516 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19832 16896
rect 19516 16831 19832 16832
rect 26944 16896 27260 16897
rect 26944 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27260 16896
rect 26944 16831 27260 16832
rect 10501 16554 10567 16557
rect 14273 16554 14339 16557
rect 10501 16552 14339 16554
rect 10501 16496 10506 16552
rect 10562 16496 14278 16552
rect 14334 16496 14339 16552
rect 10501 16494 14339 16496
rect 10501 16491 10567 16494
rect 14273 16491 14339 16494
rect 20805 16554 20871 16557
rect 23657 16554 23723 16557
rect 20805 16552 23723 16554
rect 20805 16496 20810 16552
rect 20866 16496 23662 16552
rect 23718 16496 23723 16552
rect 20805 16494 23723 16496
rect 20805 16491 20871 16494
rect 23657 16491 23723 16494
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 30925 16418 30991 16421
rect 31200 16418 32000 16448
rect 30925 16416 32000 16418
rect 30925 16360 30930 16416
rect 30986 16360 32000 16416
rect 30925 16358 32000 16360
rect 30925 16355 30991 16358
rect 5320 16352 5636 16353
rect 5320 16288 5326 16352
rect 5390 16288 5406 16352
rect 5470 16288 5486 16352
rect 5550 16288 5566 16352
rect 5630 16288 5636 16352
rect 5320 16287 5636 16288
rect 12748 16352 13064 16353
rect 12748 16288 12754 16352
rect 12818 16288 12834 16352
rect 12898 16288 12914 16352
rect 12978 16288 12994 16352
rect 13058 16288 13064 16352
rect 12748 16287 13064 16288
rect 20176 16352 20492 16353
rect 20176 16288 20182 16352
rect 20246 16288 20262 16352
rect 20326 16288 20342 16352
rect 20406 16288 20422 16352
rect 20486 16288 20492 16352
rect 20176 16287 20492 16288
rect 27604 16352 27920 16353
rect 27604 16288 27610 16352
rect 27674 16288 27690 16352
rect 27754 16288 27770 16352
rect 27834 16288 27850 16352
rect 27914 16288 27920 16352
rect 31200 16328 32000 16358
rect 27604 16287 27920 16288
rect 4660 15808 4976 15809
rect 0 15738 800 15768
rect 4660 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4976 15808
rect 4660 15743 4976 15744
rect 12088 15808 12404 15809
rect 12088 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12404 15808
rect 12088 15743 12404 15744
rect 19516 15808 19832 15809
rect 19516 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19832 15808
rect 19516 15743 19832 15744
rect 26944 15808 27260 15809
rect 26944 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27260 15808
rect 26944 15743 27260 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 30373 15738 30439 15741
rect 31200 15738 32000 15768
rect 30373 15736 32000 15738
rect 30373 15680 30378 15736
rect 30434 15680 32000 15736
rect 30373 15678 32000 15680
rect 30373 15675 30439 15678
rect 31200 15648 32000 15678
rect 5320 15264 5636 15265
rect 5320 15200 5326 15264
rect 5390 15200 5406 15264
rect 5470 15200 5486 15264
rect 5550 15200 5566 15264
rect 5630 15200 5636 15264
rect 5320 15199 5636 15200
rect 12748 15264 13064 15265
rect 12748 15200 12754 15264
rect 12818 15200 12834 15264
rect 12898 15200 12914 15264
rect 12978 15200 12994 15264
rect 13058 15200 13064 15264
rect 12748 15199 13064 15200
rect 20176 15264 20492 15265
rect 20176 15200 20182 15264
rect 20246 15200 20262 15264
rect 20326 15200 20342 15264
rect 20406 15200 20422 15264
rect 20486 15200 20492 15264
rect 20176 15199 20492 15200
rect 27604 15264 27920 15265
rect 27604 15200 27610 15264
rect 27674 15200 27690 15264
rect 27754 15200 27770 15264
rect 27834 15200 27850 15264
rect 27914 15200 27920 15264
rect 27604 15199 27920 15200
rect 1393 15192 1459 15197
rect 1393 15136 1398 15192
rect 1454 15136 1459 15192
rect 1393 15131 1459 15136
rect 0 15058 800 15088
rect 1396 15058 1456 15131
rect 0 14998 1456 15058
rect 30281 15058 30347 15061
rect 31200 15058 32000 15088
rect 30281 15056 32000 15058
rect 30281 15000 30286 15056
rect 30342 15000 32000 15056
rect 30281 14998 32000 15000
rect 0 14968 800 14998
rect 30281 14995 30347 14998
rect 31200 14968 32000 14998
rect 4660 14720 4976 14721
rect 4660 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4976 14720
rect 4660 14655 4976 14656
rect 12088 14720 12404 14721
rect 12088 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12404 14720
rect 12088 14655 12404 14656
rect 19516 14720 19832 14721
rect 19516 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19832 14720
rect 19516 14655 19832 14656
rect 26944 14720 27260 14721
rect 26944 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27260 14720
rect 26944 14655 27260 14656
rect 0 14378 800 14408
rect 933 14378 999 14381
rect 0 14376 999 14378
rect 0 14320 938 14376
rect 994 14320 999 14376
rect 0 14318 999 14320
rect 0 14288 800 14318
rect 933 14315 999 14318
rect 16481 14378 16547 14381
rect 21449 14378 21515 14381
rect 16481 14376 21515 14378
rect 16481 14320 16486 14376
rect 16542 14320 21454 14376
rect 21510 14320 21515 14376
rect 16481 14318 21515 14320
rect 16481 14315 16547 14318
rect 21449 14315 21515 14318
rect 30373 14378 30439 14381
rect 31200 14378 32000 14408
rect 30373 14376 32000 14378
rect 30373 14320 30378 14376
rect 30434 14320 32000 14376
rect 30373 14318 32000 14320
rect 30373 14315 30439 14318
rect 31200 14288 32000 14318
rect 5320 14176 5636 14177
rect 5320 14112 5326 14176
rect 5390 14112 5406 14176
rect 5470 14112 5486 14176
rect 5550 14112 5566 14176
rect 5630 14112 5636 14176
rect 5320 14111 5636 14112
rect 12748 14176 13064 14177
rect 12748 14112 12754 14176
rect 12818 14112 12834 14176
rect 12898 14112 12914 14176
rect 12978 14112 12994 14176
rect 13058 14112 13064 14176
rect 12748 14111 13064 14112
rect 20176 14176 20492 14177
rect 20176 14112 20182 14176
rect 20246 14112 20262 14176
rect 20326 14112 20342 14176
rect 20406 14112 20422 14176
rect 20486 14112 20492 14176
rect 20176 14111 20492 14112
rect 27604 14176 27920 14177
rect 27604 14112 27610 14176
rect 27674 14112 27690 14176
rect 27754 14112 27770 14176
rect 27834 14112 27850 14176
rect 27914 14112 27920 14176
rect 27604 14111 27920 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 30281 13698 30347 13701
rect 31200 13698 32000 13728
rect 30281 13696 32000 13698
rect 30281 13640 30286 13696
rect 30342 13640 32000 13696
rect 30281 13638 32000 13640
rect 30281 13635 30347 13638
rect 4660 13632 4976 13633
rect 4660 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4976 13632
rect 4660 13567 4976 13568
rect 12088 13632 12404 13633
rect 12088 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12404 13632
rect 12088 13567 12404 13568
rect 19516 13632 19832 13633
rect 19516 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19832 13632
rect 19516 13567 19832 13568
rect 26944 13632 27260 13633
rect 26944 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27260 13632
rect 31200 13608 32000 13638
rect 26944 13567 27260 13568
rect 5320 13088 5636 13089
rect 0 13018 800 13048
rect 5320 13024 5326 13088
rect 5390 13024 5406 13088
rect 5470 13024 5486 13088
rect 5550 13024 5566 13088
rect 5630 13024 5636 13088
rect 5320 13023 5636 13024
rect 12748 13088 13064 13089
rect 12748 13024 12754 13088
rect 12818 13024 12834 13088
rect 12898 13024 12914 13088
rect 12978 13024 12994 13088
rect 13058 13024 13064 13088
rect 12748 13023 13064 13024
rect 20176 13088 20492 13089
rect 20176 13024 20182 13088
rect 20246 13024 20262 13088
rect 20326 13024 20342 13088
rect 20406 13024 20422 13088
rect 20486 13024 20492 13088
rect 20176 13023 20492 13024
rect 27604 13088 27920 13089
rect 27604 13024 27610 13088
rect 27674 13024 27690 13088
rect 27754 13024 27770 13088
rect 27834 13024 27850 13088
rect 27914 13024 27920 13088
rect 27604 13023 27920 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 30373 13018 30439 13021
rect 31200 13018 32000 13048
rect 30373 13016 32000 13018
rect 30373 12960 30378 13016
rect 30434 12960 32000 13016
rect 30373 12958 32000 12960
rect 30373 12955 30439 12958
rect 31200 12928 32000 12958
rect 11053 12746 11119 12749
rect 16297 12746 16363 12749
rect 11053 12744 16363 12746
rect 11053 12688 11058 12744
rect 11114 12688 16302 12744
rect 16358 12688 16363 12744
rect 11053 12686 16363 12688
rect 11053 12683 11119 12686
rect 16297 12683 16363 12686
rect 4660 12544 4976 12545
rect 4660 12480 4666 12544
rect 4730 12480 4746 12544
rect 4810 12480 4826 12544
rect 4890 12480 4906 12544
rect 4970 12480 4976 12544
rect 4660 12479 4976 12480
rect 12088 12544 12404 12545
rect 12088 12480 12094 12544
rect 12158 12480 12174 12544
rect 12238 12480 12254 12544
rect 12318 12480 12334 12544
rect 12398 12480 12404 12544
rect 12088 12479 12404 12480
rect 19516 12544 19832 12545
rect 19516 12480 19522 12544
rect 19586 12480 19602 12544
rect 19666 12480 19682 12544
rect 19746 12480 19762 12544
rect 19826 12480 19832 12544
rect 19516 12479 19832 12480
rect 26944 12544 27260 12545
rect 26944 12480 26950 12544
rect 27014 12480 27030 12544
rect 27094 12480 27110 12544
rect 27174 12480 27190 12544
rect 27254 12480 27260 12544
rect 26944 12479 27260 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 14917 12338 14983 12341
rect 18229 12338 18295 12341
rect 14917 12336 18295 12338
rect 14917 12280 14922 12336
rect 14978 12280 18234 12336
rect 18290 12280 18295 12336
rect 14917 12278 18295 12280
rect 14917 12275 14983 12278
rect 18229 12275 18295 12278
rect 30281 12338 30347 12341
rect 31200 12338 32000 12368
rect 30281 12336 32000 12338
rect 30281 12280 30286 12336
rect 30342 12280 32000 12336
rect 30281 12278 32000 12280
rect 30281 12275 30347 12278
rect 31200 12248 32000 12278
rect 20437 12202 20503 12205
rect 21265 12202 21331 12205
rect 20437 12200 21331 12202
rect 20437 12144 20442 12200
rect 20498 12144 21270 12200
rect 21326 12144 21331 12200
rect 20437 12142 21331 12144
rect 20437 12139 20503 12142
rect 21265 12139 21331 12142
rect 5320 12000 5636 12001
rect 5320 11936 5326 12000
rect 5390 11936 5406 12000
rect 5470 11936 5486 12000
rect 5550 11936 5566 12000
rect 5630 11936 5636 12000
rect 5320 11935 5636 11936
rect 12748 12000 13064 12001
rect 12748 11936 12754 12000
rect 12818 11936 12834 12000
rect 12898 11936 12914 12000
rect 12978 11936 12994 12000
rect 13058 11936 13064 12000
rect 12748 11935 13064 11936
rect 20176 12000 20492 12001
rect 20176 11936 20182 12000
rect 20246 11936 20262 12000
rect 20326 11936 20342 12000
rect 20406 11936 20422 12000
rect 20486 11936 20492 12000
rect 20176 11935 20492 11936
rect 27604 12000 27920 12001
rect 27604 11936 27610 12000
rect 27674 11936 27690 12000
rect 27754 11936 27770 12000
rect 27834 11936 27850 12000
rect 27914 11936 27920 12000
rect 27604 11935 27920 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 30373 11658 30439 11661
rect 31200 11658 32000 11688
rect 30373 11656 32000 11658
rect 30373 11600 30378 11656
rect 30434 11600 32000 11656
rect 30373 11598 32000 11600
rect 30373 11595 30439 11598
rect 31200 11568 32000 11598
rect 4660 11456 4976 11457
rect 4660 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4976 11456
rect 4660 11391 4976 11392
rect 12088 11456 12404 11457
rect 12088 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12404 11456
rect 12088 11391 12404 11392
rect 19516 11456 19832 11457
rect 19516 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19832 11456
rect 19516 11391 19832 11392
rect 26944 11456 27260 11457
rect 26944 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27260 11456
rect 26944 11391 27260 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 30281 10978 30347 10981
rect 31200 10978 32000 11008
rect 30281 10976 32000 10978
rect 30281 10920 30286 10976
rect 30342 10920 32000 10976
rect 30281 10918 32000 10920
rect 30281 10915 30347 10918
rect 5320 10912 5636 10913
rect 5320 10848 5326 10912
rect 5390 10848 5406 10912
rect 5470 10848 5486 10912
rect 5550 10848 5566 10912
rect 5630 10848 5636 10912
rect 5320 10847 5636 10848
rect 12748 10912 13064 10913
rect 12748 10848 12754 10912
rect 12818 10848 12834 10912
rect 12898 10848 12914 10912
rect 12978 10848 12994 10912
rect 13058 10848 13064 10912
rect 12748 10847 13064 10848
rect 20176 10912 20492 10913
rect 20176 10848 20182 10912
rect 20246 10848 20262 10912
rect 20326 10848 20342 10912
rect 20406 10848 20422 10912
rect 20486 10848 20492 10912
rect 20176 10847 20492 10848
rect 27604 10912 27920 10913
rect 27604 10848 27610 10912
rect 27674 10848 27690 10912
rect 27754 10848 27770 10912
rect 27834 10848 27850 10912
rect 27914 10848 27920 10912
rect 31200 10888 32000 10918
rect 27604 10847 27920 10848
rect 4660 10368 4976 10369
rect 0 10298 800 10328
rect 4660 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4976 10368
rect 4660 10303 4976 10304
rect 12088 10368 12404 10369
rect 12088 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12404 10368
rect 12088 10303 12404 10304
rect 19516 10368 19832 10369
rect 19516 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19832 10368
rect 19516 10303 19832 10304
rect 26944 10368 27260 10369
rect 26944 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27260 10368
rect 26944 10303 27260 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 30925 10298 30991 10301
rect 31200 10298 32000 10328
rect 30925 10296 32000 10298
rect 30925 10240 30930 10296
rect 30986 10240 32000 10296
rect 30925 10238 32000 10240
rect 30925 10235 30991 10238
rect 31200 10208 32000 10238
rect 19793 10162 19859 10165
rect 20161 10162 20227 10165
rect 19793 10160 20227 10162
rect 19793 10104 19798 10160
rect 19854 10104 20166 10160
rect 20222 10104 20227 10160
rect 19793 10102 20227 10104
rect 19793 10099 19859 10102
rect 20161 10099 20227 10102
rect 5320 9824 5636 9825
rect 5320 9760 5326 9824
rect 5390 9760 5406 9824
rect 5470 9760 5486 9824
rect 5550 9760 5566 9824
rect 5630 9760 5636 9824
rect 5320 9759 5636 9760
rect 12748 9824 13064 9825
rect 12748 9760 12754 9824
rect 12818 9760 12834 9824
rect 12898 9760 12914 9824
rect 12978 9760 12994 9824
rect 13058 9760 13064 9824
rect 12748 9759 13064 9760
rect 20176 9824 20492 9825
rect 20176 9760 20182 9824
rect 20246 9760 20262 9824
rect 20326 9760 20342 9824
rect 20406 9760 20422 9824
rect 20486 9760 20492 9824
rect 20176 9759 20492 9760
rect 27604 9824 27920 9825
rect 27604 9760 27610 9824
rect 27674 9760 27690 9824
rect 27754 9760 27770 9824
rect 27834 9760 27850 9824
rect 27914 9760 27920 9824
rect 27604 9759 27920 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 30281 9618 30347 9621
rect 31200 9618 32000 9648
rect 30281 9616 32000 9618
rect 30281 9560 30286 9616
rect 30342 9560 32000 9616
rect 30281 9558 32000 9560
rect 30281 9555 30347 9558
rect 31200 9528 32000 9558
rect 20529 9482 20595 9485
rect 25313 9482 25379 9485
rect 20529 9480 25379 9482
rect 20529 9424 20534 9480
rect 20590 9424 25318 9480
rect 25374 9424 25379 9480
rect 20529 9422 25379 9424
rect 20529 9419 20595 9422
rect 25313 9419 25379 9422
rect 4660 9280 4976 9281
rect 4660 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4976 9280
rect 4660 9215 4976 9216
rect 12088 9280 12404 9281
rect 12088 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12404 9280
rect 12088 9215 12404 9216
rect 19516 9280 19832 9281
rect 19516 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19832 9280
rect 19516 9215 19832 9216
rect 26944 9280 27260 9281
rect 26944 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27260 9280
rect 26944 9215 27260 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 30373 8938 30439 8941
rect 31200 8938 32000 8968
rect 30373 8936 32000 8938
rect 30373 8880 30378 8936
rect 30434 8880 32000 8936
rect 30373 8878 32000 8880
rect 30373 8875 30439 8878
rect 31200 8848 32000 8878
rect 5993 8802 6059 8805
rect 9489 8802 9555 8805
rect 5993 8800 9555 8802
rect 5993 8744 5998 8800
rect 6054 8744 9494 8800
rect 9550 8744 9555 8800
rect 5993 8742 9555 8744
rect 5993 8739 6059 8742
rect 9489 8739 9555 8742
rect 5320 8736 5636 8737
rect 5320 8672 5326 8736
rect 5390 8672 5406 8736
rect 5470 8672 5486 8736
rect 5550 8672 5566 8736
rect 5630 8672 5636 8736
rect 5320 8671 5636 8672
rect 12748 8736 13064 8737
rect 12748 8672 12754 8736
rect 12818 8672 12834 8736
rect 12898 8672 12914 8736
rect 12978 8672 12994 8736
rect 13058 8672 13064 8736
rect 12748 8671 13064 8672
rect 20176 8736 20492 8737
rect 20176 8672 20182 8736
rect 20246 8672 20262 8736
rect 20326 8672 20342 8736
rect 20406 8672 20422 8736
rect 20486 8672 20492 8736
rect 20176 8671 20492 8672
rect 27604 8736 27920 8737
rect 27604 8672 27610 8736
rect 27674 8672 27690 8736
rect 27754 8672 27770 8736
rect 27834 8672 27850 8736
rect 27914 8672 27920 8736
rect 27604 8671 27920 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 30281 8258 30347 8261
rect 31200 8258 32000 8288
rect 30281 8256 32000 8258
rect 30281 8200 30286 8256
rect 30342 8200 32000 8256
rect 30281 8198 32000 8200
rect 30281 8195 30347 8198
rect 4660 8192 4976 8193
rect 4660 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4976 8192
rect 4660 8127 4976 8128
rect 12088 8192 12404 8193
rect 12088 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12404 8192
rect 12088 8127 12404 8128
rect 19516 8192 19832 8193
rect 19516 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19832 8192
rect 19516 8127 19832 8128
rect 26944 8192 27260 8193
rect 26944 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27260 8192
rect 31200 8168 32000 8198
rect 26944 8127 27260 8128
rect 5320 7648 5636 7649
rect 0 7578 800 7608
rect 5320 7584 5326 7648
rect 5390 7584 5406 7648
rect 5470 7584 5486 7648
rect 5550 7584 5566 7648
rect 5630 7584 5636 7648
rect 5320 7583 5636 7584
rect 12748 7648 13064 7649
rect 12748 7584 12754 7648
rect 12818 7584 12834 7648
rect 12898 7584 12914 7648
rect 12978 7584 12994 7648
rect 13058 7584 13064 7648
rect 12748 7583 13064 7584
rect 20176 7648 20492 7649
rect 20176 7584 20182 7648
rect 20246 7584 20262 7648
rect 20326 7584 20342 7648
rect 20406 7584 20422 7648
rect 20486 7584 20492 7648
rect 20176 7583 20492 7584
rect 27604 7648 27920 7649
rect 27604 7584 27610 7648
rect 27674 7584 27690 7648
rect 27754 7584 27770 7648
rect 27834 7584 27850 7648
rect 27914 7584 27920 7648
rect 27604 7583 27920 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 4660 7104 4976 7105
rect 4660 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4976 7104
rect 4660 7039 4976 7040
rect 12088 7104 12404 7105
rect 12088 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12404 7104
rect 12088 7039 12404 7040
rect 19516 7104 19832 7105
rect 19516 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19832 7104
rect 19516 7039 19832 7040
rect 26944 7104 27260 7105
rect 26944 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27260 7104
rect 26944 7039 27260 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 5320 6560 5636 6561
rect 5320 6496 5326 6560
rect 5390 6496 5406 6560
rect 5470 6496 5486 6560
rect 5550 6496 5566 6560
rect 5630 6496 5636 6560
rect 5320 6495 5636 6496
rect 12748 6560 13064 6561
rect 12748 6496 12754 6560
rect 12818 6496 12834 6560
rect 12898 6496 12914 6560
rect 12978 6496 12994 6560
rect 13058 6496 13064 6560
rect 12748 6495 13064 6496
rect 20176 6560 20492 6561
rect 20176 6496 20182 6560
rect 20246 6496 20262 6560
rect 20326 6496 20342 6560
rect 20406 6496 20422 6560
rect 20486 6496 20492 6560
rect 20176 6495 20492 6496
rect 27604 6560 27920 6561
rect 27604 6496 27610 6560
rect 27674 6496 27690 6560
rect 27754 6496 27770 6560
rect 27834 6496 27850 6560
rect 27914 6496 27920 6560
rect 27604 6495 27920 6496
rect 4660 6016 4976 6017
rect 4660 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4976 6016
rect 4660 5951 4976 5952
rect 12088 6016 12404 6017
rect 12088 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12404 6016
rect 12088 5951 12404 5952
rect 19516 6016 19832 6017
rect 19516 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19832 6016
rect 19516 5951 19832 5952
rect 26944 6016 27260 6017
rect 26944 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27260 6016
rect 26944 5951 27260 5952
rect 5320 5472 5636 5473
rect 5320 5408 5326 5472
rect 5390 5408 5406 5472
rect 5470 5408 5486 5472
rect 5550 5408 5566 5472
rect 5630 5408 5636 5472
rect 5320 5407 5636 5408
rect 12748 5472 13064 5473
rect 12748 5408 12754 5472
rect 12818 5408 12834 5472
rect 12898 5408 12914 5472
rect 12978 5408 12994 5472
rect 13058 5408 13064 5472
rect 12748 5407 13064 5408
rect 20176 5472 20492 5473
rect 20176 5408 20182 5472
rect 20246 5408 20262 5472
rect 20326 5408 20342 5472
rect 20406 5408 20422 5472
rect 20486 5408 20492 5472
rect 20176 5407 20492 5408
rect 27604 5472 27920 5473
rect 27604 5408 27610 5472
rect 27674 5408 27690 5472
rect 27754 5408 27770 5472
rect 27834 5408 27850 5472
rect 27914 5408 27920 5472
rect 27604 5407 27920 5408
rect 4660 4928 4976 4929
rect 4660 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4976 4928
rect 4660 4863 4976 4864
rect 12088 4928 12404 4929
rect 12088 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12404 4928
rect 12088 4863 12404 4864
rect 19516 4928 19832 4929
rect 19516 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19832 4928
rect 19516 4863 19832 4864
rect 26944 4928 27260 4929
rect 26944 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27260 4928
rect 26944 4863 27260 4864
rect 5320 4384 5636 4385
rect 5320 4320 5326 4384
rect 5390 4320 5406 4384
rect 5470 4320 5486 4384
rect 5550 4320 5566 4384
rect 5630 4320 5636 4384
rect 5320 4319 5636 4320
rect 12748 4384 13064 4385
rect 12748 4320 12754 4384
rect 12818 4320 12834 4384
rect 12898 4320 12914 4384
rect 12978 4320 12994 4384
rect 13058 4320 13064 4384
rect 12748 4319 13064 4320
rect 20176 4384 20492 4385
rect 20176 4320 20182 4384
rect 20246 4320 20262 4384
rect 20326 4320 20342 4384
rect 20406 4320 20422 4384
rect 20486 4320 20492 4384
rect 20176 4319 20492 4320
rect 27604 4384 27920 4385
rect 27604 4320 27610 4384
rect 27674 4320 27690 4384
rect 27754 4320 27770 4384
rect 27834 4320 27850 4384
rect 27914 4320 27920 4384
rect 27604 4319 27920 4320
rect 4660 3840 4976 3841
rect 4660 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4976 3840
rect 4660 3775 4976 3776
rect 12088 3840 12404 3841
rect 12088 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12404 3840
rect 12088 3775 12404 3776
rect 19516 3840 19832 3841
rect 19516 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19832 3840
rect 19516 3775 19832 3776
rect 26944 3840 27260 3841
rect 26944 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27260 3840
rect 26944 3775 27260 3776
rect 5320 3296 5636 3297
rect 5320 3232 5326 3296
rect 5390 3232 5406 3296
rect 5470 3232 5486 3296
rect 5550 3232 5566 3296
rect 5630 3232 5636 3296
rect 5320 3231 5636 3232
rect 12748 3296 13064 3297
rect 12748 3232 12754 3296
rect 12818 3232 12834 3296
rect 12898 3232 12914 3296
rect 12978 3232 12994 3296
rect 13058 3232 13064 3296
rect 12748 3231 13064 3232
rect 20176 3296 20492 3297
rect 20176 3232 20182 3296
rect 20246 3232 20262 3296
rect 20326 3232 20342 3296
rect 20406 3232 20422 3296
rect 20486 3232 20492 3296
rect 20176 3231 20492 3232
rect 27604 3296 27920 3297
rect 27604 3232 27610 3296
rect 27674 3232 27690 3296
rect 27754 3232 27770 3296
rect 27834 3232 27850 3296
rect 27914 3232 27920 3296
rect 27604 3231 27920 3232
rect 4660 2752 4976 2753
rect 4660 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4976 2752
rect 4660 2687 4976 2688
rect 12088 2752 12404 2753
rect 12088 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12404 2752
rect 12088 2687 12404 2688
rect 19516 2752 19832 2753
rect 19516 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19832 2752
rect 19516 2687 19832 2688
rect 26944 2752 27260 2753
rect 26944 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27260 2752
rect 26944 2687 27260 2688
rect 5320 2208 5636 2209
rect 5320 2144 5326 2208
rect 5390 2144 5406 2208
rect 5470 2144 5486 2208
rect 5550 2144 5566 2208
rect 5630 2144 5636 2208
rect 5320 2143 5636 2144
rect 12748 2208 13064 2209
rect 12748 2144 12754 2208
rect 12818 2144 12834 2208
rect 12898 2144 12914 2208
rect 12978 2144 12994 2208
rect 13058 2144 13064 2208
rect 12748 2143 13064 2144
rect 20176 2208 20492 2209
rect 20176 2144 20182 2208
rect 20246 2144 20262 2208
rect 20326 2144 20342 2208
rect 20406 2144 20422 2208
rect 20486 2144 20492 2208
rect 20176 2143 20492 2144
rect 27604 2208 27920 2209
rect 27604 2144 27610 2208
rect 27674 2144 27690 2208
rect 27754 2144 27770 2208
rect 27834 2144 27850 2208
rect 27914 2144 27920 2208
rect 27604 2143 27920 2144
<< via3 >>
rect 5326 29404 5390 29408
rect 5326 29348 5330 29404
rect 5330 29348 5386 29404
rect 5386 29348 5390 29404
rect 5326 29344 5390 29348
rect 5406 29404 5470 29408
rect 5406 29348 5410 29404
rect 5410 29348 5466 29404
rect 5466 29348 5470 29404
rect 5406 29344 5470 29348
rect 5486 29404 5550 29408
rect 5486 29348 5490 29404
rect 5490 29348 5546 29404
rect 5546 29348 5550 29404
rect 5486 29344 5550 29348
rect 5566 29404 5630 29408
rect 5566 29348 5570 29404
rect 5570 29348 5626 29404
rect 5626 29348 5630 29404
rect 5566 29344 5630 29348
rect 12754 29404 12818 29408
rect 12754 29348 12758 29404
rect 12758 29348 12814 29404
rect 12814 29348 12818 29404
rect 12754 29344 12818 29348
rect 12834 29404 12898 29408
rect 12834 29348 12838 29404
rect 12838 29348 12894 29404
rect 12894 29348 12898 29404
rect 12834 29344 12898 29348
rect 12914 29404 12978 29408
rect 12914 29348 12918 29404
rect 12918 29348 12974 29404
rect 12974 29348 12978 29404
rect 12914 29344 12978 29348
rect 12994 29404 13058 29408
rect 12994 29348 12998 29404
rect 12998 29348 13054 29404
rect 13054 29348 13058 29404
rect 12994 29344 13058 29348
rect 20182 29404 20246 29408
rect 20182 29348 20186 29404
rect 20186 29348 20242 29404
rect 20242 29348 20246 29404
rect 20182 29344 20246 29348
rect 20262 29404 20326 29408
rect 20262 29348 20266 29404
rect 20266 29348 20322 29404
rect 20322 29348 20326 29404
rect 20262 29344 20326 29348
rect 20342 29404 20406 29408
rect 20342 29348 20346 29404
rect 20346 29348 20402 29404
rect 20402 29348 20406 29404
rect 20342 29344 20406 29348
rect 20422 29404 20486 29408
rect 20422 29348 20426 29404
rect 20426 29348 20482 29404
rect 20482 29348 20486 29404
rect 20422 29344 20486 29348
rect 27610 29404 27674 29408
rect 27610 29348 27614 29404
rect 27614 29348 27670 29404
rect 27670 29348 27674 29404
rect 27610 29344 27674 29348
rect 27690 29404 27754 29408
rect 27690 29348 27694 29404
rect 27694 29348 27750 29404
rect 27750 29348 27754 29404
rect 27690 29344 27754 29348
rect 27770 29404 27834 29408
rect 27770 29348 27774 29404
rect 27774 29348 27830 29404
rect 27830 29348 27834 29404
rect 27770 29344 27834 29348
rect 27850 29404 27914 29408
rect 27850 29348 27854 29404
rect 27854 29348 27910 29404
rect 27910 29348 27914 29404
rect 27850 29344 27914 29348
rect 4666 28860 4730 28864
rect 4666 28804 4670 28860
rect 4670 28804 4726 28860
rect 4726 28804 4730 28860
rect 4666 28800 4730 28804
rect 4746 28860 4810 28864
rect 4746 28804 4750 28860
rect 4750 28804 4806 28860
rect 4806 28804 4810 28860
rect 4746 28800 4810 28804
rect 4826 28860 4890 28864
rect 4826 28804 4830 28860
rect 4830 28804 4886 28860
rect 4886 28804 4890 28860
rect 4826 28800 4890 28804
rect 4906 28860 4970 28864
rect 4906 28804 4910 28860
rect 4910 28804 4966 28860
rect 4966 28804 4970 28860
rect 4906 28800 4970 28804
rect 12094 28860 12158 28864
rect 12094 28804 12098 28860
rect 12098 28804 12154 28860
rect 12154 28804 12158 28860
rect 12094 28800 12158 28804
rect 12174 28860 12238 28864
rect 12174 28804 12178 28860
rect 12178 28804 12234 28860
rect 12234 28804 12238 28860
rect 12174 28800 12238 28804
rect 12254 28860 12318 28864
rect 12254 28804 12258 28860
rect 12258 28804 12314 28860
rect 12314 28804 12318 28860
rect 12254 28800 12318 28804
rect 12334 28860 12398 28864
rect 12334 28804 12338 28860
rect 12338 28804 12394 28860
rect 12394 28804 12398 28860
rect 12334 28800 12398 28804
rect 19522 28860 19586 28864
rect 19522 28804 19526 28860
rect 19526 28804 19582 28860
rect 19582 28804 19586 28860
rect 19522 28800 19586 28804
rect 19602 28860 19666 28864
rect 19602 28804 19606 28860
rect 19606 28804 19662 28860
rect 19662 28804 19666 28860
rect 19602 28800 19666 28804
rect 19682 28860 19746 28864
rect 19682 28804 19686 28860
rect 19686 28804 19742 28860
rect 19742 28804 19746 28860
rect 19682 28800 19746 28804
rect 19762 28860 19826 28864
rect 19762 28804 19766 28860
rect 19766 28804 19822 28860
rect 19822 28804 19826 28860
rect 19762 28800 19826 28804
rect 26950 28860 27014 28864
rect 26950 28804 26954 28860
rect 26954 28804 27010 28860
rect 27010 28804 27014 28860
rect 26950 28800 27014 28804
rect 27030 28860 27094 28864
rect 27030 28804 27034 28860
rect 27034 28804 27090 28860
rect 27090 28804 27094 28860
rect 27030 28800 27094 28804
rect 27110 28860 27174 28864
rect 27110 28804 27114 28860
rect 27114 28804 27170 28860
rect 27170 28804 27174 28860
rect 27110 28800 27174 28804
rect 27190 28860 27254 28864
rect 27190 28804 27194 28860
rect 27194 28804 27250 28860
rect 27250 28804 27254 28860
rect 27190 28800 27254 28804
rect 5326 28316 5390 28320
rect 5326 28260 5330 28316
rect 5330 28260 5386 28316
rect 5386 28260 5390 28316
rect 5326 28256 5390 28260
rect 5406 28316 5470 28320
rect 5406 28260 5410 28316
rect 5410 28260 5466 28316
rect 5466 28260 5470 28316
rect 5406 28256 5470 28260
rect 5486 28316 5550 28320
rect 5486 28260 5490 28316
rect 5490 28260 5546 28316
rect 5546 28260 5550 28316
rect 5486 28256 5550 28260
rect 5566 28316 5630 28320
rect 5566 28260 5570 28316
rect 5570 28260 5626 28316
rect 5626 28260 5630 28316
rect 5566 28256 5630 28260
rect 12754 28316 12818 28320
rect 12754 28260 12758 28316
rect 12758 28260 12814 28316
rect 12814 28260 12818 28316
rect 12754 28256 12818 28260
rect 12834 28316 12898 28320
rect 12834 28260 12838 28316
rect 12838 28260 12894 28316
rect 12894 28260 12898 28316
rect 12834 28256 12898 28260
rect 12914 28316 12978 28320
rect 12914 28260 12918 28316
rect 12918 28260 12974 28316
rect 12974 28260 12978 28316
rect 12914 28256 12978 28260
rect 12994 28316 13058 28320
rect 12994 28260 12998 28316
rect 12998 28260 13054 28316
rect 13054 28260 13058 28316
rect 12994 28256 13058 28260
rect 20182 28316 20246 28320
rect 20182 28260 20186 28316
rect 20186 28260 20242 28316
rect 20242 28260 20246 28316
rect 20182 28256 20246 28260
rect 20262 28316 20326 28320
rect 20262 28260 20266 28316
rect 20266 28260 20322 28316
rect 20322 28260 20326 28316
rect 20262 28256 20326 28260
rect 20342 28316 20406 28320
rect 20342 28260 20346 28316
rect 20346 28260 20402 28316
rect 20402 28260 20406 28316
rect 20342 28256 20406 28260
rect 20422 28316 20486 28320
rect 20422 28260 20426 28316
rect 20426 28260 20482 28316
rect 20482 28260 20486 28316
rect 20422 28256 20486 28260
rect 27610 28316 27674 28320
rect 27610 28260 27614 28316
rect 27614 28260 27670 28316
rect 27670 28260 27674 28316
rect 27610 28256 27674 28260
rect 27690 28316 27754 28320
rect 27690 28260 27694 28316
rect 27694 28260 27750 28316
rect 27750 28260 27754 28316
rect 27690 28256 27754 28260
rect 27770 28316 27834 28320
rect 27770 28260 27774 28316
rect 27774 28260 27830 28316
rect 27830 28260 27834 28316
rect 27770 28256 27834 28260
rect 27850 28316 27914 28320
rect 27850 28260 27854 28316
rect 27854 28260 27910 28316
rect 27910 28260 27914 28316
rect 27850 28256 27914 28260
rect 4666 27772 4730 27776
rect 4666 27716 4670 27772
rect 4670 27716 4726 27772
rect 4726 27716 4730 27772
rect 4666 27712 4730 27716
rect 4746 27772 4810 27776
rect 4746 27716 4750 27772
rect 4750 27716 4806 27772
rect 4806 27716 4810 27772
rect 4746 27712 4810 27716
rect 4826 27772 4890 27776
rect 4826 27716 4830 27772
rect 4830 27716 4886 27772
rect 4886 27716 4890 27772
rect 4826 27712 4890 27716
rect 4906 27772 4970 27776
rect 4906 27716 4910 27772
rect 4910 27716 4966 27772
rect 4966 27716 4970 27772
rect 4906 27712 4970 27716
rect 12094 27772 12158 27776
rect 12094 27716 12098 27772
rect 12098 27716 12154 27772
rect 12154 27716 12158 27772
rect 12094 27712 12158 27716
rect 12174 27772 12238 27776
rect 12174 27716 12178 27772
rect 12178 27716 12234 27772
rect 12234 27716 12238 27772
rect 12174 27712 12238 27716
rect 12254 27772 12318 27776
rect 12254 27716 12258 27772
rect 12258 27716 12314 27772
rect 12314 27716 12318 27772
rect 12254 27712 12318 27716
rect 12334 27772 12398 27776
rect 12334 27716 12338 27772
rect 12338 27716 12394 27772
rect 12394 27716 12398 27772
rect 12334 27712 12398 27716
rect 19522 27772 19586 27776
rect 19522 27716 19526 27772
rect 19526 27716 19582 27772
rect 19582 27716 19586 27772
rect 19522 27712 19586 27716
rect 19602 27772 19666 27776
rect 19602 27716 19606 27772
rect 19606 27716 19662 27772
rect 19662 27716 19666 27772
rect 19602 27712 19666 27716
rect 19682 27772 19746 27776
rect 19682 27716 19686 27772
rect 19686 27716 19742 27772
rect 19742 27716 19746 27772
rect 19682 27712 19746 27716
rect 19762 27772 19826 27776
rect 19762 27716 19766 27772
rect 19766 27716 19822 27772
rect 19822 27716 19826 27772
rect 19762 27712 19826 27716
rect 26950 27772 27014 27776
rect 26950 27716 26954 27772
rect 26954 27716 27010 27772
rect 27010 27716 27014 27772
rect 26950 27712 27014 27716
rect 27030 27772 27094 27776
rect 27030 27716 27034 27772
rect 27034 27716 27090 27772
rect 27090 27716 27094 27772
rect 27030 27712 27094 27716
rect 27110 27772 27174 27776
rect 27110 27716 27114 27772
rect 27114 27716 27170 27772
rect 27170 27716 27174 27772
rect 27110 27712 27174 27716
rect 27190 27772 27254 27776
rect 27190 27716 27194 27772
rect 27194 27716 27250 27772
rect 27250 27716 27254 27772
rect 27190 27712 27254 27716
rect 5326 27228 5390 27232
rect 5326 27172 5330 27228
rect 5330 27172 5386 27228
rect 5386 27172 5390 27228
rect 5326 27168 5390 27172
rect 5406 27228 5470 27232
rect 5406 27172 5410 27228
rect 5410 27172 5466 27228
rect 5466 27172 5470 27228
rect 5406 27168 5470 27172
rect 5486 27228 5550 27232
rect 5486 27172 5490 27228
rect 5490 27172 5546 27228
rect 5546 27172 5550 27228
rect 5486 27168 5550 27172
rect 5566 27228 5630 27232
rect 5566 27172 5570 27228
rect 5570 27172 5626 27228
rect 5626 27172 5630 27228
rect 5566 27168 5630 27172
rect 12754 27228 12818 27232
rect 12754 27172 12758 27228
rect 12758 27172 12814 27228
rect 12814 27172 12818 27228
rect 12754 27168 12818 27172
rect 12834 27228 12898 27232
rect 12834 27172 12838 27228
rect 12838 27172 12894 27228
rect 12894 27172 12898 27228
rect 12834 27168 12898 27172
rect 12914 27228 12978 27232
rect 12914 27172 12918 27228
rect 12918 27172 12974 27228
rect 12974 27172 12978 27228
rect 12914 27168 12978 27172
rect 12994 27228 13058 27232
rect 12994 27172 12998 27228
rect 12998 27172 13054 27228
rect 13054 27172 13058 27228
rect 12994 27168 13058 27172
rect 20182 27228 20246 27232
rect 20182 27172 20186 27228
rect 20186 27172 20242 27228
rect 20242 27172 20246 27228
rect 20182 27168 20246 27172
rect 20262 27228 20326 27232
rect 20262 27172 20266 27228
rect 20266 27172 20322 27228
rect 20322 27172 20326 27228
rect 20262 27168 20326 27172
rect 20342 27228 20406 27232
rect 20342 27172 20346 27228
rect 20346 27172 20402 27228
rect 20402 27172 20406 27228
rect 20342 27168 20406 27172
rect 20422 27228 20486 27232
rect 20422 27172 20426 27228
rect 20426 27172 20482 27228
rect 20482 27172 20486 27228
rect 20422 27168 20486 27172
rect 27610 27228 27674 27232
rect 27610 27172 27614 27228
rect 27614 27172 27670 27228
rect 27670 27172 27674 27228
rect 27610 27168 27674 27172
rect 27690 27228 27754 27232
rect 27690 27172 27694 27228
rect 27694 27172 27750 27228
rect 27750 27172 27754 27228
rect 27690 27168 27754 27172
rect 27770 27228 27834 27232
rect 27770 27172 27774 27228
rect 27774 27172 27830 27228
rect 27830 27172 27834 27228
rect 27770 27168 27834 27172
rect 27850 27228 27914 27232
rect 27850 27172 27854 27228
rect 27854 27172 27910 27228
rect 27910 27172 27914 27228
rect 27850 27168 27914 27172
rect 4666 26684 4730 26688
rect 4666 26628 4670 26684
rect 4670 26628 4726 26684
rect 4726 26628 4730 26684
rect 4666 26624 4730 26628
rect 4746 26684 4810 26688
rect 4746 26628 4750 26684
rect 4750 26628 4806 26684
rect 4806 26628 4810 26684
rect 4746 26624 4810 26628
rect 4826 26684 4890 26688
rect 4826 26628 4830 26684
rect 4830 26628 4886 26684
rect 4886 26628 4890 26684
rect 4826 26624 4890 26628
rect 4906 26684 4970 26688
rect 4906 26628 4910 26684
rect 4910 26628 4966 26684
rect 4966 26628 4970 26684
rect 4906 26624 4970 26628
rect 12094 26684 12158 26688
rect 12094 26628 12098 26684
rect 12098 26628 12154 26684
rect 12154 26628 12158 26684
rect 12094 26624 12158 26628
rect 12174 26684 12238 26688
rect 12174 26628 12178 26684
rect 12178 26628 12234 26684
rect 12234 26628 12238 26684
rect 12174 26624 12238 26628
rect 12254 26684 12318 26688
rect 12254 26628 12258 26684
rect 12258 26628 12314 26684
rect 12314 26628 12318 26684
rect 12254 26624 12318 26628
rect 12334 26684 12398 26688
rect 12334 26628 12338 26684
rect 12338 26628 12394 26684
rect 12394 26628 12398 26684
rect 12334 26624 12398 26628
rect 19522 26684 19586 26688
rect 19522 26628 19526 26684
rect 19526 26628 19582 26684
rect 19582 26628 19586 26684
rect 19522 26624 19586 26628
rect 19602 26684 19666 26688
rect 19602 26628 19606 26684
rect 19606 26628 19662 26684
rect 19662 26628 19666 26684
rect 19602 26624 19666 26628
rect 19682 26684 19746 26688
rect 19682 26628 19686 26684
rect 19686 26628 19742 26684
rect 19742 26628 19746 26684
rect 19682 26624 19746 26628
rect 19762 26684 19826 26688
rect 19762 26628 19766 26684
rect 19766 26628 19822 26684
rect 19822 26628 19826 26684
rect 19762 26624 19826 26628
rect 26950 26684 27014 26688
rect 26950 26628 26954 26684
rect 26954 26628 27010 26684
rect 27010 26628 27014 26684
rect 26950 26624 27014 26628
rect 27030 26684 27094 26688
rect 27030 26628 27034 26684
rect 27034 26628 27090 26684
rect 27090 26628 27094 26684
rect 27030 26624 27094 26628
rect 27110 26684 27174 26688
rect 27110 26628 27114 26684
rect 27114 26628 27170 26684
rect 27170 26628 27174 26684
rect 27110 26624 27174 26628
rect 27190 26684 27254 26688
rect 27190 26628 27194 26684
rect 27194 26628 27250 26684
rect 27250 26628 27254 26684
rect 27190 26624 27254 26628
rect 5326 26140 5390 26144
rect 5326 26084 5330 26140
rect 5330 26084 5386 26140
rect 5386 26084 5390 26140
rect 5326 26080 5390 26084
rect 5406 26140 5470 26144
rect 5406 26084 5410 26140
rect 5410 26084 5466 26140
rect 5466 26084 5470 26140
rect 5406 26080 5470 26084
rect 5486 26140 5550 26144
rect 5486 26084 5490 26140
rect 5490 26084 5546 26140
rect 5546 26084 5550 26140
rect 5486 26080 5550 26084
rect 5566 26140 5630 26144
rect 5566 26084 5570 26140
rect 5570 26084 5626 26140
rect 5626 26084 5630 26140
rect 5566 26080 5630 26084
rect 12754 26140 12818 26144
rect 12754 26084 12758 26140
rect 12758 26084 12814 26140
rect 12814 26084 12818 26140
rect 12754 26080 12818 26084
rect 12834 26140 12898 26144
rect 12834 26084 12838 26140
rect 12838 26084 12894 26140
rect 12894 26084 12898 26140
rect 12834 26080 12898 26084
rect 12914 26140 12978 26144
rect 12914 26084 12918 26140
rect 12918 26084 12974 26140
rect 12974 26084 12978 26140
rect 12914 26080 12978 26084
rect 12994 26140 13058 26144
rect 12994 26084 12998 26140
rect 12998 26084 13054 26140
rect 13054 26084 13058 26140
rect 12994 26080 13058 26084
rect 20182 26140 20246 26144
rect 20182 26084 20186 26140
rect 20186 26084 20242 26140
rect 20242 26084 20246 26140
rect 20182 26080 20246 26084
rect 20262 26140 20326 26144
rect 20262 26084 20266 26140
rect 20266 26084 20322 26140
rect 20322 26084 20326 26140
rect 20262 26080 20326 26084
rect 20342 26140 20406 26144
rect 20342 26084 20346 26140
rect 20346 26084 20402 26140
rect 20402 26084 20406 26140
rect 20342 26080 20406 26084
rect 20422 26140 20486 26144
rect 20422 26084 20426 26140
rect 20426 26084 20482 26140
rect 20482 26084 20486 26140
rect 20422 26080 20486 26084
rect 27610 26140 27674 26144
rect 27610 26084 27614 26140
rect 27614 26084 27670 26140
rect 27670 26084 27674 26140
rect 27610 26080 27674 26084
rect 27690 26140 27754 26144
rect 27690 26084 27694 26140
rect 27694 26084 27750 26140
rect 27750 26084 27754 26140
rect 27690 26080 27754 26084
rect 27770 26140 27834 26144
rect 27770 26084 27774 26140
rect 27774 26084 27830 26140
rect 27830 26084 27834 26140
rect 27770 26080 27834 26084
rect 27850 26140 27914 26144
rect 27850 26084 27854 26140
rect 27854 26084 27910 26140
rect 27910 26084 27914 26140
rect 27850 26080 27914 26084
rect 4666 25596 4730 25600
rect 4666 25540 4670 25596
rect 4670 25540 4726 25596
rect 4726 25540 4730 25596
rect 4666 25536 4730 25540
rect 4746 25596 4810 25600
rect 4746 25540 4750 25596
rect 4750 25540 4806 25596
rect 4806 25540 4810 25596
rect 4746 25536 4810 25540
rect 4826 25596 4890 25600
rect 4826 25540 4830 25596
rect 4830 25540 4886 25596
rect 4886 25540 4890 25596
rect 4826 25536 4890 25540
rect 4906 25596 4970 25600
rect 4906 25540 4910 25596
rect 4910 25540 4966 25596
rect 4966 25540 4970 25596
rect 4906 25536 4970 25540
rect 12094 25596 12158 25600
rect 12094 25540 12098 25596
rect 12098 25540 12154 25596
rect 12154 25540 12158 25596
rect 12094 25536 12158 25540
rect 12174 25596 12238 25600
rect 12174 25540 12178 25596
rect 12178 25540 12234 25596
rect 12234 25540 12238 25596
rect 12174 25536 12238 25540
rect 12254 25596 12318 25600
rect 12254 25540 12258 25596
rect 12258 25540 12314 25596
rect 12314 25540 12318 25596
rect 12254 25536 12318 25540
rect 12334 25596 12398 25600
rect 12334 25540 12338 25596
rect 12338 25540 12394 25596
rect 12394 25540 12398 25596
rect 12334 25536 12398 25540
rect 19522 25596 19586 25600
rect 19522 25540 19526 25596
rect 19526 25540 19582 25596
rect 19582 25540 19586 25596
rect 19522 25536 19586 25540
rect 19602 25596 19666 25600
rect 19602 25540 19606 25596
rect 19606 25540 19662 25596
rect 19662 25540 19666 25596
rect 19602 25536 19666 25540
rect 19682 25596 19746 25600
rect 19682 25540 19686 25596
rect 19686 25540 19742 25596
rect 19742 25540 19746 25596
rect 19682 25536 19746 25540
rect 19762 25596 19826 25600
rect 19762 25540 19766 25596
rect 19766 25540 19822 25596
rect 19822 25540 19826 25596
rect 19762 25536 19826 25540
rect 26950 25596 27014 25600
rect 26950 25540 26954 25596
rect 26954 25540 27010 25596
rect 27010 25540 27014 25596
rect 26950 25536 27014 25540
rect 27030 25596 27094 25600
rect 27030 25540 27034 25596
rect 27034 25540 27090 25596
rect 27090 25540 27094 25596
rect 27030 25536 27094 25540
rect 27110 25596 27174 25600
rect 27110 25540 27114 25596
rect 27114 25540 27170 25596
rect 27170 25540 27174 25596
rect 27110 25536 27174 25540
rect 27190 25596 27254 25600
rect 27190 25540 27194 25596
rect 27194 25540 27250 25596
rect 27250 25540 27254 25596
rect 27190 25536 27254 25540
rect 5326 25052 5390 25056
rect 5326 24996 5330 25052
rect 5330 24996 5386 25052
rect 5386 24996 5390 25052
rect 5326 24992 5390 24996
rect 5406 25052 5470 25056
rect 5406 24996 5410 25052
rect 5410 24996 5466 25052
rect 5466 24996 5470 25052
rect 5406 24992 5470 24996
rect 5486 25052 5550 25056
rect 5486 24996 5490 25052
rect 5490 24996 5546 25052
rect 5546 24996 5550 25052
rect 5486 24992 5550 24996
rect 5566 25052 5630 25056
rect 5566 24996 5570 25052
rect 5570 24996 5626 25052
rect 5626 24996 5630 25052
rect 5566 24992 5630 24996
rect 12754 25052 12818 25056
rect 12754 24996 12758 25052
rect 12758 24996 12814 25052
rect 12814 24996 12818 25052
rect 12754 24992 12818 24996
rect 12834 25052 12898 25056
rect 12834 24996 12838 25052
rect 12838 24996 12894 25052
rect 12894 24996 12898 25052
rect 12834 24992 12898 24996
rect 12914 25052 12978 25056
rect 12914 24996 12918 25052
rect 12918 24996 12974 25052
rect 12974 24996 12978 25052
rect 12914 24992 12978 24996
rect 12994 25052 13058 25056
rect 12994 24996 12998 25052
rect 12998 24996 13054 25052
rect 13054 24996 13058 25052
rect 12994 24992 13058 24996
rect 20182 25052 20246 25056
rect 20182 24996 20186 25052
rect 20186 24996 20242 25052
rect 20242 24996 20246 25052
rect 20182 24992 20246 24996
rect 20262 25052 20326 25056
rect 20262 24996 20266 25052
rect 20266 24996 20322 25052
rect 20322 24996 20326 25052
rect 20262 24992 20326 24996
rect 20342 25052 20406 25056
rect 20342 24996 20346 25052
rect 20346 24996 20402 25052
rect 20402 24996 20406 25052
rect 20342 24992 20406 24996
rect 20422 25052 20486 25056
rect 20422 24996 20426 25052
rect 20426 24996 20482 25052
rect 20482 24996 20486 25052
rect 20422 24992 20486 24996
rect 27610 25052 27674 25056
rect 27610 24996 27614 25052
rect 27614 24996 27670 25052
rect 27670 24996 27674 25052
rect 27610 24992 27674 24996
rect 27690 25052 27754 25056
rect 27690 24996 27694 25052
rect 27694 24996 27750 25052
rect 27750 24996 27754 25052
rect 27690 24992 27754 24996
rect 27770 25052 27834 25056
rect 27770 24996 27774 25052
rect 27774 24996 27830 25052
rect 27830 24996 27834 25052
rect 27770 24992 27834 24996
rect 27850 25052 27914 25056
rect 27850 24996 27854 25052
rect 27854 24996 27910 25052
rect 27910 24996 27914 25052
rect 27850 24992 27914 24996
rect 4666 24508 4730 24512
rect 4666 24452 4670 24508
rect 4670 24452 4726 24508
rect 4726 24452 4730 24508
rect 4666 24448 4730 24452
rect 4746 24508 4810 24512
rect 4746 24452 4750 24508
rect 4750 24452 4806 24508
rect 4806 24452 4810 24508
rect 4746 24448 4810 24452
rect 4826 24508 4890 24512
rect 4826 24452 4830 24508
rect 4830 24452 4886 24508
rect 4886 24452 4890 24508
rect 4826 24448 4890 24452
rect 4906 24508 4970 24512
rect 4906 24452 4910 24508
rect 4910 24452 4966 24508
rect 4966 24452 4970 24508
rect 4906 24448 4970 24452
rect 12094 24508 12158 24512
rect 12094 24452 12098 24508
rect 12098 24452 12154 24508
rect 12154 24452 12158 24508
rect 12094 24448 12158 24452
rect 12174 24508 12238 24512
rect 12174 24452 12178 24508
rect 12178 24452 12234 24508
rect 12234 24452 12238 24508
rect 12174 24448 12238 24452
rect 12254 24508 12318 24512
rect 12254 24452 12258 24508
rect 12258 24452 12314 24508
rect 12314 24452 12318 24508
rect 12254 24448 12318 24452
rect 12334 24508 12398 24512
rect 12334 24452 12338 24508
rect 12338 24452 12394 24508
rect 12394 24452 12398 24508
rect 12334 24448 12398 24452
rect 19522 24508 19586 24512
rect 19522 24452 19526 24508
rect 19526 24452 19582 24508
rect 19582 24452 19586 24508
rect 19522 24448 19586 24452
rect 19602 24508 19666 24512
rect 19602 24452 19606 24508
rect 19606 24452 19662 24508
rect 19662 24452 19666 24508
rect 19602 24448 19666 24452
rect 19682 24508 19746 24512
rect 19682 24452 19686 24508
rect 19686 24452 19742 24508
rect 19742 24452 19746 24508
rect 19682 24448 19746 24452
rect 19762 24508 19826 24512
rect 19762 24452 19766 24508
rect 19766 24452 19822 24508
rect 19822 24452 19826 24508
rect 19762 24448 19826 24452
rect 26950 24508 27014 24512
rect 26950 24452 26954 24508
rect 26954 24452 27010 24508
rect 27010 24452 27014 24508
rect 26950 24448 27014 24452
rect 27030 24508 27094 24512
rect 27030 24452 27034 24508
rect 27034 24452 27090 24508
rect 27090 24452 27094 24508
rect 27030 24448 27094 24452
rect 27110 24508 27174 24512
rect 27110 24452 27114 24508
rect 27114 24452 27170 24508
rect 27170 24452 27174 24508
rect 27110 24448 27174 24452
rect 27190 24508 27254 24512
rect 27190 24452 27194 24508
rect 27194 24452 27250 24508
rect 27250 24452 27254 24508
rect 27190 24448 27254 24452
rect 5326 23964 5390 23968
rect 5326 23908 5330 23964
rect 5330 23908 5386 23964
rect 5386 23908 5390 23964
rect 5326 23904 5390 23908
rect 5406 23964 5470 23968
rect 5406 23908 5410 23964
rect 5410 23908 5466 23964
rect 5466 23908 5470 23964
rect 5406 23904 5470 23908
rect 5486 23964 5550 23968
rect 5486 23908 5490 23964
rect 5490 23908 5546 23964
rect 5546 23908 5550 23964
rect 5486 23904 5550 23908
rect 5566 23964 5630 23968
rect 5566 23908 5570 23964
rect 5570 23908 5626 23964
rect 5626 23908 5630 23964
rect 5566 23904 5630 23908
rect 12754 23964 12818 23968
rect 12754 23908 12758 23964
rect 12758 23908 12814 23964
rect 12814 23908 12818 23964
rect 12754 23904 12818 23908
rect 12834 23964 12898 23968
rect 12834 23908 12838 23964
rect 12838 23908 12894 23964
rect 12894 23908 12898 23964
rect 12834 23904 12898 23908
rect 12914 23964 12978 23968
rect 12914 23908 12918 23964
rect 12918 23908 12974 23964
rect 12974 23908 12978 23964
rect 12914 23904 12978 23908
rect 12994 23964 13058 23968
rect 12994 23908 12998 23964
rect 12998 23908 13054 23964
rect 13054 23908 13058 23964
rect 12994 23904 13058 23908
rect 20182 23964 20246 23968
rect 20182 23908 20186 23964
rect 20186 23908 20242 23964
rect 20242 23908 20246 23964
rect 20182 23904 20246 23908
rect 20262 23964 20326 23968
rect 20262 23908 20266 23964
rect 20266 23908 20322 23964
rect 20322 23908 20326 23964
rect 20262 23904 20326 23908
rect 20342 23964 20406 23968
rect 20342 23908 20346 23964
rect 20346 23908 20402 23964
rect 20402 23908 20406 23964
rect 20342 23904 20406 23908
rect 20422 23964 20486 23968
rect 20422 23908 20426 23964
rect 20426 23908 20482 23964
rect 20482 23908 20486 23964
rect 20422 23904 20486 23908
rect 27610 23964 27674 23968
rect 27610 23908 27614 23964
rect 27614 23908 27670 23964
rect 27670 23908 27674 23964
rect 27610 23904 27674 23908
rect 27690 23964 27754 23968
rect 27690 23908 27694 23964
rect 27694 23908 27750 23964
rect 27750 23908 27754 23964
rect 27690 23904 27754 23908
rect 27770 23964 27834 23968
rect 27770 23908 27774 23964
rect 27774 23908 27830 23964
rect 27830 23908 27834 23964
rect 27770 23904 27834 23908
rect 27850 23964 27914 23968
rect 27850 23908 27854 23964
rect 27854 23908 27910 23964
rect 27910 23908 27914 23964
rect 27850 23904 27914 23908
rect 4666 23420 4730 23424
rect 4666 23364 4670 23420
rect 4670 23364 4726 23420
rect 4726 23364 4730 23420
rect 4666 23360 4730 23364
rect 4746 23420 4810 23424
rect 4746 23364 4750 23420
rect 4750 23364 4806 23420
rect 4806 23364 4810 23420
rect 4746 23360 4810 23364
rect 4826 23420 4890 23424
rect 4826 23364 4830 23420
rect 4830 23364 4886 23420
rect 4886 23364 4890 23420
rect 4826 23360 4890 23364
rect 4906 23420 4970 23424
rect 4906 23364 4910 23420
rect 4910 23364 4966 23420
rect 4966 23364 4970 23420
rect 4906 23360 4970 23364
rect 12094 23420 12158 23424
rect 12094 23364 12098 23420
rect 12098 23364 12154 23420
rect 12154 23364 12158 23420
rect 12094 23360 12158 23364
rect 12174 23420 12238 23424
rect 12174 23364 12178 23420
rect 12178 23364 12234 23420
rect 12234 23364 12238 23420
rect 12174 23360 12238 23364
rect 12254 23420 12318 23424
rect 12254 23364 12258 23420
rect 12258 23364 12314 23420
rect 12314 23364 12318 23420
rect 12254 23360 12318 23364
rect 12334 23420 12398 23424
rect 12334 23364 12338 23420
rect 12338 23364 12394 23420
rect 12394 23364 12398 23420
rect 12334 23360 12398 23364
rect 19522 23420 19586 23424
rect 19522 23364 19526 23420
rect 19526 23364 19582 23420
rect 19582 23364 19586 23420
rect 19522 23360 19586 23364
rect 19602 23420 19666 23424
rect 19602 23364 19606 23420
rect 19606 23364 19662 23420
rect 19662 23364 19666 23420
rect 19602 23360 19666 23364
rect 19682 23420 19746 23424
rect 19682 23364 19686 23420
rect 19686 23364 19742 23420
rect 19742 23364 19746 23420
rect 19682 23360 19746 23364
rect 19762 23420 19826 23424
rect 19762 23364 19766 23420
rect 19766 23364 19822 23420
rect 19822 23364 19826 23420
rect 19762 23360 19826 23364
rect 26950 23420 27014 23424
rect 26950 23364 26954 23420
rect 26954 23364 27010 23420
rect 27010 23364 27014 23420
rect 26950 23360 27014 23364
rect 27030 23420 27094 23424
rect 27030 23364 27034 23420
rect 27034 23364 27090 23420
rect 27090 23364 27094 23420
rect 27030 23360 27094 23364
rect 27110 23420 27174 23424
rect 27110 23364 27114 23420
rect 27114 23364 27170 23420
rect 27170 23364 27174 23420
rect 27110 23360 27174 23364
rect 27190 23420 27254 23424
rect 27190 23364 27194 23420
rect 27194 23364 27250 23420
rect 27250 23364 27254 23420
rect 27190 23360 27254 23364
rect 5326 22876 5390 22880
rect 5326 22820 5330 22876
rect 5330 22820 5386 22876
rect 5386 22820 5390 22876
rect 5326 22816 5390 22820
rect 5406 22876 5470 22880
rect 5406 22820 5410 22876
rect 5410 22820 5466 22876
rect 5466 22820 5470 22876
rect 5406 22816 5470 22820
rect 5486 22876 5550 22880
rect 5486 22820 5490 22876
rect 5490 22820 5546 22876
rect 5546 22820 5550 22876
rect 5486 22816 5550 22820
rect 5566 22876 5630 22880
rect 5566 22820 5570 22876
rect 5570 22820 5626 22876
rect 5626 22820 5630 22876
rect 5566 22816 5630 22820
rect 12754 22876 12818 22880
rect 12754 22820 12758 22876
rect 12758 22820 12814 22876
rect 12814 22820 12818 22876
rect 12754 22816 12818 22820
rect 12834 22876 12898 22880
rect 12834 22820 12838 22876
rect 12838 22820 12894 22876
rect 12894 22820 12898 22876
rect 12834 22816 12898 22820
rect 12914 22876 12978 22880
rect 12914 22820 12918 22876
rect 12918 22820 12974 22876
rect 12974 22820 12978 22876
rect 12914 22816 12978 22820
rect 12994 22876 13058 22880
rect 12994 22820 12998 22876
rect 12998 22820 13054 22876
rect 13054 22820 13058 22876
rect 12994 22816 13058 22820
rect 20182 22876 20246 22880
rect 20182 22820 20186 22876
rect 20186 22820 20242 22876
rect 20242 22820 20246 22876
rect 20182 22816 20246 22820
rect 20262 22876 20326 22880
rect 20262 22820 20266 22876
rect 20266 22820 20322 22876
rect 20322 22820 20326 22876
rect 20262 22816 20326 22820
rect 20342 22876 20406 22880
rect 20342 22820 20346 22876
rect 20346 22820 20402 22876
rect 20402 22820 20406 22876
rect 20342 22816 20406 22820
rect 20422 22876 20486 22880
rect 20422 22820 20426 22876
rect 20426 22820 20482 22876
rect 20482 22820 20486 22876
rect 20422 22816 20486 22820
rect 27610 22876 27674 22880
rect 27610 22820 27614 22876
rect 27614 22820 27670 22876
rect 27670 22820 27674 22876
rect 27610 22816 27674 22820
rect 27690 22876 27754 22880
rect 27690 22820 27694 22876
rect 27694 22820 27750 22876
rect 27750 22820 27754 22876
rect 27690 22816 27754 22820
rect 27770 22876 27834 22880
rect 27770 22820 27774 22876
rect 27774 22820 27830 22876
rect 27830 22820 27834 22876
rect 27770 22816 27834 22820
rect 27850 22876 27914 22880
rect 27850 22820 27854 22876
rect 27854 22820 27910 22876
rect 27910 22820 27914 22876
rect 27850 22816 27914 22820
rect 4666 22332 4730 22336
rect 4666 22276 4670 22332
rect 4670 22276 4726 22332
rect 4726 22276 4730 22332
rect 4666 22272 4730 22276
rect 4746 22332 4810 22336
rect 4746 22276 4750 22332
rect 4750 22276 4806 22332
rect 4806 22276 4810 22332
rect 4746 22272 4810 22276
rect 4826 22332 4890 22336
rect 4826 22276 4830 22332
rect 4830 22276 4886 22332
rect 4886 22276 4890 22332
rect 4826 22272 4890 22276
rect 4906 22332 4970 22336
rect 4906 22276 4910 22332
rect 4910 22276 4966 22332
rect 4966 22276 4970 22332
rect 4906 22272 4970 22276
rect 12094 22332 12158 22336
rect 12094 22276 12098 22332
rect 12098 22276 12154 22332
rect 12154 22276 12158 22332
rect 12094 22272 12158 22276
rect 12174 22332 12238 22336
rect 12174 22276 12178 22332
rect 12178 22276 12234 22332
rect 12234 22276 12238 22332
rect 12174 22272 12238 22276
rect 12254 22332 12318 22336
rect 12254 22276 12258 22332
rect 12258 22276 12314 22332
rect 12314 22276 12318 22332
rect 12254 22272 12318 22276
rect 12334 22332 12398 22336
rect 12334 22276 12338 22332
rect 12338 22276 12394 22332
rect 12394 22276 12398 22332
rect 12334 22272 12398 22276
rect 19522 22332 19586 22336
rect 19522 22276 19526 22332
rect 19526 22276 19582 22332
rect 19582 22276 19586 22332
rect 19522 22272 19586 22276
rect 19602 22332 19666 22336
rect 19602 22276 19606 22332
rect 19606 22276 19662 22332
rect 19662 22276 19666 22332
rect 19602 22272 19666 22276
rect 19682 22332 19746 22336
rect 19682 22276 19686 22332
rect 19686 22276 19742 22332
rect 19742 22276 19746 22332
rect 19682 22272 19746 22276
rect 19762 22332 19826 22336
rect 19762 22276 19766 22332
rect 19766 22276 19822 22332
rect 19822 22276 19826 22332
rect 19762 22272 19826 22276
rect 26950 22332 27014 22336
rect 26950 22276 26954 22332
rect 26954 22276 27010 22332
rect 27010 22276 27014 22332
rect 26950 22272 27014 22276
rect 27030 22332 27094 22336
rect 27030 22276 27034 22332
rect 27034 22276 27090 22332
rect 27090 22276 27094 22332
rect 27030 22272 27094 22276
rect 27110 22332 27174 22336
rect 27110 22276 27114 22332
rect 27114 22276 27170 22332
rect 27170 22276 27174 22332
rect 27110 22272 27174 22276
rect 27190 22332 27254 22336
rect 27190 22276 27194 22332
rect 27194 22276 27250 22332
rect 27250 22276 27254 22332
rect 27190 22272 27254 22276
rect 5326 21788 5390 21792
rect 5326 21732 5330 21788
rect 5330 21732 5386 21788
rect 5386 21732 5390 21788
rect 5326 21728 5390 21732
rect 5406 21788 5470 21792
rect 5406 21732 5410 21788
rect 5410 21732 5466 21788
rect 5466 21732 5470 21788
rect 5406 21728 5470 21732
rect 5486 21788 5550 21792
rect 5486 21732 5490 21788
rect 5490 21732 5546 21788
rect 5546 21732 5550 21788
rect 5486 21728 5550 21732
rect 5566 21788 5630 21792
rect 5566 21732 5570 21788
rect 5570 21732 5626 21788
rect 5626 21732 5630 21788
rect 5566 21728 5630 21732
rect 12754 21788 12818 21792
rect 12754 21732 12758 21788
rect 12758 21732 12814 21788
rect 12814 21732 12818 21788
rect 12754 21728 12818 21732
rect 12834 21788 12898 21792
rect 12834 21732 12838 21788
rect 12838 21732 12894 21788
rect 12894 21732 12898 21788
rect 12834 21728 12898 21732
rect 12914 21788 12978 21792
rect 12914 21732 12918 21788
rect 12918 21732 12974 21788
rect 12974 21732 12978 21788
rect 12914 21728 12978 21732
rect 12994 21788 13058 21792
rect 12994 21732 12998 21788
rect 12998 21732 13054 21788
rect 13054 21732 13058 21788
rect 12994 21728 13058 21732
rect 20182 21788 20246 21792
rect 20182 21732 20186 21788
rect 20186 21732 20242 21788
rect 20242 21732 20246 21788
rect 20182 21728 20246 21732
rect 20262 21788 20326 21792
rect 20262 21732 20266 21788
rect 20266 21732 20322 21788
rect 20322 21732 20326 21788
rect 20262 21728 20326 21732
rect 20342 21788 20406 21792
rect 20342 21732 20346 21788
rect 20346 21732 20402 21788
rect 20402 21732 20406 21788
rect 20342 21728 20406 21732
rect 20422 21788 20486 21792
rect 20422 21732 20426 21788
rect 20426 21732 20482 21788
rect 20482 21732 20486 21788
rect 20422 21728 20486 21732
rect 27610 21788 27674 21792
rect 27610 21732 27614 21788
rect 27614 21732 27670 21788
rect 27670 21732 27674 21788
rect 27610 21728 27674 21732
rect 27690 21788 27754 21792
rect 27690 21732 27694 21788
rect 27694 21732 27750 21788
rect 27750 21732 27754 21788
rect 27690 21728 27754 21732
rect 27770 21788 27834 21792
rect 27770 21732 27774 21788
rect 27774 21732 27830 21788
rect 27830 21732 27834 21788
rect 27770 21728 27834 21732
rect 27850 21788 27914 21792
rect 27850 21732 27854 21788
rect 27854 21732 27910 21788
rect 27910 21732 27914 21788
rect 27850 21728 27914 21732
rect 4666 21244 4730 21248
rect 4666 21188 4670 21244
rect 4670 21188 4726 21244
rect 4726 21188 4730 21244
rect 4666 21184 4730 21188
rect 4746 21244 4810 21248
rect 4746 21188 4750 21244
rect 4750 21188 4806 21244
rect 4806 21188 4810 21244
rect 4746 21184 4810 21188
rect 4826 21244 4890 21248
rect 4826 21188 4830 21244
rect 4830 21188 4886 21244
rect 4886 21188 4890 21244
rect 4826 21184 4890 21188
rect 4906 21244 4970 21248
rect 4906 21188 4910 21244
rect 4910 21188 4966 21244
rect 4966 21188 4970 21244
rect 4906 21184 4970 21188
rect 12094 21244 12158 21248
rect 12094 21188 12098 21244
rect 12098 21188 12154 21244
rect 12154 21188 12158 21244
rect 12094 21184 12158 21188
rect 12174 21244 12238 21248
rect 12174 21188 12178 21244
rect 12178 21188 12234 21244
rect 12234 21188 12238 21244
rect 12174 21184 12238 21188
rect 12254 21244 12318 21248
rect 12254 21188 12258 21244
rect 12258 21188 12314 21244
rect 12314 21188 12318 21244
rect 12254 21184 12318 21188
rect 12334 21244 12398 21248
rect 12334 21188 12338 21244
rect 12338 21188 12394 21244
rect 12394 21188 12398 21244
rect 12334 21184 12398 21188
rect 19522 21244 19586 21248
rect 19522 21188 19526 21244
rect 19526 21188 19582 21244
rect 19582 21188 19586 21244
rect 19522 21184 19586 21188
rect 19602 21244 19666 21248
rect 19602 21188 19606 21244
rect 19606 21188 19662 21244
rect 19662 21188 19666 21244
rect 19602 21184 19666 21188
rect 19682 21244 19746 21248
rect 19682 21188 19686 21244
rect 19686 21188 19742 21244
rect 19742 21188 19746 21244
rect 19682 21184 19746 21188
rect 19762 21244 19826 21248
rect 19762 21188 19766 21244
rect 19766 21188 19822 21244
rect 19822 21188 19826 21244
rect 19762 21184 19826 21188
rect 26950 21244 27014 21248
rect 26950 21188 26954 21244
rect 26954 21188 27010 21244
rect 27010 21188 27014 21244
rect 26950 21184 27014 21188
rect 27030 21244 27094 21248
rect 27030 21188 27034 21244
rect 27034 21188 27090 21244
rect 27090 21188 27094 21244
rect 27030 21184 27094 21188
rect 27110 21244 27174 21248
rect 27110 21188 27114 21244
rect 27114 21188 27170 21244
rect 27170 21188 27174 21244
rect 27110 21184 27174 21188
rect 27190 21244 27254 21248
rect 27190 21188 27194 21244
rect 27194 21188 27250 21244
rect 27250 21188 27254 21244
rect 27190 21184 27254 21188
rect 5326 20700 5390 20704
rect 5326 20644 5330 20700
rect 5330 20644 5386 20700
rect 5386 20644 5390 20700
rect 5326 20640 5390 20644
rect 5406 20700 5470 20704
rect 5406 20644 5410 20700
rect 5410 20644 5466 20700
rect 5466 20644 5470 20700
rect 5406 20640 5470 20644
rect 5486 20700 5550 20704
rect 5486 20644 5490 20700
rect 5490 20644 5546 20700
rect 5546 20644 5550 20700
rect 5486 20640 5550 20644
rect 5566 20700 5630 20704
rect 5566 20644 5570 20700
rect 5570 20644 5626 20700
rect 5626 20644 5630 20700
rect 5566 20640 5630 20644
rect 12754 20700 12818 20704
rect 12754 20644 12758 20700
rect 12758 20644 12814 20700
rect 12814 20644 12818 20700
rect 12754 20640 12818 20644
rect 12834 20700 12898 20704
rect 12834 20644 12838 20700
rect 12838 20644 12894 20700
rect 12894 20644 12898 20700
rect 12834 20640 12898 20644
rect 12914 20700 12978 20704
rect 12914 20644 12918 20700
rect 12918 20644 12974 20700
rect 12974 20644 12978 20700
rect 12914 20640 12978 20644
rect 12994 20700 13058 20704
rect 12994 20644 12998 20700
rect 12998 20644 13054 20700
rect 13054 20644 13058 20700
rect 12994 20640 13058 20644
rect 20182 20700 20246 20704
rect 20182 20644 20186 20700
rect 20186 20644 20242 20700
rect 20242 20644 20246 20700
rect 20182 20640 20246 20644
rect 20262 20700 20326 20704
rect 20262 20644 20266 20700
rect 20266 20644 20322 20700
rect 20322 20644 20326 20700
rect 20262 20640 20326 20644
rect 20342 20700 20406 20704
rect 20342 20644 20346 20700
rect 20346 20644 20402 20700
rect 20402 20644 20406 20700
rect 20342 20640 20406 20644
rect 20422 20700 20486 20704
rect 20422 20644 20426 20700
rect 20426 20644 20482 20700
rect 20482 20644 20486 20700
rect 20422 20640 20486 20644
rect 27610 20700 27674 20704
rect 27610 20644 27614 20700
rect 27614 20644 27670 20700
rect 27670 20644 27674 20700
rect 27610 20640 27674 20644
rect 27690 20700 27754 20704
rect 27690 20644 27694 20700
rect 27694 20644 27750 20700
rect 27750 20644 27754 20700
rect 27690 20640 27754 20644
rect 27770 20700 27834 20704
rect 27770 20644 27774 20700
rect 27774 20644 27830 20700
rect 27830 20644 27834 20700
rect 27770 20640 27834 20644
rect 27850 20700 27914 20704
rect 27850 20644 27854 20700
rect 27854 20644 27910 20700
rect 27910 20644 27914 20700
rect 27850 20640 27914 20644
rect 4666 20156 4730 20160
rect 4666 20100 4670 20156
rect 4670 20100 4726 20156
rect 4726 20100 4730 20156
rect 4666 20096 4730 20100
rect 4746 20156 4810 20160
rect 4746 20100 4750 20156
rect 4750 20100 4806 20156
rect 4806 20100 4810 20156
rect 4746 20096 4810 20100
rect 4826 20156 4890 20160
rect 4826 20100 4830 20156
rect 4830 20100 4886 20156
rect 4886 20100 4890 20156
rect 4826 20096 4890 20100
rect 4906 20156 4970 20160
rect 4906 20100 4910 20156
rect 4910 20100 4966 20156
rect 4966 20100 4970 20156
rect 4906 20096 4970 20100
rect 12094 20156 12158 20160
rect 12094 20100 12098 20156
rect 12098 20100 12154 20156
rect 12154 20100 12158 20156
rect 12094 20096 12158 20100
rect 12174 20156 12238 20160
rect 12174 20100 12178 20156
rect 12178 20100 12234 20156
rect 12234 20100 12238 20156
rect 12174 20096 12238 20100
rect 12254 20156 12318 20160
rect 12254 20100 12258 20156
rect 12258 20100 12314 20156
rect 12314 20100 12318 20156
rect 12254 20096 12318 20100
rect 12334 20156 12398 20160
rect 12334 20100 12338 20156
rect 12338 20100 12394 20156
rect 12394 20100 12398 20156
rect 12334 20096 12398 20100
rect 19522 20156 19586 20160
rect 19522 20100 19526 20156
rect 19526 20100 19582 20156
rect 19582 20100 19586 20156
rect 19522 20096 19586 20100
rect 19602 20156 19666 20160
rect 19602 20100 19606 20156
rect 19606 20100 19662 20156
rect 19662 20100 19666 20156
rect 19602 20096 19666 20100
rect 19682 20156 19746 20160
rect 19682 20100 19686 20156
rect 19686 20100 19742 20156
rect 19742 20100 19746 20156
rect 19682 20096 19746 20100
rect 19762 20156 19826 20160
rect 19762 20100 19766 20156
rect 19766 20100 19822 20156
rect 19822 20100 19826 20156
rect 19762 20096 19826 20100
rect 26950 20156 27014 20160
rect 26950 20100 26954 20156
rect 26954 20100 27010 20156
rect 27010 20100 27014 20156
rect 26950 20096 27014 20100
rect 27030 20156 27094 20160
rect 27030 20100 27034 20156
rect 27034 20100 27090 20156
rect 27090 20100 27094 20156
rect 27030 20096 27094 20100
rect 27110 20156 27174 20160
rect 27110 20100 27114 20156
rect 27114 20100 27170 20156
rect 27170 20100 27174 20156
rect 27110 20096 27174 20100
rect 27190 20156 27254 20160
rect 27190 20100 27194 20156
rect 27194 20100 27250 20156
rect 27250 20100 27254 20156
rect 27190 20096 27254 20100
rect 5326 19612 5390 19616
rect 5326 19556 5330 19612
rect 5330 19556 5386 19612
rect 5386 19556 5390 19612
rect 5326 19552 5390 19556
rect 5406 19612 5470 19616
rect 5406 19556 5410 19612
rect 5410 19556 5466 19612
rect 5466 19556 5470 19612
rect 5406 19552 5470 19556
rect 5486 19612 5550 19616
rect 5486 19556 5490 19612
rect 5490 19556 5546 19612
rect 5546 19556 5550 19612
rect 5486 19552 5550 19556
rect 5566 19612 5630 19616
rect 5566 19556 5570 19612
rect 5570 19556 5626 19612
rect 5626 19556 5630 19612
rect 5566 19552 5630 19556
rect 12754 19612 12818 19616
rect 12754 19556 12758 19612
rect 12758 19556 12814 19612
rect 12814 19556 12818 19612
rect 12754 19552 12818 19556
rect 12834 19612 12898 19616
rect 12834 19556 12838 19612
rect 12838 19556 12894 19612
rect 12894 19556 12898 19612
rect 12834 19552 12898 19556
rect 12914 19612 12978 19616
rect 12914 19556 12918 19612
rect 12918 19556 12974 19612
rect 12974 19556 12978 19612
rect 12914 19552 12978 19556
rect 12994 19612 13058 19616
rect 12994 19556 12998 19612
rect 12998 19556 13054 19612
rect 13054 19556 13058 19612
rect 12994 19552 13058 19556
rect 20182 19612 20246 19616
rect 20182 19556 20186 19612
rect 20186 19556 20242 19612
rect 20242 19556 20246 19612
rect 20182 19552 20246 19556
rect 20262 19612 20326 19616
rect 20262 19556 20266 19612
rect 20266 19556 20322 19612
rect 20322 19556 20326 19612
rect 20262 19552 20326 19556
rect 20342 19612 20406 19616
rect 20342 19556 20346 19612
rect 20346 19556 20402 19612
rect 20402 19556 20406 19612
rect 20342 19552 20406 19556
rect 20422 19612 20486 19616
rect 20422 19556 20426 19612
rect 20426 19556 20482 19612
rect 20482 19556 20486 19612
rect 20422 19552 20486 19556
rect 27610 19612 27674 19616
rect 27610 19556 27614 19612
rect 27614 19556 27670 19612
rect 27670 19556 27674 19612
rect 27610 19552 27674 19556
rect 27690 19612 27754 19616
rect 27690 19556 27694 19612
rect 27694 19556 27750 19612
rect 27750 19556 27754 19612
rect 27690 19552 27754 19556
rect 27770 19612 27834 19616
rect 27770 19556 27774 19612
rect 27774 19556 27830 19612
rect 27830 19556 27834 19612
rect 27770 19552 27834 19556
rect 27850 19612 27914 19616
rect 27850 19556 27854 19612
rect 27854 19556 27910 19612
rect 27910 19556 27914 19612
rect 27850 19552 27914 19556
rect 4666 19068 4730 19072
rect 4666 19012 4670 19068
rect 4670 19012 4726 19068
rect 4726 19012 4730 19068
rect 4666 19008 4730 19012
rect 4746 19068 4810 19072
rect 4746 19012 4750 19068
rect 4750 19012 4806 19068
rect 4806 19012 4810 19068
rect 4746 19008 4810 19012
rect 4826 19068 4890 19072
rect 4826 19012 4830 19068
rect 4830 19012 4886 19068
rect 4886 19012 4890 19068
rect 4826 19008 4890 19012
rect 4906 19068 4970 19072
rect 4906 19012 4910 19068
rect 4910 19012 4966 19068
rect 4966 19012 4970 19068
rect 4906 19008 4970 19012
rect 12094 19068 12158 19072
rect 12094 19012 12098 19068
rect 12098 19012 12154 19068
rect 12154 19012 12158 19068
rect 12094 19008 12158 19012
rect 12174 19068 12238 19072
rect 12174 19012 12178 19068
rect 12178 19012 12234 19068
rect 12234 19012 12238 19068
rect 12174 19008 12238 19012
rect 12254 19068 12318 19072
rect 12254 19012 12258 19068
rect 12258 19012 12314 19068
rect 12314 19012 12318 19068
rect 12254 19008 12318 19012
rect 12334 19068 12398 19072
rect 12334 19012 12338 19068
rect 12338 19012 12394 19068
rect 12394 19012 12398 19068
rect 12334 19008 12398 19012
rect 19522 19068 19586 19072
rect 19522 19012 19526 19068
rect 19526 19012 19582 19068
rect 19582 19012 19586 19068
rect 19522 19008 19586 19012
rect 19602 19068 19666 19072
rect 19602 19012 19606 19068
rect 19606 19012 19662 19068
rect 19662 19012 19666 19068
rect 19602 19008 19666 19012
rect 19682 19068 19746 19072
rect 19682 19012 19686 19068
rect 19686 19012 19742 19068
rect 19742 19012 19746 19068
rect 19682 19008 19746 19012
rect 19762 19068 19826 19072
rect 19762 19012 19766 19068
rect 19766 19012 19822 19068
rect 19822 19012 19826 19068
rect 19762 19008 19826 19012
rect 26950 19068 27014 19072
rect 26950 19012 26954 19068
rect 26954 19012 27010 19068
rect 27010 19012 27014 19068
rect 26950 19008 27014 19012
rect 27030 19068 27094 19072
rect 27030 19012 27034 19068
rect 27034 19012 27090 19068
rect 27090 19012 27094 19068
rect 27030 19008 27094 19012
rect 27110 19068 27174 19072
rect 27110 19012 27114 19068
rect 27114 19012 27170 19068
rect 27170 19012 27174 19068
rect 27110 19008 27174 19012
rect 27190 19068 27254 19072
rect 27190 19012 27194 19068
rect 27194 19012 27250 19068
rect 27250 19012 27254 19068
rect 27190 19008 27254 19012
rect 5326 18524 5390 18528
rect 5326 18468 5330 18524
rect 5330 18468 5386 18524
rect 5386 18468 5390 18524
rect 5326 18464 5390 18468
rect 5406 18524 5470 18528
rect 5406 18468 5410 18524
rect 5410 18468 5466 18524
rect 5466 18468 5470 18524
rect 5406 18464 5470 18468
rect 5486 18524 5550 18528
rect 5486 18468 5490 18524
rect 5490 18468 5546 18524
rect 5546 18468 5550 18524
rect 5486 18464 5550 18468
rect 5566 18524 5630 18528
rect 5566 18468 5570 18524
rect 5570 18468 5626 18524
rect 5626 18468 5630 18524
rect 5566 18464 5630 18468
rect 12754 18524 12818 18528
rect 12754 18468 12758 18524
rect 12758 18468 12814 18524
rect 12814 18468 12818 18524
rect 12754 18464 12818 18468
rect 12834 18524 12898 18528
rect 12834 18468 12838 18524
rect 12838 18468 12894 18524
rect 12894 18468 12898 18524
rect 12834 18464 12898 18468
rect 12914 18524 12978 18528
rect 12914 18468 12918 18524
rect 12918 18468 12974 18524
rect 12974 18468 12978 18524
rect 12914 18464 12978 18468
rect 12994 18524 13058 18528
rect 12994 18468 12998 18524
rect 12998 18468 13054 18524
rect 13054 18468 13058 18524
rect 12994 18464 13058 18468
rect 20182 18524 20246 18528
rect 20182 18468 20186 18524
rect 20186 18468 20242 18524
rect 20242 18468 20246 18524
rect 20182 18464 20246 18468
rect 20262 18524 20326 18528
rect 20262 18468 20266 18524
rect 20266 18468 20322 18524
rect 20322 18468 20326 18524
rect 20262 18464 20326 18468
rect 20342 18524 20406 18528
rect 20342 18468 20346 18524
rect 20346 18468 20402 18524
rect 20402 18468 20406 18524
rect 20342 18464 20406 18468
rect 20422 18524 20486 18528
rect 20422 18468 20426 18524
rect 20426 18468 20482 18524
rect 20482 18468 20486 18524
rect 20422 18464 20486 18468
rect 27610 18524 27674 18528
rect 27610 18468 27614 18524
rect 27614 18468 27670 18524
rect 27670 18468 27674 18524
rect 27610 18464 27674 18468
rect 27690 18524 27754 18528
rect 27690 18468 27694 18524
rect 27694 18468 27750 18524
rect 27750 18468 27754 18524
rect 27690 18464 27754 18468
rect 27770 18524 27834 18528
rect 27770 18468 27774 18524
rect 27774 18468 27830 18524
rect 27830 18468 27834 18524
rect 27770 18464 27834 18468
rect 27850 18524 27914 18528
rect 27850 18468 27854 18524
rect 27854 18468 27910 18524
rect 27910 18468 27914 18524
rect 27850 18464 27914 18468
rect 4666 17980 4730 17984
rect 4666 17924 4670 17980
rect 4670 17924 4726 17980
rect 4726 17924 4730 17980
rect 4666 17920 4730 17924
rect 4746 17980 4810 17984
rect 4746 17924 4750 17980
rect 4750 17924 4806 17980
rect 4806 17924 4810 17980
rect 4746 17920 4810 17924
rect 4826 17980 4890 17984
rect 4826 17924 4830 17980
rect 4830 17924 4886 17980
rect 4886 17924 4890 17980
rect 4826 17920 4890 17924
rect 4906 17980 4970 17984
rect 4906 17924 4910 17980
rect 4910 17924 4966 17980
rect 4966 17924 4970 17980
rect 4906 17920 4970 17924
rect 12094 17980 12158 17984
rect 12094 17924 12098 17980
rect 12098 17924 12154 17980
rect 12154 17924 12158 17980
rect 12094 17920 12158 17924
rect 12174 17980 12238 17984
rect 12174 17924 12178 17980
rect 12178 17924 12234 17980
rect 12234 17924 12238 17980
rect 12174 17920 12238 17924
rect 12254 17980 12318 17984
rect 12254 17924 12258 17980
rect 12258 17924 12314 17980
rect 12314 17924 12318 17980
rect 12254 17920 12318 17924
rect 12334 17980 12398 17984
rect 12334 17924 12338 17980
rect 12338 17924 12394 17980
rect 12394 17924 12398 17980
rect 12334 17920 12398 17924
rect 19522 17980 19586 17984
rect 19522 17924 19526 17980
rect 19526 17924 19582 17980
rect 19582 17924 19586 17980
rect 19522 17920 19586 17924
rect 19602 17980 19666 17984
rect 19602 17924 19606 17980
rect 19606 17924 19662 17980
rect 19662 17924 19666 17980
rect 19602 17920 19666 17924
rect 19682 17980 19746 17984
rect 19682 17924 19686 17980
rect 19686 17924 19742 17980
rect 19742 17924 19746 17980
rect 19682 17920 19746 17924
rect 19762 17980 19826 17984
rect 19762 17924 19766 17980
rect 19766 17924 19822 17980
rect 19822 17924 19826 17980
rect 19762 17920 19826 17924
rect 26950 17980 27014 17984
rect 26950 17924 26954 17980
rect 26954 17924 27010 17980
rect 27010 17924 27014 17980
rect 26950 17920 27014 17924
rect 27030 17980 27094 17984
rect 27030 17924 27034 17980
rect 27034 17924 27090 17980
rect 27090 17924 27094 17980
rect 27030 17920 27094 17924
rect 27110 17980 27174 17984
rect 27110 17924 27114 17980
rect 27114 17924 27170 17980
rect 27170 17924 27174 17980
rect 27110 17920 27174 17924
rect 27190 17980 27254 17984
rect 27190 17924 27194 17980
rect 27194 17924 27250 17980
rect 27250 17924 27254 17980
rect 27190 17920 27254 17924
rect 5326 17436 5390 17440
rect 5326 17380 5330 17436
rect 5330 17380 5386 17436
rect 5386 17380 5390 17436
rect 5326 17376 5390 17380
rect 5406 17436 5470 17440
rect 5406 17380 5410 17436
rect 5410 17380 5466 17436
rect 5466 17380 5470 17436
rect 5406 17376 5470 17380
rect 5486 17436 5550 17440
rect 5486 17380 5490 17436
rect 5490 17380 5546 17436
rect 5546 17380 5550 17436
rect 5486 17376 5550 17380
rect 5566 17436 5630 17440
rect 5566 17380 5570 17436
rect 5570 17380 5626 17436
rect 5626 17380 5630 17436
rect 5566 17376 5630 17380
rect 12754 17436 12818 17440
rect 12754 17380 12758 17436
rect 12758 17380 12814 17436
rect 12814 17380 12818 17436
rect 12754 17376 12818 17380
rect 12834 17436 12898 17440
rect 12834 17380 12838 17436
rect 12838 17380 12894 17436
rect 12894 17380 12898 17436
rect 12834 17376 12898 17380
rect 12914 17436 12978 17440
rect 12914 17380 12918 17436
rect 12918 17380 12974 17436
rect 12974 17380 12978 17436
rect 12914 17376 12978 17380
rect 12994 17436 13058 17440
rect 12994 17380 12998 17436
rect 12998 17380 13054 17436
rect 13054 17380 13058 17436
rect 12994 17376 13058 17380
rect 20182 17436 20246 17440
rect 20182 17380 20186 17436
rect 20186 17380 20242 17436
rect 20242 17380 20246 17436
rect 20182 17376 20246 17380
rect 20262 17436 20326 17440
rect 20262 17380 20266 17436
rect 20266 17380 20322 17436
rect 20322 17380 20326 17436
rect 20262 17376 20326 17380
rect 20342 17436 20406 17440
rect 20342 17380 20346 17436
rect 20346 17380 20402 17436
rect 20402 17380 20406 17436
rect 20342 17376 20406 17380
rect 20422 17436 20486 17440
rect 20422 17380 20426 17436
rect 20426 17380 20482 17436
rect 20482 17380 20486 17436
rect 20422 17376 20486 17380
rect 27610 17436 27674 17440
rect 27610 17380 27614 17436
rect 27614 17380 27670 17436
rect 27670 17380 27674 17436
rect 27610 17376 27674 17380
rect 27690 17436 27754 17440
rect 27690 17380 27694 17436
rect 27694 17380 27750 17436
rect 27750 17380 27754 17436
rect 27690 17376 27754 17380
rect 27770 17436 27834 17440
rect 27770 17380 27774 17436
rect 27774 17380 27830 17436
rect 27830 17380 27834 17436
rect 27770 17376 27834 17380
rect 27850 17436 27914 17440
rect 27850 17380 27854 17436
rect 27854 17380 27910 17436
rect 27910 17380 27914 17436
rect 27850 17376 27914 17380
rect 4666 16892 4730 16896
rect 4666 16836 4670 16892
rect 4670 16836 4726 16892
rect 4726 16836 4730 16892
rect 4666 16832 4730 16836
rect 4746 16892 4810 16896
rect 4746 16836 4750 16892
rect 4750 16836 4806 16892
rect 4806 16836 4810 16892
rect 4746 16832 4810 16836
rect 4826 16892 4890 16896
rect 4826 16836 4830 16892
rect 4830 16836 4886 16892
rect 4886 16836 4890 16892
rect 4826 16832 4890 16836
rect 4906 16892 4970 16896
rect 4906 16836 4910 16892
rect 4910 16836 4966 16892
rect 4966 16836 4970 16892
rect 4906 16832 4970 16836
rect 12094 16892 12158 16896
rect 12094 16836 12098 16892
rect 12098 16836 12154 16892
rect 12154 16836 12158 16892
rect 12094 16832 12158 16836
rect 12174 16892 12238 16896
rect 12174 16836 12178 16892
rect 12178 16836 12234 16892
rect 12234 16836 12238 16892
rect 12174 16832 12238 16836
rect 12254 16892 12318 16896
rect 12254 16836 12258 16892
rect 12258 16836 12314 16892
rect 12314 16836 12318 16892
rect 12254 16832 12318 16836
rect 12334 16892 12398 16896
rect 12334 16836 12338 16892
rect 12338 16836 12394 16892
rect 12394 16836 12398 16892
rect 12334 16832 12398 16836
rect 19522 16892 19586 16896
rect 19522 16836 19526 16892
rect 19526 16836 19582 16892
rect 19582 16836 19586 16892
rect 19522 16832 19586 16836
rect 19602 16892 19666 16896
rect 19602 16836 19606 16892
rect 19606 16836 19662 16892
rect 19662 16836 19666 16892
rect 19602 16832 19666 16836
rect 19682 16892 19746 16896
rect 19682 16836 19686 16892
rect 19686 16836 19742 16892
rect 19742 16836 19746 16892
rect 19682 16832 19746 16836
rect 19762 16892 19826 16896
rect 19762 16836 19766 16892
rect 19766 16836 19822 16892
rect 19822 16836 19826 16892
rect 19762 16832 19826 16836
rect 26950 16892 27014 16896
rect 26950 16836 26954 16892
rect 26954 16836 27010 16892
rect 27010 16836 27014 16892
rect 26950 16832 27014 16836
rect 27030 16892 27094 16896
rect 27030 16836 27034 16892
rect 27034 16836 27090 16892
rect 27090 16836 27094 16892
rect 27030 16832 27094 16836
rect 27110 16892 27174 16896
rect 27110 16836 27114 16892
rect 27114 16836 27170 16892
rect 27170 16836 27174 16892
rect 27110 16832 27174 16836
rect 27190 16892 27254 16896
rect 27190 16836 27194 16892
rect 27194 16836 27250 16892
rect 27250 16836 27254 16892
rect 27190 16832 27254 16836
rect 5326 16348 5390 16352
rect 5326 16292 5330 16348
rect 5330 16292 5386 16348
rect 5386 16292 5390 16348
rect 5326 16288 5390 16292
rect 5406 16348 5470 16352
rect 5406 16292 5410 16348
rect 5410 16292 5466 16348
rect 5466 16292 5470 16348
rect 5406 16288 5470 16292
rect 5486 16348 5550 16352
rect 5486 16292 5490 16348
rect 5490 16292 5546 16348
rect 5546 16292 5550 16348
rect 5486 16288 5550 16292
rect 5566 16348 5630 16352
rect 5566 16292 5570 16348
rect 5570 16292 5626 16348
rect 5626 16292 5630 16348
rect 5566 16288 5630 16292
rect 12754 16348 12818 16352
rect 12754 16292 12758 16348
rect 12758 16292 12814 16348
rect 12814 16292 12818 16348
rect 12754 16288 12818 16292
rect 12834 16348 12898 16352
rect 12834 16292 12838 16348
rect 12838 16292 12894 16348
rect 12894 16292 12898 16348
rect 12834 16288 12898 16292
rect 12914 16348 12978 16352
rect 12914 16292 12918 16348
rect 12918 16292 12974 16348
rect 12974 16292 12978 16348
rect 12914 16288 12978 16292
rect 12994 16348 13058 16352
rect 12994 16292 12998 16348
rect 12998 16292 13054 16348
rect 13054 16292 13058 16348
rect 12994 16288 13058 16292
rect 20182 16348 20246 16352
rect 20182 16292 20186 16348
rect 20186 16292 20242 16348
rect 20242 16292 20246 16348
rect 20182 16288 20246 16292
rect 20262 16348 20326 16352
rect 20262 16292 20266 16348
rect 20266 16292 20322 16348
rect 20322 16292 20326 16348
rect 20262 16288 20326 16292
rect 20342 16348 20406 16352
rect 20342 16292 20346 16348
rect 20346 16292 20402 16348
rect 20402 16292 20406 16348
rect 20342 16288 20406 16292
rect 20422 16348 20486 16352
rect 20422 16292 20426 16348
rect 20426 16292 20482 16348
rect 20482 16292 20486 16348
rect 20422 16288 20486 16292
rect 27610 16348 27674 16352
rect 27610 16292 27614 16348
rect 27614 16292 27670 16348
rect 27670 16292 27674 16348
rect 27610 16288 27674 16292
rect 27690 16348 27754 16352
rect 27690 16292 27694 16348
rect 27694 16292 27750 16348
rect 27750 16292 27754 16348
rect 27690 16288 27754 16292
rect 27770 16348 27834 16352
rect 27770 16292 27774 16348
rect 27774 16292 27830 16348
rect 27830 16292 27834 16348
rect 27770 16288 27834 16292
rect 27850 16348 27914 16352
rect 27850 16292 27854 16348
rect 27854 16292 27910 16348
rect 27910 16292 27914 16348
rect 27850 16288 27914 16292
rect 4666 15804 4730 15808
rect 4666 15748 4670 15804
rect 4670 15748 4726 15804
rect 4726 15748 4730 15804
rect 4666 15744 4730 15748
rect 4746 15804 4810 15808
rect 4746 15748 4750 15804
rect 4750 15748 4806 15804
rect 4806 15748 4810 15804
rect 4746 15744 4810 15748
rect 4826 15804 4890 15808
rect 4826 15748 4830 15804
rect 4830 15748 4886 15804
rect 4886 15748 4890 15804
rect 4826 15744 4890 15748
rect 4906 15804 4970 15808
rect 4906 15748 4910 15804
rect 4910 15748 4966 15804
rect 4966 15748 4970 15804
rect 4906 15744 4970 15748
rect 12094 15804 12158 15808
rect 12094 15748 12098 15804
rect 12098 15748 12154 15804
rect 12154 15748 12158 15804
rect 12094 15744 12158 15748
rect 12174 15804 12238 15808
rect 12174 15748 12178 15804
rect 12178 15748 12234 15804
rect 12234 15748 12238 15804
rect 12174 15744 12238 15748
rect 12254 15804 12318 15808
rect 12254 15748 12258 15804
rect 12258 15748 12314 15804
rect 12314 15748 12318 15804
rect 12254 15744 12318 15748
rect 12334 15804 12398 15808
rect 12334 15748 12338 15804
rect 12338 15748 12394 15804
rect 12394 15748 12398 15804
rect 12334 15744 12398 15748
rect 19522 15804 19586 15808
rect 19522 15748 19526 15804
rect 19526 15748 19582 15804
rect 19582 15748 19586 15804
rect 19522 15744 19586 15748
rect 19602 15804 19666 15808
rect 19602 15748 19606 15804
rect 19606 15748 19662 15804
rect 19662 15748 19666 15804
rect 19602 15744 19666 15748
rect 19682 15804 19746 15808
rect 19682 15748 19686 15804
rect 19686 15748 19742 15804
rect 19742 15748 19746 15804
rect 19682 15744 19746 15748
rect 19762 15804 19826 15808
rect 19762 15748 19766 15804
rect 19766 15748 19822 15804
rect 19822 15748 19826 15804
rect 19762 15744 19826 15748
rect 26950 15804 27014 15808
rect 26950 15748 26954 15804
rect 26954 15748 27010 15804
rect 27010 15748 27014 15804
rect 26950 15744 27014 15748
rect 27030 15804 27094 15808
rect 27030 15748 27034 15804
rect 27034 15748 27090 15804
rect 27090 15748 27094 15804
rect 27030 15744 27094 15748
rect 27110 15804 27174 15808
rect 27110 15748 27114 15804
rect 27114 15748 27170 15804
rect 27170 15748 27174 15804
rect 27110 15744 27174 15748
rect 27190 15804 27254 15808
rect 27190 15748 27194 15804
rect 27194 15748 27250 15804
rect 27250 15748 27254 15804
rect 27190 15744 27254 15748
rect 5326 15260 5390 15264
rect 5326 15204 5330 15260
rect 5330 15204 5386 15260
rect 5386 15204 5390 15260
rect 5326 15200 5390 15204
rect 5406 15260 5470 15264
rect 5406 15204 5410 15260
rect 5410 15204 5466 15260
rect 5466 15204 5470 15260
rect 5406 15200 5470 15204
rect 5486 15260 5550 15264
rect 5486 15204 5490 15260
rect 5490 15204 5546 15260
rect 5546 15204 5550 15260
rect 5486 15200 5550 15204
rect 5566 15260 5630 15264
rect 5566 15204 5570 15260
rect 5570 15204 5626 15260
rect 5626 15204 5630 15260
rect 5566 15200 5630 15204
rect 12754 15260 12818 15264
rect 12754 15204 12758 15260
rect 12758 15204 12814 15260
rect 12814 15204 12818 15260
rect 12754 15200 12818 15204
rect 12834 15260 12898 15264
rect 12834 15204 12838 15260
rect 12838 15204 12894 15260
rect 12894 15204 12898 15260
rect 12834 15200 12898 15204
rect 12914 15260 12978 15264
rect 12914 15204 12918 15260
rect 12918 15204 12974 15260
rect 12974 15204 12978 15260
rect 12914 15200 12978 15204
rect 12994 15260 13058 15264
rect 12994 15204 12998 15260
rect 12998 15204 13054 15260
rect 13054 15204 13058 15260
rect 12994 15200 13058 15204
rect 20182 15260 20246 15264
rect 20182 15204 20186 15260
rect 20186 15204 20242 15260
rect 20242 15204 20246 15260
rect 20182 15200 20246 15204
rect 20262 15260 20326 15264
rect 20262 15204 20266 15260
rect 20266 15204 20322 15260
rect 20322 15204 20326 15260
rect 20262 15200 20326 15204
rect 20342 15260 20406 15264
rect 20342 15204 20346 15260
rect 20346 15204 20402 15260
rect 20402 15204 20406 15260
rect 20342 15200 20406 15204
rect 20422 15260 20486 15264
rect 20422 15204 20426 15260
rect 20426 15204 20482 15260
rect 20482 15204 20486 15260
rect 20422 15200 20486 15204
rect 27610 15260 27674 15264
rect 27610 15204 27614 15260
rect 27614 15204 27670 15260
rect 27670 15204 27674 15260
rect 27610 15200 27674 15204
rect 27690 15260 27754 15264
rect 27690 15204 27694 15260
rect 27694 15204 27750 15260
rect 27750 15204 27754 15260
rect 27690 15200 27754 15204
rect 27770 15260 27834 15264
rect 27770 15204 27774 15260
rect 27774 15204 27830 15260
rect 27830 15204 27834 15260
rect 27770 15200 27834 15204
rect 27850 15260 27914 15264
rect 27850 15204 27854 15260
rect 27854 15204 27910 15260
rect 27910 15204 27914 15260
rect 27850 15200 27914 15204
rect 4666 14716 4730 14720
rect 4666 14660 4670 14716
rect 4670 14660 4726 14716
rect 4726 14660 4730 14716
rect 4666 14656 4730 14660
rect 4746 14716 4810 14720
rect 4746 14660 4750 14716
rect 4750 14660 4806 14716
rect 4806 14660 4810 14716
rect 4746 14656 4810 14660
rect 4826 14716 4890 14720
rect 4826 14660 4830 14716
rect 4830 14660 4886 14716
rect 4886 14660 4890 14716
rect 4826 14656 4890 14660
rect 4906 14716 4970 14720
rect 4906 14660 4910 14716
rect 4910 14660 4966 14716
rect 4966 14660 4970 14716
rect 4906 14656 4970 14660
rect 12094 14716 12158 14720
rect 12094 14660 12098 14716
rect 12098 14660 12154 14716
rect 12154 14660 12158 14716
rect 12094 14656 12158 14660
rect 12174 14716 12238 14720
rect 12174 14660 12178 14716
rect 12178 14660 12234 14716
rect 12234 14660 12238 14716
rect 12174 14656 12238 14660
rect 12254 14716 12318 14720
rect 12254 14660 12258 14716
rect 12258 14660 12314 14716
rect 12314 14660 12318 14716
rect 12254 14656 12318 14660
rect 12334 14716 12398 14720
rect 12334 14660 12338 14716
rect 12338 14660 12394 14716
rect 12394 14660 12398 14716
rect 12334 14656 12398 14660
rect 19522 14716 19586 14720
rect 19522 14660 19526 14716
rect 19526 14660 19582 14716
rect 19582 14660 19586 14716
rect 19522 14656 19586 14660
rect 19602 14716 19666 14720
rect 19602 14660 19606 14716
rect 19606 14660 19662 14716
rect 19662 14660 19666 14716
rect 19602 14656 19666 14660
rect 19682 14716 19746 14720
rect 19682 14660 19686 14716
rect 19686 14660 19742 14716
rect 19742 14660 19746 14716
rect 19682 14656 19746 14660
rect 19762 14716 19826 14720
rect 19762 14660 19766 14716
rect 19766 14660 19822 14716
rect 19822 14660 19826 14716
rect 19762 14656 19826 14660
rect 26950 14716 27014 14720
rect 26950 14660 26954 14716
rect 26954 14660 27010 14716
rect 27010 14660 27014 14716
rect 26950 14656 27014 14660
rect 27030 14716 27094 14720
rect 27030 14660 27034 14716
rect 27034 14660 27090 14716
rect 27090 14660 27094 14716
rect 27030 14656 27094 14660
rect 27110 14716 27174 14720
rect 27110 14660 27114 14716
rect 27114 14660 27170 14716
rect 27170 14660 27174 14716
rect 27110 14656 27174 14660
rect 27190 14716 27254 14720
rect 27190 14660 27194 14716
rect 27194 14660 27250 14716
rect 27250 14660 27254 14716
rect 27190 14656 27254 14660
rect 5326 14172 5390 14176
rect 5326 14116 5330 14172
rect 5330 14116 5386 14172
rect 5386 14116 5390 14172
rect 5326 14112 5390 14116
rect 5406 14172 5470 14176
rect 5406 14116 5410 14172
rect 5410 14116 5466 14172
rect 5466 14116 5470 14172
rect 5406 14112 5470 14116
rect 5486 14172 5550 14176
rect 5486 14116 5490 14172
rect 5490 14116 5546 14172
rect 5546 14116 5550 14172
rect 5486 14112 5550 14116
rect 5566 14172 5630 14176
rect 5566 14116 5570 14172
rect 5570 14116 5626 14172
rect 5626 14116 5630 14172
rect 5566 14112 5630 14116
rect 12754 14172 12818 14176
rect 12754 14116 12758 14172
rect 12758 14116 12814 14172
rect 12814 14116 12818 14172
rect 12754 14112 12818 14116
rect 12834 14172 12898 14176
rect 12834 14116 12838 14172
rect 12838 14116 12894 14172
rect 12894 14116 12898 14172
rect 12834 14112 12898 14116
rect 12914 14172 12978 14176
rect 12914 14116 12918 14172
rect 12918 14116 12974 14172
rect 12974 14116 12978 14172
rect 12914 14112 12978 14116
rect 12994 14172 13058 14176
rect 12994 14116 12998 14172
rect 12998 14116 13054 14172
rect 13054 14116 13058 14172
rect 12994 14112 13058 14116
rect 20182 14172 20246 14176
rect 20182 14116 20186 14172
rect 20186 14116 20242 14172
rect 20242 14116 20246 14172
rect 20182 14112 20246 14116
rect 20262 14172 20326 14176
rect 20262 14116 20266 14172
rect 20266 14116 20322 14172
rect 20322 14116 20326 14172
rect 20262 14112 20326 14116
rect 20342 14172 20406 14176
rect 20342 14116 20346 14172
rect 20346 14116 20402 14172
rect 20402 14116 20406 14172
rect 20342 14112 20406 14116
rect 20422 14172 20486 14176
rect 20422 14116 20426 14172
rect 20426 14116 20482 14172
rect 20482 14116 20486 14172
rect 20422 14112 20486 14116
rect 27610 14172 27674 14176
rect 27610 14116 27614 14172
rect 27614 14116 27670 14172
rect 27670 14116 27674 14172
rect 27610 14112 27674 14116
rect 27690 14172 27754 14176
rect 27690 14116 27694 14172
rect 27694 14116 27750 14172
rect 27750 14116 27754 14172
rect 27690 14112 27754 14116
rect 27770 14172 27834 14176
rect 27770 14116 27774 14172
rect 27774 14116 27830 14172
rect 27830 14116 27834 14172
rect 27770 14112 27834 14116
rect 27850 14172 27914 14176
rect 27850 14116 27854 14172
rect 27854 14116 27910 14172
rect 27910 14116 27914 14172
rect 27850 14112 27914 14116
rect 4666 13628 4730 13632
rect 4666 13572 4670 13628
rect 4670 13572 4726 13628
rect 4726 13572 4730 13628
rect 4666 13568 4730 13572
rect 4746 13628 4810 13632
rect 4746 13572 4750 13628
rect 4750 13572 4806 13628
rect 4806 13572 4810 13628
rect 4746 13568 4810 13572
rect 4826 13628 4890 13632
rect 4826 13572 4830 13628
rect 4830 13572 4886 13628
rect 4886 13572 4890 13628
rect 4826 13568 4890 13572
rect 4906 13628 4970 13632
rect 4906 13572 4910 13628
rect 4910 13572 4966 13628
rect 4966 13572 4970 13628
rect 4906 13568 4970 13572
rect 12094 13628 12158 13632
rect 12094 13572 12098 13628
rect 12098 13572 12154 13628
rect 12154 13572 12158 13628
rect 12094 13568 12158 13572
rect 12174 13628 12238 13632
rect 12174 13572 12178 13628
rect 12178 13572 12234 13628
rect 12234 13572 12238 13628
rect 12174 13568 12238 13572
rect 12254 13628 12318 13632
rect 12254 13572 12258 13628
rect 12258 13572 12314 13628
rect 12314 13572 12318 13628
rect 12254 13568 12318 13572
rect 12334 13628 12398 13632
rect 12334 13572 12338 13628
rect 12338 13572 12394 13628
rect 12394 13572 12398 13628
rect 12334 13568 12398 13572
rect 19522 13628 19586 13632
rect 19522 13572 19526 13628
rect 19526 13572 19582 13628
rect 19582 13572 19586 13628
rect 19522 13568 19586 13572
rect 19602 13628 19666 13632
rect 19602 13572 19606 13628
rect 19606 13572 19662 13628
rect 19662 13572 19666 13628
rect 19602 13568 19666 13572
rect 19682 13628 19746 13632
rect 19682 13572 19686 13628
rect 19686 13572 19742 13628
rect 19742 13572 19746 13628
rect 19682 13568 19746 13572
rect 19762 13628 19826 13632
rect 19762 13572 19766 13628
rect 19766 13572 19822 13628
rect 19822 13572 19826 13628
rect 19762 13568 19826 13572
rect 26950 13628 27014 13632
rect 26950 13572 26954 13628
rect 26954 13572 27010 13628
rect 27010 13572 27014 13628
rect 26950 13568 27014 13572
rect 27030 13628 27094 13632
rect 27030 13572 27034 13628
rect 27034 13572 27090 13628
rect 27090 13572 27094 13628
rect 27030 13568 27094 13572
rect 27110 13628 27174 13632
rect 27110 13572 27114 13628
rect 27114 13572 27170 13628
rect 27170 13572 27174 13628
rect 27110 13568 27174 13572
rect 27190 13628 27254 13632
rect 27190 13572 27194 13628
rect 27194 13572 27250 13628
rect 27250 13572 27254 13628
rect 27190 13568 27254 13572
rect 5326 13084 5390 13088
rect 5326 13028 5330 13084
rect 5330 13028 5386 13084
rect 5386 13028 5390 13084
rect 5326 13024 5390 13028
rect 5406 13084 5470 13088
rect 5406 13028 5410 13084
rect 5410 13028 5466 13084
rect 5466 13028 5470 13084
rect 5406 13024 5470 13028
rect 5486 13084 5550 13088
rect 5486 13028 5490 13084
rect 5490 13028 5546 13084
rect 5546 13028 5550 13084
rect 5486 13024 5550 13028
rect 5566 13084 5630 13088
rect 5566 13028 5570 13084
rect 5570 13028 5626 13084
rect 5626 13028 5630 13084
rect 5566 13024 5630 13028
rect 12754 13084 12818 13088
rect 12754 13028 12758 13084
rect 12758 13028 12814 13084
rect 12814 13028 12818 13084
rect 12754 13024 12818 13028
rect 12834 13084 12898 13088
rect 12834 13028 12838 13084
rect 12838 13028 12894 13084
rect 12894 13028 12898 13084
rect 12834 13024 12898 13028
rect 12914 13084 12978 13088
rect 12914 13028 12918 13084
rect 12918 13028 12974 13084
rect 12974 13028 12978 13084
rect 12914 13024 12978 13028
rect 12994 13084 13058 13088
rect 12994 13028 12998 13084
rect 12998 13028 13054 13084
rect 13054 13028 13058 13084
rect 12994 13024 13058 13028
rect 20182 13084 20246 13088
rect 20182 13028 20186 13084
rect 20186 13028 20242 13084
rect 20242 13028 20246 13084
rect 20182 13024 20246 13028
rect 20262 13084 20326 13088
rect 20262 13028 20266 13084
rect 20266 13028 20322 13084
rect 20322 13028 20326 13084
rect 20262 13024 20326 13028
rect 20342 13084 20406 13088
rect 20342 13028 20346 13084
rect 20346 13028 20402 13084
rect 20402 13028 20406 13084
rect 20342 13024 20406 13028
rect 20422 13084 20486 13088
rect 20422 13028 20426 13084
rect 20426 13028 20482 13084
rect 20482 13028 20486 13084
rect 20422 13024 20486 13028
rect 27610 13084 27674 13088
rect 27610 13028 27614 13084
rect 27614 13028 27670 13084
rect 27670 13028 27674 13084
rect 27610 13024 27674 13028
rect 27690 13084 27754 13088
rect 27690 13028 27694 13084
rect 27694 13028 27750 13084
rect 27750 13028 27754 13084
rect 27690 13024 27754 13028
rect 27770 13084 27834 13088
rect 27770 13028 27774 13084
rect 27774 13028 27830 13084
rect 27830 13028 27834 13084
rect 27770 13024 27834 13028
rect 27850 13084 27914 13088
rect 27850 13028 27854 13084
rect 27854 13028 27910 13084
rect 27910 13028 27914 13084
rect 27850 13024 27914 13028
rect 4666 12540 4730 12544
rect 4666 12484 4670 12540
rect 4670 12484 4726 12540
rect 4726 12484 4730 12540
rect 4666 12480 4730 12484
rect 4746 12540 4810 12544
rect 4746 12484 4750 12540
rect 4750 12484 4806 12540
rect 4806 12484 4810 12540
rect 4746 12480 4810 12484
rect 4826 12540 4890 12544
rect 4826 12484 4830 12540
rect 4830 12484 4886 12540
rect 4886 12484 4890 12540
rect 4826 12480 4890 12484
rect 4906 12540 4970 12544
rect 4906 12484 4910 12540
rect 4910 12484 4966 12540
rect 4966 12484 4970 12540
rect 4906 12480 4970 12484
rect 12094 12540 12158 12544
rect 12094 12484 12098 12540
rect 12098 12484 12154 12540
rect 12154 12484 12158 12540
rect 12094 12480 12158 12484
rect 12174 12540 12238 12544
rect 12174 12484 12178 12540
rect 12178 12484 12234 12540
rect 12234 12484 12238 12540
rect 12174 12480 12238 12484
rect 12254 12540 12318 12544
rect 12254 12484 12258 12540
rect 12258 12484 12314 12540
rect 12314 12484 12318 12540
rect 12254 12480 12318 12484
rect 12334 12540 12398 12544
rect 12334 12484 12338 12540
rect 12338 12484 12394 12540
rect 12394 12484 12398 12540
rect 12334 12480 12398 12484
rect 19522 12540 19586 12544
rect 19522 12484 19526 12540
rect 19526 12484 19582 12540
rect 19582 12484 19586 12540
rect 19522 12480 19586 12484
rect 19602 12540 19666 12544
rect 19602 12484 19606 12540
rect 19606 12484 19662 12540
rect 19662 12484 19666 12540
rect 19602 12480 19666 12484
rect 19682 12540 19746 12544
rect 19682 12484 19686 12540
rect 19686 12484 19742 12540
rect 19742 12484 19746 12540
rect 19682 12480 19746 12484
rect 19762 12540 19826 12544
rect 19762 12484 19766 12540
rect 19766 12484 19822 12540
rect 19822 12484 19826 12540
rect 19762 12480 19826 12484
rect 26950 12540 27014 12544
rect 26950 12484 26954 12540
rect 26954 12484 27010 12540
rect 27010 12484 27014 12540
rect 26950 12480 27014 12484
rect 27030 12540 27094 12544
rect 27030 12484 27034 12540
rect 27034 12484 27090 12540
rect 27090 12484 27094 12540
rect 27030 12480 27094 12484
rect 27110 12540 27174 12544
rect 27110 12484 27114 12540
rect 27114 12484 27170 12540
rect 27170 12484 27174 12540
rect 27110 12480 27174 12484
rect 27190 12540 27254 12544
rect 27190 12484 27194 12540
rect 27194 12484 27250 12540
rect 27250 12484 27254 12540
rect 27190 12480 27254 12484
rect 5326 11996 5390 12000
rect 5326 11940 5330 11996
rect 5330 11940 5386 11996
rect 5386 11940 5390 11996
rect 5326 11936 5390 11940
rect 5406 11996 5470 12000
rect 5406 11940 5410 11996
rect 5410 11940 5466 11996
rect 5466 11940 5470 11996
rect 5406 11936 5470 11940
rect 5486 11996 5550 12000
rect 5486 11940 5490 11996
rect 5490 11940 5546 11996
rect 5546 11940 5550 11996
rect 5486 11936 5550 11940
rect 5566 11996 5630 12000
rect 5566 11940 5570 11996
rect 5570 11940 5626 11996
rect 5626 11940 5630 11996
rect 5566 11936 5630 11940
rect 12754 11996 12818 12000
rect 12754 11940 12758 11996
rect 12758 11940 12814 11996
rect 12814 11940 12818 11996
rect 12754 11936 12818 11940
rect 12834 11996 12898 12000
rect 12834 11940 12838 11996
rect 12838 11940 12894 11996
rect 12894 11940 12898 11996
rect 12834 11936 12898 11940
rect 12914 11996 12978 12000
rect 12914 11940 12918 11996
rect 12918 11940 12974 11996
rect 12974 11940 12978 11996
rect 12914 11936 12978 11940
rect 12994 11996 13058 12000
rect 12994 11940 12998 11996
rect 12998 11940 13054 11996
rect 13054 11940 13058 11996
rect 12994 11936 13058 11940
rect 20182 11996 20246 12000
rect 20182 11940 20186 11996
rect 20186 11940 20242 11996
rect 20242 11940 20246 11996
rect 20182 11936 20246 11940
rect 20262 11996 20326 12000
rect 20262 11940 20266 11996
rect 20266 11940 20322 11996
rect 20322 11940 20326 11996
rect 20262 11936 20326 11940
rect 20342 11996 20406 12000
rect 20342 11940 20346 11996
rect 20346 11940 20402 11996
rect 20402 11940 20406 11996
rect 20342 11936 20406 11940
rect 20422 11996 20486 12000
rect 20422 11940 20426 11996
rect 20426 11940 20482 11996
rect 20482 11940 20486 11996
rect 20422 11936 20486 11940
rect 27610 11996 27674 12000
rect 27610 11940 27614 11996
rect 27614 11940 27670 11996
rect 27670 11940 27674 11996
rect 27610 11936 27674 11940
rect 27690 11996 27754 12000
rect 27690 11940 27694 11996
rect 27694 11940 27750 11996
rect 27750 11940 27754 11996
rect 27690 11936 27754 11940
rect 27770 11996 27834 12000
rect 27770 11940 27774 11996
rect 27774 11940 27830 11996
rect 27830 11940 27834 11996
rect 27770 11936 27834 11940
rect 27850 11996 27914 12000
rect 27850 11940 27854 11996
rect 27854 11940 27910 11996
rect 27910 11940 27914 11996
rect 27850 11936 27914 11940
rect 4666 11452 4730 11456
rect 4666 11396 4670 11452
rect 4670 11396 4726 11452
rect 4726 11396 4730 11452
rect 4666 11392 4730 11396
rect 4746 11452 4810 11456
rect 4746 11396 4750 11452
rect 4750 11396 4806 11452
rect 4806 11396 4810 11452
rect 4746 11392 4810 11396
rect 4826 11452 4890 11456
rect 4826 11396 4830 11452
rect 4830 11396 4886 11452
rect 4886 11396 4890 11452
rect 4826 11392 4890 11396
rect 4906 11452 4970 11456
rect 4906 11396 4910 11452
rect 4910 11396 4966 11452
rect 4966 11396 4970 11452
rect 4906 11392 4970 11396
rect 12094 11452 12158 11456
rect 12094 11396 12098 11452
rect 12098 11396 12154 11452
rect 12154 11396 12158 11452
rect 12094 11392 12158 11396
rect 12174 11452 12238 11456
rect 12174 11396 12178 11452
rect 12178 11396 12234 11452
rect 12234 11396 12238 11452
rect 12174 11392 12238 11396
rect 12254 11452 12318 11456
rect 12254 11396 12258 11452
rect 12258 11396 12314 11452
rect 12314 11396 12318 11452
rect 12254 11392 12318 11396
rect 12334 11452 12398 11456
rect 12334 11396 12338 11452
rect 12338 11396 12394 11452
rect 12394 11396 12398 11452
rect 12334 11392 12398 11396
rect 19522 11452 19586 11456
rect 19522 11396 19526 11452
rect 19526 11396 19582 11452
rect 19582 11396 19586 11452
rect 19522 11392 19586 11396
rect 19602 11452 19666 11456
rect 19602 11396 19606 11452
rect 19606 11396 19662 11452
rect 19662 11396 19666 11452
rect 19602 11392 19666 11396
rect 19682 11452 19746 11456
rect 19682 11396 19686 11452
rect 19686 11396 19742 11452
rect 19742 11396 19746 11452
rect 19682 11392 19746 11396
rect 19762 11452 19826 11456
rect 19762 11396 19766 11452
rect 19766 11396 19822 11452
rect 19822 11396 19826 11452
rect 19762 11392 19826 11396
rect 26950 11452 27014 11456
rect 26950 11396 26954 11452
rect 26954 11396 27010 11452
rect 27010 11396 27014 11452
rect 26950 11392 27014 11396
rect 27030 11452 27094 11456
rect 27030 11396 27034 11452
rect 27034 11396 27090 11452
rect 27090 11396 27094 11452
rect 27030 11392 27094 11396
rect 27110 11452 27174 11456
rect 27110 11396 27114 11452
rect 27114 11396 27170 11452
rect 27170 11396 27174 11452
rect 27110 11392 27174 11396
rect 27190 11452 27254 11456
rect 27190 11396 27194 11452
rect 27194 11396 27250 11452
rect 27250 11396 27254 11452
rect 27190 11392 27254 11396
rect 5326 10908 5390 10912
rect 5326 10852 5330 10908
rect 5330 10852 5386 10908
rect 5386 10852 5390 10908
rect 5326 10848 5390 10852
rect 5406 10908 5470 10912
rect 5406 10852 5410 10908
rect 5410 10852 5466 10908
rect 5466 10852 5470 10908
rect 5406 10848 5470 10852
rect 5486 10908 5550 10912
rect 5486 10852 5490 10908
rect 5490 10852 5546 10908
rect 5546 10852 5550 10908
rect 5486 10848 5550 10852
rect 5566 10908 5630 10912
rect 5566 10852 5570 10908
rect 5570 10852 5626 10908
rect 5626 10852 5630 10908
rect 5566 10848 5630 10852
rect 12754 10908 12818 10912
rect 12754 10852 12758 10908
rect 12758 10852 12814 10908
rect 12814 10852 12818 10908
rect 12754 10848 12818 10852
rect 12834 10908 12898 10912
rect 12834 10852 12838 10908
rect 12838 10852 12894 10908
rect 12894 10852 12898 10908
rect 12834 10848 12898 10852
rect 12914 10908 12978 10912
rect 12914 10852 12918 10908
rect 12918 10852 12974 10908
rect 12974 10852 12978 10908
rect 12914 10848 12978 10852
rect 12994 10908 13058 10912
rect 12994 10852 12998 10908
rect 12998 10852 13054 10908
rect 13054 10852 13058 10908
rect 12994 10848 13058 10852
rect 20182 10908 20246 10912
rect 20182 10852 20186 10908
rect 20186 10852 20242 10908
rect 20242 10852 20246 10908
rect 20182 10848 20246 10852
rect 20262 10908 20326 10912
rect 20262 10852 20266 10908
rect 20266 10852 20322 10908
rect 20322 10852 20326 10908
rect 20262 10848 20326 10852
rect 20342 10908 20406 10912
rect 20342 10852 20346 10908
rect 20346 10852 20402 10908
rect 20402 10852 20406 10908
rect 20342 10848 20406 10852
rect 20422 10908 20486 10912
rect 20422 10852 20426 10908
rect 20426 10852 20482 10908
rect 20482 10852 20486 10908
rect 20422 10848 20486 10852
rect 27610 10908 27674 10912
rect 27610 10852 27614 10908
rect 27614 10852 27670 10908
rect 27670 10852 27674 10908
rect 27610 10848 27674 10852
rect 27690 10908 27754 10912
rect 27690 10852 27694 10908
rect 27694 10852 27750 10908
rect 27750 10852 27754 10908
rect 27690 10848 27754 10852
rect 27770 10908 27834 10912
rect 27770 10852 27774 10908
rect 27774 10852 27830 10908
rect 27830 10852 27834 10908
rect 27770 10848 27834 10852
rect 27850 10908 27914 10912
rect 27850 10852 27854 10908
rect 27854 10852 27910 10908
rect 27910 10852 27914 10908
rect 27850 10848 27914 10852
rect 4666 10364 4730 10368
rect 4666 10308 4670 10364
rect 4670 10308 4726 10364
rect 4726 10308 4730 10364
rect 4666 10304 4730 10308
rect 4746 10364 4810 10368
rect 4746 10308 4750 10364
rect 4750 10308 4806 10364
rect 4806 10308 4810 10364
rect 4746 10304 4810 10308
rect 4826 10364 4890 10368
rect 4826 10308 4830 10364
rect 4830 10308 4886 10364
rect 4886 10308 4890 10364
rect 4826 10304 4890 10308
rect 4906 10364 4970 10368
rect 4906 10308 4910 10364
rect 4910 10308 4966 10364
rect 4966 10308 4970 10364
rect 4906 10304 4970 10308
rect 12094 10364 12158 10368
rect 12094 10308 12098 10364
rect 12098 10308 12154 10364
rect 12154 10308 12158 10364
rect 12094 10304 12158 10308
rect 12174 10364 12238 10368
rect 12174 10308 12178 10364
rect 12178 10308 12234 10364
rect 12234 10308 12238 10364
rect 12174 10304 12238 10308
rect 12254 10364 12318 10368
rect 12254 10308 12258 10364
rect 12258 10308 12314 10364
rect 12314 10308 12318 10364
rect 12254 10304 12318 10308
rect 12334 10364 12398 10368
rect 12334 10308 12338 10364
rect 12338 10308 12394 10364
rect 12394 10308 12398 10364
rect 12334 10304 12398 10308
rect 19522 10364 19586 10368
rect 19522 10308 19526 10364
rect 19526 10308 19582 10364
rect 19582 10308 19586 10364
rect 19522 10304 19586 10308
rect 19602 10364 19666 10368
rect 19602 10308 19606 10364
rect 19606 10308 19662 10364
rect 19662 10308 19666 10364
rect 19602 10304 19666 10308
rect 19682 10364 19746 10368
rect 19682 10308 19686 10364
rect 19686 10308 19742 10364
rect 19742 10308 19746 10364
rect 19682 10304 19746 10308
rect 19762 10364 19826 10368
rect 19762 10308 19766 10364
rect 19766 10308 19822 10364
rect 19822 10308 19826 10364
rect 19762 10304 19826 10308
rect 26950 10364 27014 10368
rect 26950 10308 26954 10364
rect 26954 10308 27010 10364
rect 27010 10308 27014 10364
rect 26950 10304 27014 10308
rect 27030 10364 27094 10368
rect 27030 10308 27034 10364
rect 27034 10308 27090 10364
rect 27090 10308 27094 10364
rect 27030 10304 27094 10308
rect 27110 10364 27174 10368
rect 27110 10308 27114 10364
rect 27114 10308 27170 10364
rect 27170 10308 27174 10364
rect 27110 10304 27174 10308
rect 27190 10364 27254 10368
rect 27190 10308 27194 10364
rect 27194 10308 27250 10364
rect 27250 10308 27254 10364
rect 27190 10304 27254 10308
rect 5326 9820 5390 9824
rect 5326 9764 5330 9820
rect 5330 9764 5386 9820
rect 5386 9764 5390 9820
rect 5326 9760 5390 9764
rect 5406 9820 5470 9824
rect 5406 9764 5410 9820
rect 5410 9764 5466 9820
rect 5466 9764 5470 9820
rect 5406 9760 5470 9764
rect 5486 9820 5550 9824
rect 5486 9764 5490 9820
rect 5490 9764 5546 9820
rect 5546 9764 5550 9820
rect 5486 9760 5550 9764
rect 5566 9820 5630 9824
rect 5566 9764 5570 9820
rect 5570 9764 5626 9820
rect 5626 9764 5630 9820
rect 5566 9760 5630 9764
rect 12754 9820 12818 9824
rect 12754 9764 12758 9820
rect 12758 9764 12814 9820
rect 12814 9764 12818 9820
rect 12754 9760 12818 9764
rect 12834 9820 12898 9824
rect 12834 9764 12838 9820
rect 12838 9764 12894 9820
rect 12894 9764 12898 9820
rect 12834 9760 12898 9764
rect 12914 9820 12978 9824
rect 12914 9764 12918 9820
rect 12918 9764 12974 9820
rect 12974 9764 12978 9820
rect 12914 9760 12978 9764
rect 12994 9820 13058 9824
rect 12994 9764 12998 9820
rect 12998 9764 13054 9820
rect 13054 9764 13058 9820
rect 12994 9760 13058 9764
rect 20182 9820 20246 9824
rect 20182 9764 20186 9820
rect 20186 9764 20242 9820
rect 20242 9764 20246 9820
rect 20182 9760 20246 9764
rect 20262 9820 20326 9824
rect 20262 9764 20266 9820
rect 20266 9764 20322 9820
rect 20322 9764 20326 9820
rect 20262 9760 20326 9764
rect 20342 9820 20406 9824
rect 20342 9764 20346 9820
rect 20346 9764 20402 9820
rect 20402 9764 20406 9820
rect 20342 9760 20406 9764
rect 20422 9820 20486 9824
rect 20422 9764 20426 9820
rect 20426 9764 20482 9820
rect 20482 9764 20486 9820
rect 20422 9760 20486 9764
rect 27610 9820 27674 9824
rect 27610 9764 27614 9820
rect 27614 9764 27670 9820
rect 27670 9764 27674 9820
rect 27610 9760 27674 9764
rect 27690 9820 27754 9824
rect 27690 9764 27694 9820
rect 27694 9764 27750 9820
rect 27750 9764 27754 9820
rect 27690 9760 27754 9764
rect 27770 9820 27834 9824
rect 27770 9764 27774 9820
rect 27774 9764 27830 9820
rect 27830 9764 27834 9820
rect 27770 9760 27834 9764
rect 27850 9820 27914 9824
rect 27850 9764 27854 9820
rect 27854 9764 27910 9820
rect 27910 9764 27914 9820
rect 27850 9760 27914 9764
rect 4666 9276 4730 9280
rect 4666 9220 4670 9276
rect 4670 9220 4726 9276
rect 4726 9220 4730 9276
rect 4666 9216 4730 9220
rect 4746 9276 4810 9280
rect 4746 9220 4750 9276
rect 4750 9220 4806 9276
rect 4806 9220 4810 9276
rect 4746 9216 4810 9220
rect 4826 9276 4890 9280
rect 4826 9220 4830 9276
rect 4830 9220 4886 9276
rect 4886 9220 4890 9276
rect 4826 9216 4890 9220
rect 4906 9276 4970 9280
rect 4906 9220 4910 9276
rect 4910 9220 4966 9276
rect 4966 9220 4970 9276
rect 4906 9216 4970 9220
rect 12094 9276 12158 9280
rect 12094 9220 12098 9276
rect 12098 9220 12154 9276
rect 12154 9220 12158 9276
rect 12094 9216 12158 9220
rect 12174 9276 12238 9280
rect 12174 9220 12178 9276
rect 12178 9220 12234 9276
rect 12234 9220 12238 9276
rect 12174 9216 12238 9220
rect 12254 9276 12318 9280
rect 12254 9220 12258 9276
rect 12258 9220 12314 9276
rect 12314 9220 12318 9276
rect 12254 9216 12318 9220
rect 12334 9276 12398 9280
rect 12334 9220 12338 9276
rect 12338 9220 12394 9276
rect 12394 9220 12398 9276
rect 12334 9216 12398 9220
rect 19522 9276 19586 9280
rect 19522 9220 19526 9276
rect 19526 9220 19582 9276
rect 19582 9220 19586 9276
rect 19522 9216 19586 9220
rect 19602 9276 19666 9280
rect 19602 9220 19606 9276
rect 19606 9220 19662 9276
rect 19662 9220 19666 9276
rect 19602 9216 19666 9220
rect 19682 9276 19746 9280
rect 19682 9220 19686 9276
rect 19686 9220 19742 9276
rect 19742 9220 19746 9276
rect 19682 9216 19746 9220
rect 19762 9276 19826 9280
rect 19762 9220 19766 9276
rect 19766 9220 19822 9276
rect 19822 9220 19826 9276
rect 19762 9216 19826 9220
rect 26950 9276 27014 9280
rect 26950 9220 26954 9276
rect 26954 9220 27010 9276
rect 27010 9220 27014 9276
rect 26950 9216 27014 9220
rect 27030 9276 27094 9280
rect 27030 9220 27034 9276
rect 27034 9220 27090 9276
rect 27090 9220 27094 9276
rect 27030 9216 27094 9220
rect 27110 9276 27174 9280
rect 27110 9220 27114 9276
rect 27114 9220 27170 9276
rect 27170 9220 27174 9276
rect 27110 9216 27174 9220
rect 27190 9276 27254 9280
rect 27190 9220 27194 9276
rect 27194 9220 27250 9276
rect 27250 9220 27254 9276
rect 27190 9216 27254 9220
rect 5326 8732 5390 8736
rect 5326 8676 5330 8732
rect 5330 8676 5386 8732
rect 5386 8676 5390 8732
rect 5326 8672 5390 8676
rect 5406 8732 5470 8736
rect 5406 8676 5410 8732
rect 5410 8676 5466 8732
rect 5466 8676 5470 8732
rect 5406 8672 5470 8676
rect 5486 8732 5550 8736
rect 5486 8676 5490 8732
rect 5490 8676 5546 8732
rect 5546 8676 5550 8732
rect 5486 8672 5550 8676
rect 5566 8732 5630 8736
rect 5566 8676 5570 8732
rect 5570 8676 5626 8732
rect 5626 8676 5630 8732
rect 5566 8672 5630 8676
rect 12754 8732 12818 8736
rect 12754 8676 12758 8732
rect 12758 8676 12814 8732
rect 12814 8676 12818 8732
rect 12754 8672 12818 8676
rect 12834 8732 12898 8736
rect 12834 8676 12838 8732
rect 12838 8676 12894 8732
rect 12894 8676 12898 8732
rect 12834 8672 12898 8676
rect 12914 8732 12978 8736
rect 12914 8676 12918 8732
rect 12918 8676 12974 8732
rect 12974 8676 12978 8732
rect 12914 8672 12978 8676
rect 12994 8732 13058 8736
rect 12994 8676 12998 8732
rect 12998 8676 13054 8732
rect 13054 8676 13058 8732
rect 12994 8672 13058 8676
rect 20182 8732 20246 8736
rect 20182 8676 20186 8732
rect 20186 8676 20242 8732
rect 20242 8676 20246 8732
rect 20182 8672 20246 8676
rect 20262 8732 20326 8736
rect 20262 8676 20266 8732
rect 20266 8676 20322 8732
rect 20322 8676 20326 8732
rect 20262 8672 20326 8676
rect 20342 8732 20406 8736
rect 20342 8676 20346 8732
rect 20346 8676 20402 8732
rect 20402 8676 20406 8732
rect 20342 8672 20406 8676
rect 20422 8732 20486 8736
rect 20422 8676 20426 8732
rect 20426 8676 20482 8732
rect 20482 8676 20486 8732
rect 20422 8672 20486 8676
rect 27610 8732 27674 8736
rect 27610 8676 27614 8732
rect 27614 8676 27670 8732
rect 27670 8676 27674 8732
rect 27610 8672 27674 8676
rect 27690 8732 27754 8736
rect 27690 8676 27694 8732
rect 27694 8676 27750 8732
rect 27750 8676 27754 8732
rect 27690 8672 27754 8676
rect 27770 8732 27834 8736
rect 27770 8676 27774 8732
rect 27774 8676 27830 8732
rect 27830 8676 27834 8732
rect 27770 8672 27834 8676
rect 27850 8732 27914 8736
rect 27850 8676 27854 8732
rect 27854 8676 27910 8732
rect 27910 8676 27914 8732
rect 27850 8672 27914 8676
rect 4666 8188 4730 8192
rect 4666 8132 4670 8188
rect 4670 8132 4726 8188
rect 4726 8132 4730 8188
rect 4666 8128 4730 8132
rect 4746 8188 4810 8192
rect 4746 8132 4750 8188
rect 4750 8132 4806 8188
rect 4806 8132 4810 8188
rect 4746 8128 4810 8132
rect 4826 8188 4890 8192
rect 4826 8132 4830 8188
rect 4830 8132 4886 8188
rect 4886 8132 4890 8188
rect 4826 8128 4890 8132
rect 4906 8188 4970 8192
rect 4906 8132 4910 8188
rect 4910 8132 4966 8188
rect 4966 8132 4970 8188
rect 4906 8128 4970 8132
rect 12094 8188 12158 8192
rect 12094 8132 12098 8188
rect 12098 8132 12154 8188
rect 12154 8132 12158 8188
rect 12094 8128 12158 8132
rect 12174 8188 12238 8192
rect 12174 8132 12178 8188
rect 12178 8132 12234 8188
rect 12234 8132 12238 8188
rect 12174 8128 12238 8132
rect 12254 8188 12318 8192
rect 12254 8132 12258 8188
rect 12258 8132 12314 8188
rect 12314 8132 12318 8188
rect 12254 8128 12318 8132
rect 12334 8188 12398 8192
rect 12334 8132 12338 8188
rect 12338 8132 12394 8188
rect 12394 8132 12398 8188
rect 12334 8128 12398 8132
rect 19522 8188 19586 8192
rect 19522 8132 19526 8188
rect 19526 8132 19582 8188
rect 19582 8132 19586 8188
rect 19522 8128 19586 8132
rect 19602 8188 19666 8192
rect 19602 8132 19606 8188
rect 19606 8132 19662 8188
rect 19662 8132 19666 8188
rect 19602 8128 19666 8132
rect 19682 8188 19746 8192
rect 19682 8132 19686 8188
rect 19686 8132 19742 8188
rect 19742 8132 19746 8188
rect 19682 8128 19746 8132
rect 19762 8188 19826 8192
rect 19762 8132 19766 8188
rect 19766 8132 19822 8188
rect 19822 8132 19826 8188
rect 19762 8128 19826 8132
rect 26950 8188 27014 8192
rect 26950 8132 26954 8188
rect 26954 8132 27010 8188
rect 27010 8132 27014 8188
rect 26950 8128 27014 8132
rect 27030 8188 27094 8192
rect 27030 8132 27034 8188
rect 27034 8132 27090 8188
rect 27090 8132 27094 8188
rect 27030 8128 27094 8132
rect 27110 8188 27174 8192
rect 27110 8132 27114 8188
rect 27114 8132 27170 8188
rect 27170 8132 27174 8188
rect 27110 8128 27174 8132
rect 27190 8188 27254 8192
rect 27190 8132 27194 8188
rect 27194 8132 27250 8188
rect 27250 8132 27254 8188
rect 27190 8128 27254 8132
rect 5326 7644 5390 7648
rect 5326 7588 5330 7644
rect 5330 7588 5386 7644
rect 5386 7588 5390 7644
rect 5326 7584 5390 7588
rect 5406 7644 5470 7648
rect 5406 7588 5410 7644
rect 5410 7588 5466 7644
rect 5466 7588 5470 7644
rect 5406 7584 5470 7588
rect 5486 7644 5550 7648
rect 5486 7588 5490 7644
rect 5490 7588 5546 7644
rect 5546 7588 5550 7644
rect 5486 7584 5550 7588
rect 5566 7644 5630 7648
rect 5566 7588 5570 7644
rect 5570 7588 5626 7644
rect 5626 7588 5630 7644
rect 5566 7584 5630 7588
rect 12754 7644 12818 7648
rect 12754 7588 12758 7644
rect 12758 7588 12814 7644
rect 12814 7588 12818 7644
rect 12754 7584 12818 7588
rect 12834 7644 12898 7648
rect 12834 7588 12838 7644
rect 12838 7588 12894 7644
rect 12894 7588 12898 7644
rect 12834 7584 12898 7588
rect 12914 7644 12978 7648
rect 12914 7588 12918 7644
rect 12918 7588 12974 7644
rect 12974 7588 12978 7644
rect 12914 7584 12978 7588
rect 12994 7644 13058 7648
rect 12994 7588 12998 7644
rect 12998 7588 13054 7644
rect 13054 7588 13058 7644
rect 12994 7584 13058 7588
rect 20182 7644 20246 7648
rect 20182 7588 20186 7644
rect 20186 7588 20242 7644
rect 20242 7588 20246 7644
rect 20182 7584 20246 7588
rect 20262 7644 20326 7648
rect 20262 7588 20266 7644
rect 20266 7588 20322 7644
rect 20322 7588 20326 7644
rect 20262 7584 20326 7588
rect 20342 7644 20406 7648
rect 20342 7588 20346 7644
rect 20346 7588 20402 7644
rect 20402 7588 20406 7644
rect 20342 7584 20406 7588
rect 20422 7644 20486 7648
rect 20422 7588 20426 7644
rect 20426 7588 20482 7644
rect 20482 7588 20486 7644
rect 20422 7584 20486 7588
rect 27610 7644 27674 7648
rect 27610 7588 27614 7644
rect 27614 7588 27670 7644
rect 27670 7588 27674 7644
rect 27610 7584 27674 7588
rect 27690 7644 27754 7648
rect 27690 7588 27694 7644
rect 27694 7588 27750 7644
rect 27750 7588 27754 7644
rect 27690 7584 27754 7588
rect 27770 7644 27834 7648
rect 27770 7588 27774 7644
rect 27774 7588 27830 7644
rect 27830 7588 27834 7644
rect 27770 7584 27834 7588
rect 27850 7644 27914 7648
rect 27850 7588 27854 7644
rect 27854 7588 27910 7644
rect 27910 7588 27914 7644
rect 27850 7584 27914 7588
rect 4666 7100 4730 7104
rect 4666 7044 4670 7100
rect 4670 7044 4726 7100
rect 4726 7044 4730 7100
rect 4666 7040 4730 7044
rect 4746 7100 4810 7104
rect 4746 7044 4750 7100
rect 4750 7044 4806 7100
rect 4806 7044 4810 7100
rect 4746 7040 4810 7044
rect 4826 7100 4890 7104
rect 4826 7044 4830 7100
rect 4830 7044 4886 7100
rect 4886 7044 4890 7100
rect 4826 7040 4890 7044
rect 4906 7100 4970 7104
rect 4906 7044 4910 7100
rect 4910 7044 4966 7100
rect 4966 7044 4970 7100
rect 4906 7040 4970 7044
rect 12094 7100 12158 7104
rect 12094 7044 12098 7100
rect 12098 7044 12154 7100
rect 12154 7044 12158 7100
rect 12094 7040 12158 7044
rect 12174 7100 12238 7104
rect 12174 7044 12178 7100
rect 12178 7044 12234 7100
rect 12234 7044 12238 7100
rect 12174 7040 12238 7044
rect 12254 7100 12318 7104
rect 12254 7044 12258 7100
rect 12258 7044 12314 7100
rect 12314 7044 12318 7100
rect 12254 7040 12318 7044
rect 12334 7100 12398 7104
rect 12334 7044 12338 7100
rect 12338 7044 12394 7100
rect 12394 7044 12398 7100
rect 12334 7040 12398 7044
rect 19522 7100 19586 7104
rect 19522 7044 19526 7100
rect 19526 7044 19582 7100
rect 19582 7044 19586 7100
rect 19522 7040 19586 7044
rect 19602 7100 19666 7104
rect 19602 7044 19606 7100
rect 19606 7044 19662 7100
rect 19662 7044 19666 7100
rect 19602 7040 19666 7044
rect 19682 7100 19746 7104
rect 19682 7044 19686 7100
rect 19686 7044 19742 7100
rect 19742 7044 19746 7100
rect 19682 7040 19746 7044
rect 19762 7100 19826 7104
rect 19762 7044 19766 7100
rect 19766 7044 19822 7100
rect 19822 7044 19826 7100
rect 19762 7040 19826 7044
rect 26950 7100 27014 7104
rect 26950 7044 26954 7100
rect 26954 7044 27010 7100
rect 27010 7044 27014 7100
rect 26950 7040 27014 7044
rect 27030 7100 27094 7104
rect 27030 7044 27034 7100
rect 27034 7044 27090 7100
rect 27090 7044 27094 7100
rect 27030 7040 27094 7044
rect 27110 7100 27174 7104
rect 27110 7044 27114 7100
rect 27114 7044 27170 7100
rect 27170 7044 27174 7100
rect 27110 7040 27174 7044
rect 27190 7100 27254 7104
rect 27190 7044 27194 7100
rect 27194 7044 27250 7100
rect 27250 7044 27254 7100
rect 27190 7040 27254 7044
rect 5326 6556 5390 6560
rect 5326 6500 5330 6556
rect 5330 6500 5386 6556
rect 5386 6500 5390 6556
rect 5326 6496 5390 6500
rect 5406 6556 5470 6560
rect 5406 6500 5410 6556
rect 5410 6500 5466 6556
rect 5466 6500 5470 6556
rect 5406 6496 5470 6500
rect 5486 6556 5550 6560
rect 5486 6500 5490 6556
rect 5490 6500 5546 6556
rect 5546 6500 5550 6556
rect 5486 6496 5550 6500
rect 5566 6556 5630 6560
rect 5566 6500 5570 6556
rect 5570 6500 5626 6556
rect 5626 6500 5630 6556
rect 5566 6496 5630 6500
rect 12754 6556 12818 6560
rect 12754 6500 12758 6556
rect 12758 6500 12814 6556
rect 12814 6500 12818 6556
rect 12754 6496 12818 6500
rect 12834 6556 12898 6560
rect 12834 6500 12838 6556
rect 12838 6500 12894 6556
rect 12894 6500 12898 6556
rect 12834 6496 12898 6500
rect 12914 6556 12978 6560
rect 12914 6500 12918 6556
rect 12918 6500 12974 6556
rect 12974 6500 12978 6556
rect 12914 6496 12978 6500
rect 12994 6556 13058 6560
rect 12994 6500 12998 6556
rect 12998 6500 13054 6556
rect 13054 6500 13058 6556
rect 12994 6496 13058 6500
rect 20182 6556 20246 6560
rect 20182 6500 20186 6556
rect 20186 6500 20242 6556
rect 20242 6500 20246 6556
rect 20182 6496 20246 6500
rect 20262 6556 20326 6560
rect 20262 6500 20266 6556
rect 20266 6500 20322 6556
rect 20322 6500 20326 6556
rect 20262 6496 20326 6500
rect 20342 6556 20406 6560
rect 20342 6500 20346 6556
rect 20346 6500 20402 6556
rect 20402 6500 20406 6556
rect 20342 6496 20406 6500
rect 20422 6556 20486 6560
rect 20422 6500 20426 6556
rect 20426 6500 20482 6556
rect 20482 6500 20486 6556
rect 20422 6496 20486 6500
rect 27610 6556 27674 6560
rect 27610 6500 27614 6556
rect 27614 6500 27670 6556
rect 27670 6500 27674 6556
rect 27610 6496 27674 6500
rect 27690 6556 27754 6560
rect 27690 6500 27694 6556
rect 27694 6500 27750 6556
rect 27750 6500 27754 6556
rect 27690 6496 27754 6500
rect 27770 6556 27834 6560
rect 27770 6500 27774 6556
rect 27774 6500 27830 6556
rect 27830 6500 27834 6556
rect 27770 6496 27834 6500
rect 27850 6556 27914 6560
rect 27850 6500 27854 6556
rect 27854 6500 27910 6556
rect 27910 6500 27914 6556
rect 27850 6496 27914 6500
rect 4666 6012 4730 6016
rect 4666 5956 4670 6012
rect 4670 5956 4726 6012
rect 4726 5956 4730 6012
rect 4666 5952 4730 5956
rect 4746 6012 4810 6016
rect 4746 5956 4750 6012
rect 4750 5956 4806 6012
rect 4806 5956 4810 6012
rect 4746 5952 4810 5956
rect 4826 6012 4890 6016
rect 4826 5956 4830 6012
rect 4830 5956 4886 6012
rect 4886 5956 4890 6012
rect 4826 5952 4890 5956
rect 4906 6012 4970 6016
rect 4906 5956 4910 6012
rect 4910 5956 4966 6012
rect 4966 5956 4970 6012
rect 4906 5952 4970 5956
rect 12094 6012 12158 6016
rect 12094 5956 12098 6012
rect 12098 5956 12154 6012
rect 12154 5956 12158 6012
rect 12094 5952 12158 5956
rect 12174 6012 12238 6016
rect 12174 5956 12178 6012
rect 12178 5956 12234 6012
rect 12234 5956 12238 6012
rect 12174 5952 12238 5956
rect 12254 6012 12318 6016
rect 12254 5956 12258 6012
rect 12258 5956 12314 6012
rect 12314 5956 12318 6012
rect 12254 5952 12318 5956
rect 12334 6012 12398 6016
rect 12334 5956 12338 6012
rect 12338 5956 12394 6012
rect 12394 5956 12398 6012
rect 12334 5952 12398 5956
rect 19522 6012 19586 6016
rect 19522 5956 19526 6012
rect 19526 5956 19582 6012
rect 19582 5956 19586 6012
rect 19522 5952 19586 5956
rect 19602 6012 19666 6016
rect 19602 5956 19606 6012
rect 19606 5956 19662 6012
rect 19662 5956 19666 6012
rect 19602 5952 19666 5956
rect 19682 6012 19746 6016
rect 19682 5956 19686 6012
rect 19686 5956 19742 6012
rect 19742 5956 19746 6012
rect 19682 5952 19746 5956
rect 19762 6012 19826 6016
rect 19762 5956 19766 6012
rect 19766 5956 19822 6012
rect 19822 5956 19826 6012
rect 19762 5952 19826 5956
rect 26950 6012 27014 6016
rect 26950 5956 26954 6012
rect 26954 5956 27010 6012
rect 27010 5956 27014 6012
rect 26950 5952 27014 5956
rect 27030 6012 27094 6016
rect 27030 5956 27034 6012
rect 27034 5956 27090 6012
rect 27090 5956 27094 6012
rect 27030 5952 27094 5956
rect 27110 6012 27174 6016
rect 27110 5956 27114 6012
rect 27114 5956 27170 6012
rect 27170 5956 27174 6012
rect 27110 5952 27174 5956
rect 27190 6012 27254 6016
rect 27190 5956 27194 6012
rect 27194 5956 27250 6012
rect 27250 5956 27254 6012
rect 27190 5952 27254 5956
rect 5326 5468 5390 5472
rect 5326 5412 5330 5468
rect 5330 5412 5386 5468
rect 5386 5412 5390 5468
rect 5326 5408 5390 5412
rect 5406 5468 5470 5472
rect 5406 5412 5410 5468
rect 5410 5412 5466 5468
rect 5466 5412 5470 5468
rect 5406 5408 5470 5412
rect 5486 5468 5550 5472
rect 5486 5412 5490 5468
rect 5490 5412 5546 5468
rect 5546 5412 5550 5468
rect 5486 5408 5550 5412
rect 5566 5468 5630 5472
rect 5566 5412 5570 5468
rect 5570 5412 5626 5468
rect 5626 5412 5630 5468
rect 5566 5408 5630 5412
rect 12754 5468 12818 5472
rect 12754 5412 12758 5468
rect 12758 5412 12814 5468
rect 12814 5412 12818 5468
rect 12754 5408 12818 5412
rect 12834 5468 12898 5472
rect 12834 5412 12838 5468
rect 12838 5412 12894 5468
rect 12894 5412 12898 5468
rect 12834 5408 12898 5412
rect 12914 5468 12978 5472
rect 12914 5412 12918 5468
rect 12918 5412 12974 5468
rect 12974 5412 12978 5468
rect 12914 5408 12978 5412
rect 12994 5468 13058 5472
rect 12994 5412 12998 5468
rect 12998 5412 13054 5468
rect 13054 5412 13058 5468
rect 12994 5408 13058 5412
rect 20182 5468 20246 5472
rect 20182 5412 20186 5468
rect 20186 5412 20242 5468
rect 20242 5412 20246 5468
rect 20182 5408 20246 5412
rect 20262 5468 20326 5472
rect 20262 5412 20266 5468
rect 20266 5412 20322 5468
rect 20322 5412 20326 5468
rect 20262 5408 20326 5412
rect 20342 5468 20406 5472
rect 20342 5412 20346 5468
rect 20346 5412 20402 5468
rect 20402 5412 20406 5468
rect 20342 5408 20406 5412
rect 20422 5468 20486 5472
rect 20422 5412 20426 5468
rect 20426 5412 20482 5468
rect 20482 5412 20486 5468
rect 20422 5408 20486 5412
rect 27610 5468 27674 5472
rect 27610 5412 27614 5468
rect 27614 5412 27670 5468
rect 27670 5412 27674 5468
rect 27610 5408 27674 5412
rect 27690 5468 27754 5472
rect 27690 5412 27694 5468
rect 27694 5412 27750 5468
rect 27750 5412 27754 5468
rect 27690 5408 27754 5412
rect 27770 5468 27834 5472
rect 27770 5412 27774 5468
rect 27774 5412 27830 5468
rect 27830 5412 27834 5468
rect 27770 5408 27834 5412
rect 27850 5468 27914 5472
rect 27850 5412 27854 5468
rect 27854 5412 27910 5468
rect 27910 5412 27914 5468
rect 27850 5408 27914 5412
rect 4666 4924 4730 4928
rect 4666 4868 4670 4924
rect 4670 4868 4726 4924
rect 4726 4868 4730 4924
rect 4666 4864 4730 4868
rect 4746 4924 4810 4928
rect 4746 4868 4750 4924
rect 4750 4868 4806 4924
rect 4806 4868 4810 4924
rect 4746 4864 4810 4868
rect 4826 4924 4890 4928
rect 4826 4868 4830 4924
rect 4830 4868 4886 4924
rect 4886 4868 4890 4924
rect 4826 4864 4890 4868
rect 4906 4924 4970 4928
rect 4906 4868 4910 4924
rect 4910 4868 4966 4924
rect 4966 4868 4970 4924
rect 4906 4864 4970 4868
rect 12094 4924 12158 4928
rect 12094 4868 12098 4924
rect 12098 4868 12154 4924
rect 12154 4868 12158 4924
rect 12094 4864 12158 4868
rect 12174 4924 12238 4928
rect 12174 4868 12178 4924
rect 12178 4868 12234 4924
rect 12234 4868 12238 4924
rect 12174 4864 12238 4868
rect 12254 4924 12318 4928
rect 12254 4868 12258 4924
rect 12258 4868 12314 4924
rect 12314 4868 12318 4924
rect 12254 4864 12318 4868
rect 12334 4924 12398 4928
rect 12334 4868 12338 4924
rect 12338 4868 12394 4924
rect 12394 4868 12398 4924
rect 12334 4864 12398 4868
rect 19522 4924 19586 4928
rect 19522 4868 19526 4924
rect 19526 4868 19582 4924
rect 19582 4868 19586 4924
rect 19522 4864 19586 4868
rect 19602 4924 19666 4928
rect 19602 4868 19606 4924
rect 19606 4868 19662 4924
rect 19662 4868 19666 4924
rect 19602 4864 19666 4868
rect 19682 4924 19746 4928
rect 19682 4868 19686 4924
rect 19686 4868 19742 4924
rect 19742 4868 19746 4924
rect 19682 4864 19746 4868
rect 19762 4924 19826 4928
rect 19762 4868 19766 4924
rect 19766 4868 19822 4924
rect 19822 4868 19826 4924
rect 19762 4864 19826 4868
rect 26950 4924 27014 4928
rect 26950 4868 26954 4924
rect 26954 4868 27010 4924
rect 27010 4868 27014 4924
rect 26950 4864 27014 4868
rect 27030 4924 27094 4928
rect 27030 4868 27034 4924
rect 27034 4868 27090 4924
rect 27090 4868 27094 4924
rect 27030 4864 27094 4868
rect 27110 4924 27174 4928
rect 27110 4868 27114 4924
rect 27114 4868 27170 4924
rect 27170 4868 27174 4924
rect 27110 4864 27174 4868
rect 27190 4924 27254 4928
rect 27190 4868 27194 4924
rect 27194 4868 27250 4924
rect 27250 4868 27254 4924
rect 27190 4864 27254 4868
rect 5326 4380 5390 4384
rect 5326 4324 5330 4380
rect 5330 4324 5386 4380
rect 5386 4324 5390 4380
rect 5326 4320 5390 4324
rect 5406 4380 5470 4384
rect 5406 4324 5410 4380
rect 5410 4324 5466 4380
rect 5466 4324 5470 4380
rect 5406 4320 5470 4324
rect 5486 4380 5550 4384
rect 5486 4324 5490 4380
rect 5490 4324 5546 4380
rect 5546 4324 5550 4380
rect 5486 4320 5550 4324
rect 5566 4380 5630 4384
rect 5566 4324 5570 4380
rect 5570 4324 5626 4380
rect 5626 4324 5630 4380
rect 5566 4320 5630 4324
rect 12754 4380 12818 4384
rect 12754 4324 12758 4380
rect 12758 4324 12814 4380
rect 12814 4324 12818 4380
rect 12754 4320 12818 4324
rect 12834 4380 12898 4384
rect 12834 4324 12838 4380
rect 12838 4324 12894 4380
rect 12894 4324 12898 4380
rect 12834 4320 12898 4324
rect 12914 4380 12978 4384
rect 12914 4324 12918 4380
rect 12918 4324 12974 4380
rect 12974 4324 12978 4380
rect 12914 4320 12978 4324
rect 12994 4380 13058 4384
rect 12994 4324 12998 4380
rect 12998 4324 13054 4380
rect 13054 4324 13058 4380
rect 12994 4320 13058 4324
rect 20182 4380 20246 4384
rect 20182 4324 20186 4380
rect 20186 4324 20242 4380
rect 20242 4324 20246 4380
rect 20182 4320 20246 4324
rect 20262 4380 20326 4384
rect 20262 4324 20266 4380
rect 20266 4324 20322 4380
rect 20322 4324 20326 4380
rect 20262 4320 20326 4324
rect 20342 4380 20406 4384
rect 20342 4324 20346 4380
rect 20346 4324 20402 4380
rect 20402 4324 20406 4380
rect 20342 4320 20406 4324
rect 20422 4380 20486 4384
rect 20422 4324 20426 4380
rect 20426 4324 20482 4380
rect 20482 4324 20486 4380
rect 20422 4320 20486 4324
rect 27610 4380 27674 4384
rect 27610 4324 27614 4380
rect 27614 4324 27670 4380
rect 27670 4324 27674 4380
rect 27610 4320 27674 4324
rect 27690 4380 27754 4384
rect 27690 4324 27694 4380
rect 27694 4324 27750 4380
rect 27750 4324 27754 4380
rect 27690 4320 27754 4324
rect 27770 4380 27834 4384
rect 27770 4324 27774 4380
rect 27774 4324 27830 4380
rect 27830 4324 27834 4380
rect 27770 4320 27834 4324
rect 27850 4380 27914 4384
rect 27850 4324 27854 4380
rect 27854 4324 27910 4380
rect 27910 4324 27914 4380
rect 27850 4320 27914 4324
rect 4666 3836 4730 3840
rect 4666 3780 4670 3836
rect 4670 3780 4726 3836
rect 4726 3780 4730 3836
rect 4666 3776 4730 3780
rect 4746 3836 4810 3840
rect 4746 3780 4750 3836
rect 4750 3780 4806 3836
rect 4806 3780 4810 3836
rect 4746 3776 4810 3780
rect 4826 3836 4890 3840
rect 4826 3780 4830 3836
rect 4830 3780 4886 3836
rect 4886 3780 4890 3836
rect 4826 3776 4890 3780
rect 4906 3836 4970 3840
rect 4906 3780 4910 3836
rect 4910 3780 4966 3836
rect 4966 3780 4970 3836
rect 4906 3776 4970 3780
rect 12094 3836 12158 3840
rect 12094 3780 12098 3836
rect 12098 3780 12154 3836
rect 12154 3780 12158 3836
rect 12094 3776 12158 3780
rect 12174 3836 12238 3840
rect 12174 3780 12178 3836
rect 12178 3780 12234 3836
rect 12234 3780 12238 3836
rect 12174 3776 12238 3780
rect 12254 3836 12318 3840
rect 12254 3780 12258 3836
rect 12258 3780 12314 3836
rect 12314 3780 12318 3836
rect 12254 3776 12318 3780
rect 12334 3836 12398 3840
rect 12334 3780 12338 3836
rect 12338 3780 12394 3836
rect 12394 3780 12398 3836
rect 12334 3776 12398 3780
rect 19522 3836 19586 3840
rect 19522 3780 19526 3836
rect 19526 3780 19582 3836
rect 19582 3780 19586 3836
rect 19522 3776 19586 3780
rect 19602 3836 19666 3840
rect 19602 3780 19606 3836
rect 19606 3780 19662 3836
rect 19662 3780 19666 3836
rect 19602 3776 19666 3780
rect 19682 3836 19746 3840
rect 19682 3780 19686 3836
rect 19686 3780 19742 3836
rect 19742 3780 19746 3836
rect 19682 3776 19746 3780
rect 19762 3836 19826 3840
rect 19762 3780 19766 3836
rect 19766 3780 19822 3836
rect 19822 3780 19826 3836
rect 19762 3776 19826 3780
rect 26950 3836 27014 3840
rect 26950 3780 26954 3836
rect 26954 3780 27010 3836
rect 27010 3780 27014 3836
rect 26950 3776 27014 3780
rect 27030 3836 27094 3840
rect 27030 3780 27034 3836
rect 27034 3780 27090 3836
rect 27090 3780 27094 3836
rect 27030 3776 27094 3780
rect 27110 3836 27174 3840
rect 27110 3780 27114 3836
rect 27114 3780 27170 3836
rect 27170 3780 27174 3836
rect 27110 3776 27174 3780
rect 27190 3836 27254 3840
rect 27190 3780 27194 3836
rect 27194 3780 27250 3836
rect 27250 3780 27254 3836
rect 27190 3776 27254 3780
rect 5326 3292 5390 3296
rect 5326 3236 5330 3292
rect 5330 3236 5386 3292
rect 5386 3236 5390 3292
rect 5326 3232 5390 3236
rect 5406 3292 5470 3296
rect 5406 3236 5410 3292
rect 5410 3236 5466 3292
rect 5466 3236 5470 3292
rect 5406 3232 5470 3236
rect 5486 3292 5550 3296
rect 5486 3236 5490 3292
rect 5490 3236 5546 3292
rect 5546 3236 5550 3292
rect 5486 3232 5550 3236
rect 5566 3292 5630 3296
rect 5566 3236 5570 3292
rect 5570 3236 5626 3292
rect 5626 3236 5630 3292
rect 5566 3232 5630 3236
rect 12754 3292 12818 3296
rect 12754 3236 12758 3292
rect 12758 3236 12814 3292
rect 12814 3236 12818 3292
rect 12754 3232 12818 3236
rect 12834 3292 12898 3296
rect 12834 3236 12838 3292
rect 12838 3236 12894 3292
rect 12894 3236 12898 3292
rect 12834 3232 12898 3236
rect 12914 3292 12978 3296
rect 12914 3236 12918 3292
rect 12918 3236 12974 3292
rect 12974 3236 12978 3292
rect 12914 3232 12978 3236
rect 12994 3292 13058 3296
rect 12994 3236 12998 3292
rect 12998 3236 13054 3292
rect 13054 3236 13058 3292
rect 12994 3232 13058 3236
rect 20182 3292 20246 3296
rect 20182 3236 20186 3292
rect 20186 3236 20242 3292
rect 20242 3236 20246 3292
rect 20182 3232 20246 3236
rect 20262 3292 20326 3296
rect 20262 3236 20266 3292
rect 20266 3236 20322 3292
rect 20322 3236 20326 3292
rect 20262 3232 20326 3236
rect 20342 3292 20406 3296
rect 20342 3236 20346 3292
rect 20346 3236 20402 3292
rect 20402 3236 20406 3292
rect 20342 3232 20406 3236
rect 20422 3292 20486 3296
rect 20422 3236 20426 3292
rect 20426 3236 20482 3292
rect 20482 3236 20486 3292
rect 20422 3232 20486 3236
rect 27610 3292 27674 3296
rect 27610 3236 27614 3292
rect 27614 3236 27670 3292
rect 27670 3236 27674 3292
rect 27610 3232 27674 3236
rect 27690 3292 27754 3296
rect 27690 3236 27694 3292
rect 27694 3236 27750 3292
rect 27750 3236 27754 3292
rect 27690 3232 27754 3236
rect 27770 3292 27834 3296
rect 27770 3236 27774 3292
rect 27774 3236 27830 3292
rect 27830 3236 27834 3292
rect 27770 3232 27834 3236
rect 27850 3292 27914 3296
rect 27850 3236 27854 3292
rect 27854 3236 27910 3292
rect 27910 3236 27914 3292
rect 27850 3232 27914 3236
rect 4666 2748 4730 2752
rect 4666 2692 4670 2748
rect 4670 2692 4726 2748
rect 4726 2692 4730 2748
rect 4666 2688 4730 2692
rect 4746 2748 4810 2752
rect 4746 2692 4750 2748
rect 4750 2692 4806 2748
rect 4806 2692 4810 2748
rect 4746 2688 4810 2692
rect 4826 2748 4890 2752
rect 4826 2692 4830 2748
rect 4830 2692 4886 2748
rect 4886 2692 4890 2748
rect 4826 2688 4890 2692
rect 4906 2748 4970 2752
rect 4906 2692 4910 2748
rect 4910 2692 4966 2748
rect 4966 2692 4970 2748
rect 4906 2688 4970 2692
rect 12094 2748 12158 2752
rect 12094 2692 12098 2748
rect 12098 2692 12154 2748
rect 12154 2692 12158 2748
rect 12094 2688 12158 2692
rect 12174 2748 12238 2752
rect 12174 2692 12178 2748
rect 12178 2692 12234 2748
rect 12234 2692 12238 2748
rect 12174 2688 12238 2692
rect 12254 2748 12318 2752
rect 12254 2692 12258 2748
rect 12258 2692 12314 2748
rect 12314 2692 12318 2748
rect 12254 2688 12318 2692
rect 12334 2748 12398 2752
rect 12334 2692 12338 2748
rect 12338 2692 12394 2748
rect 12394 2692 12398 2748
rect 12334 2688 12398 2692
rect 19522 2748 19586 2752
rect 19522 2692 19526 2748
rect 19526 2692 19582 2748
rect 19582 2692 19586 2748
rect 19522 2688 19586 2692
rect 19602 2748 19666 2752
rect 19602 2692 19606 2748
rect 19606 2692 19662 2748
rect 19662 2692 19666 2748
rect 19602 2688 19666 2692
rect 19682 2748 19746 2752
rect 19682 2692 19686 2748
rect 19686 2692 19742 2748
rect 19742 2692 19746 2748
rect 19682 2688 19746 2692
rect 19762 2748 19826 2752
rect 19762 2692 19766 2748
rect 19766 2692 19822 2748
rect 19822 2692 19826 2748
rect 19762 2688 19826 2692
rect 26950 2748 27014 2752
rect 26950 2692 26954 2748
rect 26954 2692 27010 2748
rect 27010 2692 27014 2748
rect 26950 2688 27014 2692
rect 27030 2748 27094 2752
rect 27030 2692 27034 2748
rect 27034 2692 27090 2748
rect 27090 2692 27094 2748
rect 27030 2688 27094 2692
rect 27110 2748 27174 2752
rect 27110 2692 27114 2748
rect 27114 2692 27170 2748
rect 27170 2692 27174 2748
rect 27110 2688 27174 2692
rect 27190 2748 27254 2752
rect 27190 2692 27194 2748
rect 27194 2692 27250 2748
rect 27250 2692 27254 2748
rect 27190 2688 27254 2692
rect 5326 2204 5390 2208
rect 5326 2148 5330 2204
rect 5330 2148 5386 2204
rect 5386 2148 5390 2204
rect 5326 2144 5390 2148
rect 5406 2204 5470 2208
rect 5406 2148 5410 2204
rect 5410 2148 5466 2204
rect 5466 2148 5470 2204
rect 5406 2144 5470 2148
rect 5486 2204 5550 2208
rect 5486 2148 5490 2204
rect 5490 2148 5546 2204
rect 5546 2148 5550 2204
rect 5486 2144 5550 2148
rect 5566 2204 5630 2208
rect 5566 2148 5570 2204
rect 5570 2148 5626 2204
rect 5626 2148 5630 2204
rect 5566 2144 5630 2148
rect 12754 2204 12818 2208
rect 12754 2148 12758 2204
rect 12758 2148 12814 2204
rect 12814 2148 12818 2204
rect 12754 2144 12818 2148
rect 12834 2204 12898 2208
rect 12834 2148 12838 2204
rect 12838 2148 12894 2204
rect 12894 2148 12898 2204
rect 12834 2144 12898 2148
rect 12914 2204 12978 2208
rect 12914 2148 12918 2204
rect 12918 2148 12974 2204
rect 12974 2148 12978 2204
rect 12914 2144 12978 2148
rect 12994 2204 13058 2208
rect 12994 2148 12998 2204
rect 12998 2148 13054 2204
rect 13054 2148 13058 2204
rect 12994 2144 13058 2148
rect 20182 2204 20246 2208
rect 20182 2148 20186 2204
rect 20186 2148 20242 2204
rect 20242 2148 20246 2204
rect 20182 2144 20246 2148
rect 20262 2204 20326 2208
rect 20262 2148 20266 2204
rect 20266 2148 20322 2204
rect 20322 2148 20326 2204
rect 20262 2144 20326 2148
rect 20342 2204 20406 2208
rect 20342 2148 20346 2204
rect 20346 2148 20402 2204
rect 20402 2148 20406 2204
rect 20342 2144 20406 2148
rect 20422 2204 20486 2208
rect 20422 2148 20426 2204
rect 20426 2148 20482 2204
rect 20482 2148 20486 2204
rect 20422 2144 20486 2148
rect 27610 2204 27674 2208
rect 27610 2148 27614 2204
rect 27614 2148 27670 2204
rect 27670 2148 27674 2204
rect 27610 2144 27674 2148
rect 27690 2204 27754 2208
rect 27690 2148 27694 2204
rect 27694 2148 27750 2204
rect 27750 2148 27754 2204
rect 27690 2144 27754 2148
rect 27770 2204 27834 2208
rect 27770 2148 27774 2204
rect 27774 2148 27830 2204
rect 27830 2148 27834 2204
rect 27770 2144 27834 2148
rect 27850 2204 27914 2208
rect 27850 2148 27854 2204
rect 27854 2148 27910 2204
rect 27910 2148 27914 2204
rect 27850 2144 27914 2148
<< metal4 >>
rect 4658 28864 4978 29424
rect 4658 28800 4666 28864
rect 4730 28800 4746 28864
rect 4810 28800 4826 28864
rect 4890 28800 4906 28864
rect 4970 28800 4978 28864
rect 4658 27776 4978 28800
rect 4658 27712 4666 27776
rect 4730 27712 4746 27776
rect 4810 27712 4826 27776
rect 4890 27712 4906 27776
rect 4970 27712 4978 27776
rect 4658 26688 4978 27712
rect 4658 26624 4666 26688
rect 4730 26624 4746 26688
rect 4810 26624 4826 26688
rect 4890 26624 4906 26688
rect 4970 26624 4978 26688
rect 4658 26094 4978 26624
rect 4658 25858 4700 26094
rect 4936 25858 4978 26094
rect 4658 25600 4978 25858
rect 4658 25536 4666 25600
rect 4730 25536 4746 25600
rect 4810 25536 4826 25600
rect 4890 25536 4906 25600
rect 4970 25536 4978 25600
rect 4658 24512 4978 25536
rect 4658 24448 4666 24512
rect 4730 24448 4746 24512
rect 4810 24448 4826 24512
rect 4890 24448 4906 24512
rect 4970 24448 4978 24512
rect 4658 23424 4978 24448
rect 4658 23360 4666 23424
rect 4730 23360 4746 23424
rect 4810 23360 4826 23424
rect 4890 23360 4906 23424
rect 4970 23360 4978 23424
rect 4658 22336 4978 23360
rect 4658 22272 4666 22336
rect 4730 22272 4746 22336
rect 4810 22272 4826 22336
rect 4890 22272 4906 22336
rect 4970 22272 4978 22336
rect 4658 21248 4978 22272
rect 4658 21184 4666 21248
rect 4730 21184 4746 21248
rect 4810 21184 4826 21248
rect 4890 21184 4906 21248
rect 4970 21184 4978 21248
rect 4658 20160 4978 21184
rect 4658 20096 4666 20160
rect 4730 20096 4746 20160
rect 4810 20096 4826 20160
rect 4890 20096 4906 20160
rect 4970 20096 4978 20160
rect 4658 19294 4978 20096
rect 4658 19072 4700 19294
rect 4936 19072 4978 19294
rect 4658 19008 4666 19072
rect 4730 19008 4746 19058
rect 4810 19008 4826 19058
rect 4890 19008 4906 19058
rect 4970 19008 4978 19072
rect 4658 17984 4978 19008
rect 4658 17920 4666 17984
rect 4730 17920 4746 17984
rect 4810 17920 4826 17984
rect 4890 17920 4906 17984
rect 4970 17920 4978 17984
rect 4658 16896 4978 17920
rect 4658 16832 4666 16896
rect 4730 16832 4746 16896
rect 4810 16832 4826 16896
rect 4890 16832 4906 16896
rect 4970 16832 4978 16896
rect 4658 15808 4978 16832
rect 4658 15744 4666 15808
rect 4730 15744 4746 15808
rect 4810 15744 4826 15808
rect 4890 15744 4906 15808
rect 4970 15744 4978 15808
rect 4658 14720 4978 15744
rect 4658 14656 4666 14720
rect 4730 14656 4746 14720
rect 4810 14656 4826 14720
rect 4890 14656 4906 14720
rect 4970 14656 4978 14720
rect 4658 13632 4978 14656
rect 4658 13568 4666 13632
rect 4730 13568 4746 13632
rect 4810 13568 4826 13632
rect 4890 13568 4906 13632
rect 4970 13568 4978 13632
rect 4658 12544 4978 13568
rect 4658 12480 4666 12544
rect 4730 12494 4746 12544
rect 4810 12494 4826 12544
rect 4890 12494 4906 12544
rect 4970 12480 4978 12544
rect 4658 12258 4700 12480
rect 4936 12258 4978 12480
rect 4658 11456 4978 12258
rect 4658 11392 4666 11456
rect 4730 11392 4746 11456
rect 4810 11392 4826 11456
rect 4890 11392 4906 11456
rect 4970 11392 4978 11456
rect 4658 10368 4978 11392
rect 4658 10304 4666 10368
rect 4730 10304 4746 10368
rect 4810 10304 4826 10368
rect 4890 10304 4906 10368
rect 4970 10304 4978 10368
rect 4658 9280 4978 10304
rect 4658 9216 4666 9280
rect 4730 9216 4746 9280
rect 4810 9216 4826 9280
rect 4890 9216 4906 9280
rect 4970 9216 4978 9280
rect 4658 8192 4978 9216
rect 4658 8128 4666 8192
rect 4730 8128 4746 8192
rect 4810 8128 4826 8192
rect 4890 8128 4906 8192
rect 4970 8128 4978 8192
rect 4658 7104 4978 8128
rect 4658 7040 4666 7104
rect 4730 7040 4746 7104
rect 4810 7040 4826 7104
rect 4890 7040 4906 7104
rect 4970 7040 4978 7104
rect 4658 6016 4978 7040
rect 4658 5952 4666 6016
rect 4730 5952 4746 6016
rect 4810 5952 4826 6016
rect 4890 5952 4906 6016
rect 4970 5952 4978 6016
rect 4658 5694 4978 5952
rect 4658 5458 4700 5694
rect 4936 5458 4978 5694
rect 4658 4928 4978 5458
rect 4658 4864 4666 4928
rect 4730 4864 4746 4928
rect 4810 4864 4826 4928
rect 4890 4864 4906 4928
rect 4970 4864 4978 4928
rect 4658 3840 4978 4864
rect 4658 3776 4666 3840
rect 4730 3776 4746 3840
rect 4810 3776 4826 3840
rect 4890 3776 4906 3840
rect 4970 3776 4978 3840
rect 4658 2752 4978 3776
rect 4658 2688 4666 2752
rect 4730 2688 4746 2752
rect 4810 2688 4826 2752
rect 4890 2688 4906 2752
rect 4970 2688 4978 2752
rect 4658 2128 4978 2688
rect 5318 29408 5638 29424
rect 5318 29344 5326 29408
rect 5390 29344 5406 29408
rect 5470 29344 5486 29408
rect 5550 29344 5566 29408
rect 5630 29344 5638 29408
rect 5318 28320 5638 29344
rect 5318 28256 5326 28320
rect 5390 28256 5406 28320
rect 5470 28256 5486 28320
rect 5550 28256 5566 28320
rect 5630 28256 5638 28320
rect 5318 27232 5638 28256
rect 5318 27168 5326 27232
rect 5390 27168 5406 27232
rect 5470 27168 5486 27232
rect 5550 27168 5566 27232
rect 5630 27168 5638 27232
rect 5318 26754 5638 27168
rect 5318 26518 5360 26754
rect 5596 26518 5638 26754
rect 5318 26144 5638 26518
rect 5318 26080 5326 26144
rect 5390 26080 5406 26144
rect 5470 26080 5486 26144
rect 5550 26080 5566 26144
rect 5630 26080 5638 26144
rect 5318 25056 5638 26080
rect 5318 24992 5326 25056
rect 5390 24992 5406 25056
rect 5470 24992 5486 25056
rect 5550 24992 5566 25056
rect 5630 24992 5638 25056
rect 5318 23968 5638 24992
rect 5318 23904 5326 23968
rect 5390 23904 5406 23968
rect 5470 23904 5486 23968
rect 5550 23904 5566 23968
rect 5630 23904 5638 23968
rect 5318 22880 5638 23904
rect 5318 22816 5326 22880
rect 5390 22816 5406 22880
rect 5470 22816 5486 22880
rect 5550 22816 5566 22880
rect 5630 22816 5638 22880
rect 5318 21792 5638 22816
rect 5318 21728 5326 21792
rect 5390 21728 5406 21792
rect 5470 21728 5486 21792
rect 5550 21728 5566 21792
rect 5630 21728 5638 21792
rect 5318 20704 5638 21728
rect 5318 20640 5326 20704
rect 5390 20640 5406 20704
rect 5470 20640 5486 20704
rect 5550 20640 5566 20704
rect 5630 20640 5638 20704
rect 5318 19954 5638 20640
rect 5318 19718 5360 19954
rect 5596 19718 5638 19954
rect 5318 19616 5638 19718
rect 5318 19552 5326 19616
rect 5390 19552 5406 19616
rect 5470 19552 5486 19616
rect 5550 19552 5566 19616
rect 5630 19552 5638 19616
rect 5318 18528 5638 19552
rect 5318 18464 5326 18528
rect 5390 18464 5406 18528
rect 5470 18464 5486 18528
rect 5550 18464 5566 18528
rect 5630 18464 5638 18528
rect 5318 17440 5638 18464
rect 5318 17376 5326 17440
rect 5390 17376 5406 17440
rect 5470 17376 5486 17440
rect 5550 17376 5566 17440
rect 5630 17376 5638 17440
rect 5318 16352 5638 17376
rect 5318 16288 5326 16352
rect 5390 16288 5406 16352
rect 5470 16288 5486 16352
rect 5550 16288 5566 16352
rect 5630 16288 5638 16352
rect 5318 15264 5638 16288
rect 5318 15200 5326 15264
rect 5390 15200 5406 15264
rect 5470 15200 5486 15264
rect 5550 15200 5566 15264
rect 5630 15200 5638 15264
rect 5318 14176 5638 15200
rect 5318 14112 5326 14176
rect 5390 14112 5406 14176
rect 5470 14112 5486 14176
rect 5550 14112 5566 14176
rect 5630 14112 5638 14176
rect 5318 13154 5638 14112
rect 5318 13088 5360 13154
rect 5596 13088 5638 13154
rect 5318 13024 5326 13088
rect 5630 13024 5638 13088
rect 5318 12918 5360 13024
rect 5596 12918 5638 13024
rect 5318 12000 5638 12918
rect 5318 11936 5326 12000
rect 5390 11936 5406 12000
rect 5470 11936 5486 12000
rect 5550 11936 5566 12000
rect 5630 11936 5638 12000
rect 5318 10912 5638 11936
rect 5318 10848 5326 10912
rect 5390 10848 5406 10912
rect 5470 10848 5486 10912
rect 5550 10848 5566 10912
rect 5630 10848 5638 10912
rect 5318 9824 5638 10848
rect 5318 9760 5326 9824
rect 5390 9760 5406 9824
rect 5470 9760 5486 9824
rect 5550 9760 5566 9824
rect 5630 9760 5638 9824
rect 5318 8736 5638 9760
rect 5318 8672 5326 8736
rect 5390 8672 5406 8736
rect 5470 8672 5486 8736
rect 5550 8672 5566 8736
rect 5630 8672 5638 8736
rect 5318 7648 5638 8672
rect 5318 7584 5326 7648
rect 5390 7584 5406 7648
rect 5470 7584 5486 7648
rect 5550 7584 5566 7648
rect 5630 7584 5638 7648
rect 5318 6560 5638 7584
rect 5318 6496 5326 6560
rect 5390 6496 5406 6560
rect 5470 6496 5486 6560
rect 5550 6496 5566 6560
rect 5630 6496 5638 6560
rect 5318 6354 5638 6496
rect 5318 6118 5360 6354
rect 5596 6118 5638 6354
rect 5318 5472 5638 6118
rect 5318 5408 5326 5472
rect 5390 5408 5406 5472
rect 5470 5408 5486 5472
rect 5550 5408 5566 5472
rect 5630 5408 5638 5472
rect 5318 4384 5638 5408
rect 5318 4320 5326 4384
rect 5390 4320 5406 4384
rect 5470 4320 5486 4384
rect 5550 4320 5566 4384
rect 5630 4320 5638 4384
rect 5318 3296 5638 4320
rect 5318 3232 5326 3296
rect 5390 3232 5406 3296
rect 5470 3232 5486 3296
rect 5550 3232 5566 3296
rect 5630 3232 5638 3296
rect 5318 2208 5638 3232
rect 5318 2144 5326 2208
rect 5390 2144 5406 2208
rect 5470 2144 5486 2208
rect 5550 2144 5566 2208
rect 5630 2144 5638 2208
rect 5318 2128 5638 2144
rect 12086 28864 12406 29424
rect 12086 28800 12094 28864
rect 12158 28800 12174 28864
rect 12238 28800 12254 28864
rect 12318 28800 12334 28864
rect 12398 28800 12406 28864
rect 12086 27776 12406 28800
rect 12086 27712 12094 27776
rect 12158 27712 12174 27776
rect 12238 27712 12254 27776
rect 12318 27712 12334 27776
rect 12398 27712 12406 27776
rect 12086 26688 12406 27712
rect 12086 26624 12094 26688
rect 12158 26624 12174 26688
rect 12238 26624 12254 26688
rect 12318 26624 12334 26688
rect 12398 26624 12406 26688
rect 12086 26094 12406 26624
rect 12086 25858 12128 26094
rect 12364 25858 12406 26094
rect 12086 25600 12406 25858
rect 12086 25536 12094 25600
rect 12158 25536 12174 25600
rect 12238 25536 12254 25600
rect 12318 25536 12334 25600
rect 12398 25536 12406 25600
rect 12086 24512 12406 25536
rect 12086 24448 12094 24512
rect 12158 24448 12174 24512
rect 12238 24448 12254 24512
rect 12318 24448 12334 24512
rect 12398 24448 12406 24512
rect 12086 23424 12406 24448
rect 12086 23360 12094 23424
rect 12158 23360 12174 23424
rect 12238 23360 12254 23424
rect 12318 23360 12334 23424
rect 12398 23360 12406 23424
rect 12086 22336 12406 23360
rect 12086 22272 12094 22336
rect 12158 22272 12174 22336
rect 12238 22272 12254 22336
rect 12318 22272 12334 22336
rect 12398 22272 12406 22336
rect 12086 21248 12406 22272
rect 12086 21184 12094 21248
rect 12158 21184 12174 21248
rect 12238 21184 12254 21248
rect 12318 21184 12334 21248
rect 12398 21184 12406 21248
rect 12086 20160 12406 21184
rect 12086 20096 12094 20160
rect 12158 20096 12174 20160
rect 12238 20096 12254 20160
rect 12318 20096 12334 20160
rect 12398 20096 12406 20160
rect 12086 19294 12406 20096
rect 12086 19072 12128 19294
rect 12364 19072 12406 19294
rect 12086 19008 12094 19072
rect 12158 19008 12174 19058
rect 12238 19008 12254 19058
rect 12318 19008 12334 19058
rect 12398 19008 12406 19072
rect 12086 17984 12406 19008
rect 12086 17920 12094 17984
rect 12158 17920 12174 17984
rect 12238 17920 12254 17984
rect 12318 17920 12334 17984
rect 12398 17920 12406 17984
rect 12086 16896 12406 17920
rect 12086 16832 12094 16896
rect 12158 16832 12174 16896
rect 12238 16832 12254 16896
rect 12318 16832 12334 16896
rect 12398 16832 12406 16896
rect 12086 15808 12406 16832
rect 12086 15744 12094 15808
rect 12158 15744 12174 15808
rect 12238 15744 12254 15808
rect 12318 15744 12334 15808
rect 12398 15744 12406 15808
rect 12086 14720 12406 15744
rect 12086 14656 12094 14720
rect 12158 14656 12174 14720
rect 12238 14656 12254 14720
rect 12318 14656 12334 14720
rect 12398 14656 12406 14720
rect 12086 13632 12406 14656
rect 12086 13568 12094 13632
rect 12158 13568 12174 13632
rect 12238 13568 12254 13632
rect 12318 13568 12334 13632
rect 12398 13568 12406 13632
rect 12086 12544 12406 13568
rect 12086 12480 12094 12544
rect 12158 12494 12174 12544
rect 12238 12494 12254 12544
rect 12318 12494 12334 12544
rect 12398 12480 12406 12544
rect 12086 12258 12128 12480
rect 12364 12258 12406 12480
rect 12086 11456 12406 12258
rect 12086 11392 12094 11456
rect 12158 11392 12174 11456
rect 12238 11392 12254 11456
rect 12318 11392 12334 11456
rect 12398 11392 12406 11456
rect 12086 10368 12406 11392
rect 12086 10304 12094 10368
rect 12158 10304 12174 10368
rect 12238 10304 12254 10368
rect 12318 10304 12334 10368
rect 12398 10304 12406 10368
rect 12086 9280 12406 10304
rect 12086 9216 12094 9280
rect 12158 9216 12174 9280
rect 12238 9216 12254 9280
rect 12318 9216 12334 9280
rect 12398 9216 12406 9280
rect 12086 8192 12406 9216
rect 12086 8128 12094 8192
rect 12158 8128 12174 8192
rect 12238 8128 12254 8192
rect 12318 8128 12334 8192
rect 12398 8128 12406 8192
rect 12086 7104 12406 8128
rect 12086 7040 12094 7104
rect 12158 7040 12174 7104
rect 12238 7040 12254 7104
rect 12318 7040 12334 7104
rect 12398 7040 12406 7104
rect 12086 6016 12406 7040
rect 12086 5952 12094 6016
rect 12158 5952 12174 6016
rect 12238 5952 12254 6016
rect 12318 5952 12334 6016
rect 12398 5952 12406 6016
rect 12086 5694 12406 5952
rect 12086 5458 12128 5694
rect 12364 5458 12406 5694
rect 12086 4928 12406 5458
rect 12086 4864 12094 4928
rect 12158 4864 12174 4928
rect 12238 4864 12254 4928
rect 12318 4864 12334 4928
rect 12398 4864 12406 4928
rect 12086 3840 12406 4864
rect 12086 3776 12094 3840
rect 12158 3776 12174 3840
rect 12238 3776 12254 3840
rect 12318 3776 12334 3840
rect 12398 3776 12406 3840
rect 12086 2752 12406 3776
rect 12086 2688 12094 2752
rect 12158 2688 12174 2752
rect 12238 2688 12254 2752
rect 12318 2688 12334 2752
rect 12398 2688 12406 2752
rect 12086 2128 12406 2688
rect 12746 29408 13066 29424
rect 12746 29344 12754 29408
rect 12818 29344 12834 29408
rect 12898 29344 12914 29408
rect 12978 29344 12994 29408
rect 13058 29344 13066 29408
rect 12746 28320 13066 29344
rect 12746 28256 12754 28320
rect 12818 28256 12834 28320
rect 12898 28256 12914 28320
rect 12978 28256 12994 28320
rect 13058 28256 13066 28320
rect 12746 27232 13066 28256
rect 12746 27168 12754 27232
rect 12818 27168 12834 27232
rect 12898 27168 12914 27232
rect 12978 27168 12994 27232
rect 13058 27168 13066 27232
rect 12746 26754 13066 27168
rect 12746 26518 12788 26754
rect 13024 26518 13066 26754
rect 12746 26144 13066 26518
rect 12746 26080 12754 26144
rect 12818 26080 12834 26144
rect 12898 26080 12914 26144
rect 12978 26080 12994 26144
rect 13058 26080 13066 26144
rect 12746 25056 13066 26080
rect 12746 24992 12754 25056
rect 12818 24992 12834 25056
rect 12898 24992 12914 25056
rect 12978 24992 12994 25056
rect 13058 24992 13066 25056
rect 12746 23968 13066 24992
rect 12746 23904 12754 23968
rect 12818 23904 12834 23968
rect 12898 23904 12914 23968
rect 12978 23904 12994 23968
rect 13058 23904 13066 23968
rect 12746 22880 13066 23904
rect 12746 22816 12754 22880
rect 12818 22816 12834 22880
rect 12898 22816 12914 22880
rect 12978 22816 12994 22880
rect 13058 22816 13066 22880
rect 12746 21792 13066 22816
rect 12746 21728 12754 21792
rect 12818 21728 12834 21792
rect 12898 21728 12914 21792
rect 12978 21728 12994 21792
rect 13058 21728 13066 21792
rect 12746 20704 13066 21728
rect 12746 20640 12754 20704
rect 12818 20640 12834 20704
rect 12898 20640 12914 20704
rect 12978 20640 12994 20704
rect 13058 20640 13066 20704
rect 12746 19954 13066 20640
rect 12746 19718 12788 19954
rect 13024 19718 13066 19954
rect 12746 19616 13066 19718
rect 12746 19552 12754 19616
rect 12818 19552 12834 19616
rect 12898 19552 12914 19616
rect 12978 19552 12994 19616
rect 13058 19552 13066 19616
rect 12746 18528 13066 19552
rect 12746 18464 12754 18528
rect 12818 18464 12834 18528
rect 12898 18464 12914 18528
rect 12978 18464 12994 18528
rect 13058 18464 13066 18528
rect 12746 17440 13066 18464
rect 12746 17376 12754 17440
rect 12818 17376 12834 17440
rect 12898 17376 12914 17440
rect 12978 17376 12994 17440
rect 13058 17376 13066 17440
rect 12746 16352 13066 17376
rect 12746 16288 12754 16352
rect 12818 16288 12834 16352
rect 12898 16288 12914 16352
rect 12978 16288 12994 16352
rect 13058 16288 13066 16352
rect 12746 15264 13066 16288
rect 12746 15200 12754 15264
rect 12818 15200 12834 15264
rect 12898 15200 12914 15264
rect 12978 15200 12994 15264
rect 13058 15200 13066 15264
rect 12746 14176 13066 15200
rect 12746 14112 12754 14176
rect 12818 14112 12834 14176
rect 12898 14112 12914 14176
rect 12978 14112 12994 14176
rect 13058 14112 13066 14176
rect 12746 13154 13066 14112
rect 12746 13088 12788 13154
rect 13024 13088 13066 13154
rect 12746 13024 12754 13088
rect 13058 13024 13066 13088
rect 12746 12918 12788 13024
rect 13024 12918 13066 13024
rect 12746 12000 13066 12918
rect 12746 11936 12754 12000
rect 12818 11936 12834 12000
rect 12898 11936 12914 12000
rect 12978 11936 12994 12000
rect 13058 11936 13066 12000
rect 12746 10912 13066 11936
rect 12746 10848 12754 10912
rect 12818 10848 12834 10912
rect 12898 10848 12914 10912
rect 12978 10848 12994 10912
rect 13058 10848 13066 10912
rect 12746 9824 13066 10848
rect 12746 9760 12754 9824
rect 12818 9760 12834 9824
rect 12898 9760 12914 9824
rect 12978 9760 12994 9824
rect 13058 9760 13066 9824
rect 12746 8736 13066 9760
rect 12746 8672 12754 8736
rect 12818 8672 12834 8736
rect 12898 8672 12914 8736
rect 12978 8672 12994 8736
rect 13058 8672 13066 8736
rect 12746 7648 13066 8672
rect 12746 7584 12754 7648
rect 12818 7584 12834 7648
rect 12898 7584 12914 7648
rect 12978 7584 12994 7648
rect 13058 7584 13066 7648
rect 12746 6560 13066 7584
rect 12746 6496 12754 6560
rect 12818 6496 12834 6560
rect 12898 6496 12914 6560
rect 12978 6496 12994 6560
rect 13058 6496 13066 6560
rect 12746 6354 13066 6496
rect 12746 6118 12788 6354
rect 13024 6118 13066 6354
rect 12746 5472 13066 6118
rect 12746 5408 12754 5472
rect 12818 5408 12834 5472
rect 12898 5408 12914 5472
rect 12978 5408 12994 5472
rect 13058 5408 13066 5472
rect 12746 4384 13066 5408
rect 12746 4320 12754 4384
rect 12818 4320 12834 4384
rect 12898 4320 12914 4384
rect 12978 4320 12994 4384
rect 13058 4320 13066 4384
rect 12746 3296 13066 4320
rect 12746 3232 12754 3296
rect 12818 3232 12834 3296
rect 12898 3232 12914 3296
rect 12978 3232 12994 3296
rect 13058 3232 13066 3296
rect 12746 2208 13066 3232
rect 12746 2144 12754 2208
rect 12818 2144 12834 2208
rect 12898 2144 12914 2208
rect 12978 2144 12994 2208
rect 13058 2144 13066 2208
rect 12746 2128 13066 2144
rect 19514 28864 19834 29424
rect 19514 28800 19522 28864
rect 19586 28800 19602 28864
rect 19666 28800 19682 28864
rect 19746 28800 19762 28864
rect 19826 28800 19834 28864
rect 19514 27776 19834 28800
rect 19514 27712 19522 27776
rect 19586 27712 19602 27776
rect 19666 27712 19682 27776
rect 19746 27712 19762 27776
rect 19826 27712 19834 27776
rect 19514 26688 19834 27712
rect 19514 26624 19522 26688
rect 19586 26624 19602 26688
rect 19666 26624 19682 26688
rect 19746 26624 19762 26688
rect 19826 26624 19834 26688
rect 19514 26094 19834 26624
rect 19514 25858 19556 26094
rect 19792 25858 19834 26094
rect 19514 25600 19834 25858
rect 19514 25536 19522 25600
rect 19586 25536 19602 25600
rect 19666 25536 19682 25600
rect 19746 25536 19762 25600
rect 19826 25536 19834 25600
rect 19514 24512 19834 25536
rect 19514 24448 19522 24512
rect 19586 24448 19602 24512
rect 19666 24448 19682 24512
rect 19746 24448 19762 24512
rect 19826 24448 19834 24512
rect 19514 23424 19834 24448
rect 19514 23360 19522 23424
rect 19586 23360 19602 23424
rect 19666 23360 19682 23424
rect 19746 23360 19762 23424
rect 19826 23360 19834 23424
rect 19514 22336 19834 23360
rect 19514 22272 19522 22336
rect 19586 22272 19602 22336
rect 19666 22272 19682 22336
rect 19746 22272 19762 22336
rect 19826 22272 19834 22336
rect 19514 21248 19834 22272
rect 19514 21184 19522 21248
rect 19586 21184 19602 21248
rect 19666 21184 19682 21248
rect 19746 21184 19762 21248
rect 19826 21184 19834 21248
rect 19514 20160 19834 21184
rect 19514 20096 19522 20160
rect 19586 20096 19602 20160
rect 19666 20096 19682 20160
rect 19746 20096 19762 20160
rect 19826 20096 19834 20160
rect 19514 19294 19834 20096
rect 19514 19072 19556 19294
rect 19792 19072 19834 19294
rect 19514 19008 19522 19072
rect 19586 19008 19602 19058
rect 19666 19008 19682 19058
rect 19746 19008 19762 19058
rect 19826 19008 19834 19072
rect 19514 17984 19834 19008
rect 19514 17920 19522 17984
rect 19586 17920 19602 17984
rect 19666 17920 19682 17984
rect 19746 17920 19762 17984
rect 19826 17920 19834 17984
rect 19514 16896 19834 17920
rect 19514 16832 19522 16896
rect 19586 16832 19602 16896
rect 19666 16832 19682 16896
rect 19746 16832 19762 16896
rect 19826 16832 19834 16896
rect 19514 15808 19834 16832
rect 19514 15744 19522 15808
rect 19586 15744 19602 15808
rect 19666 15744 19682 15808
rect 19746 15744 19762 15808
rect 19826 15744 19834 15808
rect 19514 14720 19834 15744
rect 19514 14656 19522 14720
rect 19586 14656 19602 14720
rect 19666 14656 19682 14720
rect 19746 14656 19762 14720
rect 19826 14656 19834 14720
rect 19514 13632 19834 14656
rect 19514 13568 19522 13632
rect 19586 13568 19602 13632
rect 19666 13568 19682 13632
rect 19746 13568 19762 13632
rect 19826 13568 19834 13632
rect 19514 12544 19834 13568
rect 19514 12480 19522 12544
rect 19586 12494 19602 12544
rect 19666 12494 19682 12544
rect 19746 12494 19762 12544
rect 19826 12480 19834 12544
rect 19514 12258 19556 12480
rect 19792 12258 19834 12480
rect 19514 11456 19834 12258
rect 19514 11392 19522 11456
rect 19586 11392 19602 11456
rect 19666 11392 19682 11456
rect 19746 11392 19762 11456
rect 19826 11392 19834 11456
rect 19514 10368 19834 11392
rect 19514 10304 19522 10368
rect 19586 10304 19602 10368
rect 19666 10304 19682 10368
rect 19746 10304 19762 10368
rect 19826 10304 19834 10368
rect 19514 9280 19834 10304
rect 19514 9216 19522 9280
rect 19586 9216 19602 9280
rect 19666 9216 19682 9280
rect 19746 9216 19762 9280
rect 19826 9216 19834 9280
rect 19514 8192 19834 9216
rect 19514 8128 19522 8192
rect 19586 8128 19602 8192
rect 19666 8128 19682 8192
rect 19746 8128 19762 8192
rect 19826 8128 19834 8192
rect 19514 7104 19834 8128
rect 19514 7040 19522 7104
rect 19586 7040 19602 7104
rect 19666 7040 19682 7104
rect 19746 7040 19762 7104
rect 19826 7040 19834 7104
rect 19514 6016 19834 7040
rect 19514 5952 19522 6016
rect 19586 5952 19602 6016
rect 19666 5952 19682 6016
rect 19746 5952 19762 6016
rect 19826 5952 19834 6016
rect 19514 5694 19834 5952
rect 19514 5458 19556 5694
rect 19792 5458 19834 5694
rect 19514 4928 19834 5458
rect 19514 4864 19522 4928
rect 19586 4864 19602 4928
rect 19666 4864 19682 4928
rect 19746 4864 19762 4928
rect 19826 4864 19834 4928
rect 19514 3840 19834 4864
rect 19514 3776 19522 3840
rect 19586 3776 19602 3840
rect 19666 3776 19682 3840
rect 19746 3776 19762 3840
rect 19826 3776 19834 3840
rect 19514 2752 19834 3776
rect 19514 2688 19522 2752
rect 19586 2688 19602 2752
rect 19666 2688 19682 2752
rect 19746 2688 19762 2752
rect 19826 2688 19834 2752
rect 19514 2128 19834 2688
rect 20174 29408 20494 29424
rect 20174 29344 20182 29408
rect 20246 29344 20262 29408
rect 20326 29344 20342 29408
rect 20406 29344 20422 29408
rect 20486 29344 20494 29408
rect 20174 28320 20494 29344
rect 20174 28256 20182 28320
rect 20246 28256 20262 28320
rect 20326 28256 20342 28320
rect 20406 28256 20422 28320
rect 20486 28256 20494 28320
rect 20174 27232 20494 28256
rect 20174 27168 20182 27232
rect 20246 27168 20262 27232
rect 20326 27168 20342 27232
rect 20406 27168 20422 27232
rect 20486 27168 20494 27232
rect 20174 26754 20494 27168
rect 20174 26518 20216 26754
rect 20452 26518 20494 26754
rect 20174 26144 20494 26518
rect 20174 26080 20182 26144
rect 20246 26080 20262 26144
rect 20326 26080 20342 26144
rect 20406 26080 20422 26144
rect 20486 26080 20494 26144
rect 20174 25056 20494 26080
rect 20174 24992 20182 25056
rect 20246 24992 20262 25056
rect 20326 24992 20342 25056
rect 20406 24992 20422 25056
rect 20486 24992 20494 25056
rect 20174 23968 20494 24992
rect 20174 23904 20182 23968
rect 20246 23904 20262 23968
rect 20326 23904 20342 23968
rect 20406 23904 20422 23968
rect 20486 23904 20494 23968
rect 20174 22880 20494 23904
rect 20174 22816 20182 22880
rect 20246 22816 20262 22880
rect 20326 22816 20342 22880
rect 20406 22816 20422 22880
rect 20486 22816 20494 22880
rect 20174 21792 20494 22816
rect 20174 21728 20182 21792
rect 20246 21728 20262 21792
rect 20326 21728 20342 21792
rect 20406 21728 20422 21792
rect 20486 21728 20494 21792
rect 20174 20704 20494 21728
rect 20174 20640 20182 20704
rect 20246 20640 20262 20704
rect 20326 20640 20342 20704
rect 20406 20640 20422 20704
rect 20486 20640 20494 20704
rect 20174 19954 20494 20640
rect 20174 19718 20216 19954
rect 20452 19718 20494 19954
rect 20174 19616 20494 19718
rect 20174 19552 20182 19616
rect 20246 19552 20262 19616
rect 20326 19552 20342 19616
rect 20406 19552 20422 19616
rect 20486 19552 20494 19616
rect 20174 18528 20494 19552
rect 20174 18464 20182 18528
rect 20246 18464 20262 18528
rect 20326 18464 20342 18528
rect 20406 18464 20422 18528
rect 20486 18464 20494 18528
rect 20174 17440 20494 18464
rect 20174 17376 20182 17440
rect 20246 17376 20262 17440
rect 20326 17376 20342 17440
rect 20406 17376 20422 17440
rect 20486 17376 20494 17440
rect 20174 16352 20494 17376
rect 20174 16288 20182 16352
rect 20246 16288 20262 16352
rect 20326 16288 20342 16352
rect 20406 16288 20422 16352
rect 20486 16288 20494 16352
rect 20174 15264 20494 16288
rect 20174 15200 20182 15264
rect 20246 15200 20262 15264
rect 20326 15200 20342 15264
rect 20406 15200 20422 15264
rect 20486 15200 20494 15264
rect 20174 14176 20494 15200
rect 20174 14112 20182 14176
rect 20246 14112 20262 14176
rect 20326 14112 20342 14176
rect 20406 14112 20422 14176
rect 20486 14112 20494 14176
rect 20174 13154 20494 14112
rect 20174 13088 20216 13154
rect 20452 13088 20494 13154
rect 20174 13024 20182 13088
rect 20486 13024 20494 13088
rect 20174 12918 20216 13024
rect 20452 12918 20494 13024
rect 20174 12000 20494 12918
rect 20174 11936 20182 12000
rect 20246 11936 20262 12000
rect 20326 11936 20342 12000
rect 20406 11936 20422 12000
rect 20486 11936 20494 12000
rect 20174 10912 20494 11936
rect 20174 10848 20182 10912
rect 20246 10848 20262 10912
rect 20326 10848 20342 10912
rect 20406 10848 20422 10912
rect 20486 10848 20494 10912
rect 20174 9824 20494 10848
rect 20174 9760 20182 9824
rect 20246 9760 20262 9824
rect 20326 9760 20342 9824
rect 20406 9760 20422 9824
rect 20486 9760 20494 9824
rect 20174 8736 20494 9760
rect 20174 8672 20182 8736
rect 20246 8672 20262 8736
rect 20326 8672 20342 8736
rect 20406 8672 20422 8736
rect 20486 8672 20494 8736
rect 20174 7648 20494 8672
rect 20174 7584 20182 7648
rect 20246 7584 20262 7648
rect 20326 7584 20342 7648
rect 20406 7584 20422 7648
rect 20486 7584 20494 7648
rect 20174 6560 20494 7584
rect 20174 6496 20182 6560
rect 20246 6496 20262 6560
rect 20326 6496 20342 6560
rect 20406 6496 20422 6560
rect 20486 6496 20494 6560
rect 20174 6354 20494 6496
rect 20174 6118 20216 6354
rect 20452 6118 20494 6354
rect 20174 5472 20494 6118
rect 20174 5408 20182 5472
rect 20246 5408 20262 5472
rect 20326 5408 20342 5472
rect 20406 5408 20422 5472
rect 20486 5408 20494 5472
rect 20174 4384 20494 5408
rect 20174 4320 20182 4384
rect 20246 4320 20262 4384
rect 20326 4320 20342 4384
rect 20406 4320 20422 4384
rect 20486 4320 20494 4384
rect 20174 3296 20494 4320
rect 20174 3232 20182 3296
rect 20246 3232 20262 3296
rect 20326 3232 20342 3296
rect 20406 3232 20422 3296
rect 20486 3232 20494 3296
rect 20174 2208 20494 3232
rect 20174 2144 20182 2208
rect 20246 2144 20262 2208
rect 20326 2144 20342 2208
rect 20406 2144 20422 2208
rect 20486 2144 20494 2208
rect 20174 2128 20494 2144
rect 26942 28864 27262 29424
rect 26942 28800 26950 28864
rect 27014 28800 27030 28864
rect 27094 28800 27110 28864
rect 27174 28800 27190 28864
rect 27254 28800 27262 28864
rect 26942 27776 27262 28800
rect 26942 27712 26950 27776
rect 27014 27712 27030 27776
rect 27094 27712 27110 27776
rect 27174 27712 27190 27776
rect 27254 27712 27262 27776
rect 26942 26688 27262 27712
rect 26942 26624 26950 26688
rect 27014 26624 27030 26688
rect 27094 26624 27110 26688
rect 27174 26624 27190 26688
rect 27254 26624 27262 26688
rect 26942 26094 27262 26624
rect 26942 25858 26984 26094
rect 27220 25858 27262 26094
rect 26942 25600 27262 25858
rect 26942 25536 26950 25600
rect 27014 25536 27030 25600
rect 27094 25536 27110 25600
rect 27174 25536 27190 25600
rect 27254 25536 27262 25600
rect 26942 24512 27262 25536
rect 26942 24448 26950 24512
rect 27014 24448 27030 24512
rect 27094 24448 27110 24512
rect 27174 24448 27190 24512
rect 27254 24448 27262 24512
rect 26942 23424 27262 24448
rect 26942 23360 26950 23424
rect 27014 23360 27030 23424
rect 27094 23360 27110 23424
rect 27174 23360 27190 23424
rect 27254 23360 27262 23424
rect 26942 22336 27262 23360
rect 26942 22272 26950 22336
rect 27014 22272 27030 22336
rect 27094 22272 27110 22336
rect 27174 22272 27190 22336
rect 27254 22272 27262 22336
rect 26942 21248 27262 22272
rect 26942 21184 26950 21248
rect 27014 21184 27030 21248
rect 27094 21184 27110 21248
rect 27174 21184 27190 21248
rect 27254 21184 27262 21248
rect 26942 20160 27262 21184
rect 26942 20096 26950 20160
rect 27014 20096 27030 20160
rect 27094 20096 27110 20160
rect 27174 20096 27190 20160
rect 27254 20096 27262 20160
rect 26942 19294 27262 20096
rect 26942 19072 26984 19294
rect 27220 19072 27262 19294
rect 26942 19008 26950 19072
rect 27014 19008 27030 19058
rect 27094 19008 27110 19058
rect 27174 19008 27190 19058
rect 27254 19008 27262 19072
rect 26942 17984 27262 19008
rect 26942 17920 26950 17984
rect 27014 17920 27030 17984
rect 27094 17920 27110 17984
rect 27174 17920 27190 17984
rect 27254 17920 27262 17984
rect 26942 16896 27262 17920
rect 26942 16832 26950 16896
rect 27014 16832 27030 16896
rect 27094 16832 27110 16896
rect 27174 16832 27190 16896
rect 27254 16832 27262 16896
rect 26942 15808 27262 16832
rect 26942 15744 26950 15808
rect 27014 15744 27030 15808
rect 27094 15744 27110 15808
rect 27174 15744 27190 15808
rect 27254 15744 27262 15808
rect 26942 14720 27262 15744
rect 26942 14656 26950 14720
rect 27014 14656 27030 14720
rect 27094 14656 27110 14720
rect 27174 14656 27190 14720
rect 27254 14656 27262 14720
rect 26942 13632 27262 14656
rect 26942 13568 26950 13632
rect 27014 13568 27030 13632
rect 27094 13568 27110 13632
rect 27174 13568 27190 13632
rect 27254 13568 27262 13632
rect 26942 12544 27262 13568
rect 26942 12480 26950 12544
rect 27014 12494 27030 12544
rect 27094 12494 27110 12544
rect 27174 12494 27190 12544
rect 27254 12480 27262 12544
rect 26942 12258 26984 12480
rect 27220 12258 27262 12480
rect 26942 11456 27262 12258
rect 26942 11392 26950 11456
rect 27014 11392 27030 11456
rect 27094 11392 27110 11456
rect 27174 11392 27190 11456
rect 27254 11392 27262 11456
rect 26942 10368 27262 11392
rect 26942 10304 26950 10368
rect 27014 10304 27030 10368
rect 27094 10304 27110 10368
rect 27174 10304 27190 10368
rect 27254 10304 27262 10368
rect 26942 9280 27262 10304
rect 26942 9216 26950 9280
rect 27014 9216 27030 9280
rect 27094 9216 27110 9280
rect 27174 9216 27190 9280
rect 27254 9216 27262 9280
rect 26942 8192 27262 9216
rect 26942 8128 26950 8192
rect 27014 8128 27030 8192
rect 27094 8128 27110 8192
rect 27174 8128 27190 8192
rect 27254 8128 27262 8192
rect 26942 7104 27262 8128
rect 26942 7040 26950 7104
rect 27014 7040 27030 7104
rect 27094 7040 27110 7104
rect 27174 7040 27190 7104
rect 27254 7040 27262 7104
rect 26942 6016 27262 7040
rect 26942 5952 26950 6016
rect 27014 5952 27030 6016
rect 27094 5952 27110 6016
rect 27174 5952 27190 6016
rect 27254 5952 27262 6016
rect 26942 5694 27262 5952
rect 26942 5458 26984 5694
rect 27220 5458 27262 5694
rect 26942 4928 27262 5458
rect 26942 4864 26950 4928
rect 27014 4864 27030 4928
rect 27094 4864 27110 4928
rect 27174 4864 27190 4928
rect 27254 4864 27262 4928
rect 26942 3840 27262 4864
rect 26942 3776 26950 3840
rect 27014 3776 27030 3840
rect 27094 3776 27110 3840
rect 27174 3776 27190 3840
rect 27254 3776 27262 3840
rect 26942 2752 27262 3776
rect 26942 2688 26950 2752
rect 27014 2688 27030 2752
rect 27094 2688 27110 2752
rect 27174 2688 27190 2752
rect 27254 2688 27262 2752
rect 26942 2128 27262 2688
rect 27602 29408 27922 29424
rect 27602 29344 27610 29408
rect 27674 29344 27690 29408
rect 27754 29344 27770 29408
rect 27834 29344 27850 29408
rect 27914 29344 27922 29408
rect 27602 28320 27922 29344
rect 27602 28256 27610 28320
rect 27674 28256 27690 28320
rect 27754 28256 27770 28320
rect 27834 28256 27850 28320
rect 27914 28256 27922 28320
rect 27602 27232 27922 28256
rect 27602 27168 27610 27232
rect 27674 27168 27690 27232
rect 27754 27168 27770 27232
rect 27834 27168 27850 27232
rect 27914 27168 27922 27232
rect 27602 26754 27922 27168
rect 27602 26518 27644 26754
rect 27880 26518 27922 26754
rect 27602 26144 27922 26518
rect 27602 26080 27610 26144
rect 27674 26080 27690 26144
rect 27754 26080 27770 26144
rect 27834 26080 27850 26144
rect 27914 26080 27922 26144
rect 27602 25056 27922 26080
rect 27602 24992 27610 25056
rect 27674 24992 27690 25056
rect 27754 24992 27770 25056
rect 27834 24992 27850 25056
rect 27914 24992 27922 25056
rect 27602 23968 27922 24992
rect 27602 23904 27610 23968
rect 27674 23904 27690 23968
rect 27754 23904 27770 23968
rect 27834 23904 27850 23968
rect 27914 23904 27922 23968
rect 27602 22880 27922 23904
rect 27602 22816 27610 22880
rect 27674 22816 27690 22880
rect 27754 22816 27770 22880
rect 27834 22816 27850 22880
rect 27914 22816 27922 22880
rect 27602 21792 27922 22816
rect 27602 21728 27610 21792
rect 27674 21728 27690 21792
rect 27754 21728 27770 21792
rect 27834 21728 27850 21792
rect 27914 21728 27922 21792
rect 27602 20704 27922 21728
rect 27602 20640 27610 20704
rect 27674 20640 27690 20704
rect 27754 20640 27770 20704
rect 27834 20640 27850 20704
rect 27914 20640 27922 20704
rect 27602 19954 27922 20640
rect 27602 19718 27644 19954
rect 27880 19718 27922 19954
rect 27602 19616 27922 19718
rect 27602 19552 27610 19616
rect 27674 19552 27690 19616
rect 27754 19552 27770 19616
rect 27834 19552 27850 19616
rect 27914 19552 27922 19616
rect 27602 18528 27922 19552
rect 27602 18464 27610 18528
rect 27674 18464 27690 18528
rect 27754 18464 27770 18528
rect 27834 18464 27850 18528
rect 27914 18464 27922 18528
rect 27602 17440 27922 18464
rect 27602 17376 27610 17440
rect 27674 17376 27690 17440
rect 27754 17376 27770 17440
rect 27834 17376 27850 17440
rect 27914 17376 27922 17440
rect 27602 16352 27922 17376
rect 27602 16288 27610 16352
rect 27674 16288 27690 16352
rect 27754 16288 27770 16352
rect 27834 16288 27850 16352
rect 27914 16288 27922 16352
rect 27602 15264 27922 16288
rect 27602 15200 27610 15264
rect 27674 15200 27690 15264
rect 27754 15200 27770 15264
rect 27834 15200 27850 15264
rect 27914 15200 27922 15264
rect 27602 14176 27922 15200
rect 27602 14112 27610 14176
rect 27674 14112 27690 14176
rect 27754 14112 27770 14176
rect 27834 14112 27850 14176
rect 27914 14112 27922 14176
rect 27602 13154 27922 14112
rect 27602 13088 27644 13154
rect 27880 13088 27922 13154
rect 27602 13024 27610 13088
rect 27914 13024 27922 13088
rect 27602 12918 27644 13024
rect 27880 12918 27922 13024
rect 27602 12000 27922 12918
rect 27602 11936 27610 12000
rect 27674 11936 27690 12000
rect 27754 11936 27770 12000
rect 27834 11936 27850 12000
rect 27914 11936 27922 12000
rect 27602 10912 27922 11936
rect 27602 10848 27610 10912
rect 27674 10848 27690 10912
rect 27754 10848 27770 10912
rect 27834 10848 27850 10912
rect 27914 10848 27922 10912
rect 27602 9824 27922 10848
rect 27602 9760 27610 9824
rect 27674 9760 27690 9824
rect 27754 9760 27770 9824
rect 27834 9760 27850 9824
rect 27914 9760 27922 9824
rect 27602 8736 27922 9760
rect 27602 8672 27610 8736
rect 27674 8672 27690 8736
rect 27754 8672 27770 8736
rect 27834 8672 27850 8736
rect 27914 8672 27922 8736
rect 27602 7648 27922 8672
rect 27602 7584 27610 7648
rect 27674 7584 27690 7648
rect 27754 7584 27770 7648
rect 27834 7584 27850 7648
rect 27914 7584 27922 7648
rect 27602 6560 27922 7584
rect 27602 6496 27610 6560
rect 27674 6496 27690 6560
rect 27754 6496 27770 6560
rect 27834 6496 27850 6560
rect 27914 6496 27922 6560
rect 27602 6354 27922 6496
rect 27602 6118 27644 6354
rect 27880 6118 27922 6354
rect 27602 5472 27922 6118
rect 27602 5408 27610 5472
rect 27674 5408 27690 5472
rect 27754 5408 27770 5472
rect 27834 5408 27850 5472
rect 27914 5408 27922 5472
rect 27602 4384 27922 5408
rect 27602 4320 27610 4384
rect 27674 4320 27690 4384
rect 27754 4320 27770 4384
rect 27834 4320 27850 4384
rect 27914 4320 27922 4384
rect 27602 3296 27922 4320
rect 27602 3232 27610 3296
rect 27674 3232 27690 3296
rect 27754 3232 27770 3296
rect 27834 3232 27850 3296
rect 27914 3232 27922 3296
rect 27602 2208 27922 3232
rect 27602 2144 27610 2208
rect 27674 2144 27690 2208
rect 27754 2144 27770 2208
rect 27834 2144 27850 2208
rect 27914 2144 27922 2208
rect 27602 2128 27922 2144
<< via4 >>
rect 4700 25858 4936 26094
rect 4700 19072 4936 19294
rect 4700 19058 4730 19072
rect 4730 19058 4746 19072
rect 4746 19058 4810 19072
rect 4810 19058 4826 19072
rect 4826 19058 4890 19072
rect 4890 19058 4906 19072
rect 4906 19058 4936 19072
rect 4700 12480 4730 12494
rect 4730 12480 4746 12494
rect 4746 12480 4810 12494
rect 4810 12480 4826 12494
rect 4826 12480 4890 12494
rect 4890 12480 4906 12494
rect 4906 12480 4936 12494
rect 4700 12258 4936 12480
rect 4700 5458 4936 5694
rect 5360 26518 5596 26754
rect 5360 19718 5596 19954
rect 5360 13088 5596 13154
rect 5360 13024 5390 13088
rect 5390 13024 5406 13088
rect 5406 13024 5470 13088
rect 5470 13024 5486 13088
rect 5486 13024 5550 13088
rect 5550 13024 5566 13088
rect 5566 13024 5596 13088
rect 5360 12918 5596 13024
rect 5360 6118 5596 6354
rect 12128 25858 12364 26094
rect 12128 19072 12364 19294
rect 12128 19058 12158 19072
rect 12158 19058 12174 19072
rect 12174 19058 12238 19072
rect 12238 19058 12254 19072
rect 12254 19058 12318 19072
rect 12318 19058 12334 19072
rect 12334 19058 12364 19072
rect 12128 12480 12158 12494
rect 12158 12480 12174 12494
rect 12174 12480 12238 12494
rect 12238 12480 12254 12494
rect 12254 12480 12318 12494
rect 12318 12480 12334 12494
rect 12334 12480 12364 12494
rect 12128 12258 12364 12480
rect 12128 5458 12364 5694
rect 12788 26518 13024 26754
rect 12788 19718 13024 19954
rect 12788 13088 13024 13154
rect 12788 13024 12818 13088
rect 12818 13024 12834 13088
rect 12834 13024 12898 13088
rect 12898 13024 12914 13088
rect 12914 13024 12978 13088
rect 12978 13024 12994 13088
rect 12994 13024 13024 13088
rect 12788 12918 13024 13024
rect 12788 6118 13024 6354
rect 19556 25858 19792 26094
rect 19556 19072 19792 19294
rect 19556 19058 19586 19072
rect 19586 19058 19602 19072
rect 19602 19058 19666 19072
rect 19666 19058 19682 19072
rect 19682 19058 19746 19072
rect 19746 19058 19762 19072
rect 19762 19058 19792 19072
rect 19556 12480 19586 12494
rect 19586 12480 19602 12494
rect 19602 12480 19666 12494
rect 19666 12480 19682 12494
rect 19682 12480 19746 12494
rect 19746 12480 19762 12494
rect 19762 12480 19792 12494
rect 19556 12258 19792 12480
rect 19556 5458 19792 5694
rect 20216 26518 20452 26754
rect 20216 19718 20452 19954
rect 20216 13088 20452 13154
rect 20216 13024 20246 13088
rect 20246 13024 20262 13088
rect 20262 13024 20326 13088
rect 20326 13024 20342 13088
rect 20342 13024 20406 13088
rect 20406 13024 20422 13088
rect 20422 13024 20452 13088
rect 20216 12918 20452 13024
rect 20216 6118 20452 6354
rect 26984 25858 27220 26094
rect 26984 19072 27220 19294
rect 26984 19058 27014 19072
rect 27014 19058 27030 19072
rect 27030 19058 27094 19072
rect 27094 19058 27110 19072
rect 27110 19058 27174 19072
rect 27174 19058 27190 19072
rect 27190 19058 27220 19072
rect 26984 12480 27014 12494
rect 27014 12480 27030 12494
rect 27030 12480 27094 12494
rect 27094 12480 27110 12494
rect 27110 12480 27174 12494
rect 27174 12480 27190 12494
rect 27190 12480 27220 12494
rect 26984 12258 27220 12480
rect 26984 5458 27220 5694
rect 27644 26518 27880 26754
rect 27644 19718 27880 19954
rect 27644 13088 27880 13154
rect 27644 13024 27674 13088
rect 27674 13024 27690 13088
rect 27690 13024 27754 13088
rect 27754 13024 27770 13088
rect 27770 13024 27834 13088
rect 27834 13024 27850 13088
rect 27850 13024 27880 13088
rect 27644 12918 27880 13024
rect 27644 6118 27880 6354
<< metal5 >>
rect 1056 26754 30868 26796
rect 1056 26518 5360 26754
rect 5596 26518 12788 26754
rect 13024 26518 20216 26754
rect 20452 26518 27644 26754
rect 27880 26518 30868 26754
rect 1056 26476 30868 26518
rect 1056 26094 30868 26136
rect 1056 25858 4700 26094
rect 4936 25858 12128 26094
rect 12364 25858 19556 26094
rect 19792 25858 26984 26094
rect 27220 25858 30868 26094
rect 1056 25816 30868 25858
rect 1056 19954 30868 19996
rect 1056 19718 5360 19954
rect 5596 19718 12788 19954
rect 13024 19718 20216 19954
rect 20452 19718 27644 19954
rect 27880 19718 30868 19954
rect 1056 19676 30868 19718
rect 1056 19294 30868 19336
rect 1056 19058 4700 19294
rect 4936 19058 12128 19294
rect 12364 19058 19556 19294
rect 19792 19058 26984 19294
rect 27220 19058 30868 19294
rect 1056 19016 30868 19058
rect 1056 13154 30868 13196
rect 1056 12918 5360 13154
rect 5596 12918 12788 13154
rect 13024 12918 20216 13154
rect 20452 12918 27644 13154
rect 27880 12918 30868 13154
rect 1056 12876 30868 12918
rect 1056 12494 30868 12536
rect 1056 12258 4700 12494
rect 4936 12258 12128 12494
rect 12364 12258 19556 12494
rect 19792 12258 26984 12494
rect 27220 12258 30868 12494
rect 1056 12216 30868 12258
rect 1056 6354 30868 6396
rect 1056 6118 5360 6354
rect 5596 6118 12788 6354
rect 13024 6118 20216 6354
rect 20452 6118 27644 6354
rect 27880 6118 30868 6354
rect 1056 6076 30868 6118
rect 1056 5694 30868 5736
rect 1056 5458 4700 5694
rect 4936 5458 12128 5694
rect 12364 5458 19556 5694
rect 19792 5458 26984 5694
rect 27220 5458 30868 5694
rect 1056 5416 30868 5458
use sky130_fd_sc_hd__inv_2  _0542_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16008 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0543_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16192 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15456 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0545_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 13616 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0546_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0547_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0548_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15272 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14720 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0550_
timestamp 1698431365
transform 1 0 14352 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0551_
timestamp 1698431365
transform -1 0 13984 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0552_
timestamp 1698431365
transform 1 0 17388 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0553_
timestamp 1698431365
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0554_
timestamp 1698431365
transform 1 0 24840 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0555_
timestamp 1698431365
transform 1 0 23644 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0556_
timestamp 1698431365
transform -1 0 25300 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0557_
timestamp 1698431365
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0558_
timestamp 1698431365
transform 1 0 21896 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0559_
timestamp 1698431365
transform 1 0 21528 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0560_
timestamp 1698431365
transform 1 0 19412 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1698431365
transform -1 0 19136 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 21344 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0563_
timestamp 1698431365
transform 1 0 17848 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0564_
timestamp 1698431365
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0565_
timestamp 1698431365
transform 1 0 15824 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0566_
timestamp 1698431365
transform -1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_2  _0567_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14904 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_2  _0568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14352 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 15364 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0571_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14168 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21344 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0573_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 23092 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0574_
timestamp 1698431365
transform -1 0 23828 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0575_
timestamp 1698431365
transform 1 0 21252 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0576_
timestamp 1698431365
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0577_
timestamp 1698431365
transform 1 0 17756 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0578_
timestamp 1698431365
transform 1 0 18584 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0579_
timestamp 1698431365
transform -1 0 15088 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0580_
timestamp 1698431365
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0581_
timestamp 1698431365
transform 1 0 7544 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0582_
timestamp 1698431365
transform -1 0 8832 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0583_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 7176 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0584_
timestamp 1698431365
transform -1 0 6164 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0585_
timestamp 1698431365
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0586_
timestamp 1698431365
transform 1 0 12236 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12604 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _0588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13156 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0589_
timestamp 1698431365
transform -1 0 11408 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0590_
timestamp 1698431365
transform -1 0 26404 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0591_
timestamp 1698431365
transform 1 0 23552 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0592_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 23644 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0593_
timestamp 1698431365
transform 1 0 19688 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0594_
timestamp 1698431365
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 20332 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 21436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0598_
timestamp 1698431365
transform 1 0 23276 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0599_
timestamp 1698431365
transform 1 0 23368 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0600_
timestamp 1698431365
transform 1 0 24288 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0601_
timestamp 1698431365
transform 1 0 24012 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0602_
timestamp 1698431365
transform -1 0 24932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0603_
timestamp 1698431365
transform 1 0 24564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0604_
timestamp 1698431365
transform 1 0 25668 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0605_
timestamp 1698431365
transform -1 0 27048 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0606_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 24932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1698431365
transform 1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0608_
timestamp 1698431365
transform 1 0 23092 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0609_
timestamp 1698431365
transform -1 0 24196 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0610_
timestamp 1698431365
transform 1 0 23828 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0611_
timestamp 1698431365
transform -1 0 24932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0612_
timestamp 1698431365
transform -1 0 24104 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0613_
timestamp 1698431365
transform 1 0 24472 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0614_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0615_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14996 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0616_
timestamp 1698431365
transform 1 0 17940 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0617_
timestamp 1698431365
transform -1 0 18768 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0618_
timestamp 1698431365
transform -1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0619_
timestamp 1698431365
transform 1 0 21252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0620_
timestamp 1698431365
transform -1 0 22356 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0621_
timestamp 1698431365
transform -1 0 22172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0622_
timestamp 1698431365
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0623_
timestamp 1698431365
transform -1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19504 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0625_
timestamp 1698431365
transform 1 0 16744 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0626_
timestamp 1698431365
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0627_
timestamp 1698431365
transform 1 0 16744 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0628_
timestamp 1698431365
transform 1 0 17296 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0629_
timestamp 1698431365
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0630_
timestamp 1698431365
transform -1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0631_
timestamp 1698431365
transform -1 0 18860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0632_
timestamp 1698431365
transform 1 0 18768 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0633_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 17664 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0634_
timestamp 1698431365
transform 1 0 19872 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0635_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 20332 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1698431365
transform 1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0637_
timestamp 1698431365
transform 1 0 20792 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1698431365
transform -1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0639_
timestamp 1698431365
transform 1 0 16928 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0640_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17020 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1698431365
transform -1 0 19136 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0643_
timestamp 1698431365
transform -1 0 17480 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1698431365
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1698431365
transform -1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0646_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14168 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0647_
timestamp 1698431365
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16836 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0649_
timestamp 1698431365
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0650_
timestamp 1698431365
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0651_
timestamp 1698431365
transform -1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0652_
timestamp 1698431365
transform 1 0 7728 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0653_
timestamp 1698431365
transform 1 0 8280 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0654_
timestamp 1698431365
transform 1 0 8832 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0655_
timestamp 1698431365
transform 1 0 7820 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0656_
timestamp 1698431365
transform 1 0 7820 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0657_
timestamp 1698431365
transform 1 0 7268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 1698431365
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1698431365
transform 1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0660_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 7360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0661_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 6348 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0662_
timestamp 1698431365
transform 1 0 7360 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0663_
timestamp 1698431365
transform 1 0 8188 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0664_
timestamp 1698431365
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0665_
timestamp 1698431365
transform 1 0 11040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0666_
timestamp 1698431365
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0667_
timestamp 1698431365
transform 1 0 13156 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0668_
timestamp 1698431365
transform 1 0 13156 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0669_
timestamp 1698431365
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1698431365
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0671_
timestamp 1698431365
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0672_
timestamp 1698431365
transform -1 0 13800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0673_
timestamp 1698431365
transform -1 0 13248 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1698431365
transform -1 0 13064 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0675_
timestamp 1698431365
transform -1 0 11040 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0676_
timestamp 1698431365
transform -1 0 10304 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0677_
timestamp 1698431365
transform 1 0 9292 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0678_
timestamp 1698431365
transform -1 0 12052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0679_
timestamp 1698431365
transform -1 0 11316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0680_
timestamp 1698431365
transform 1 0 10028 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0681_
timestamp 1698431365
transform -1 0 7360 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0682_
timestamp 1698431365
transform 1 0 8280 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0683_
timestamp 1698431365
transform 1 0 8280 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0684_
timestamp 1698431365
transform -1 0 9476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0685_
timestamp 1698431365
transform 1 0 6808 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1698431365
transform 1 0 5336 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1698431365
transform 1 0 5336 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0688_
timestamp 1698431365
transform 1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0689_
timestamp 1698431365
transform 1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0690_
timestamp 1698431365
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0691_
timestamp 1698431365
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1698431365
transform 1 0 7176 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0693_
timestamp 1698431365
transform 1 0 6532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0694_
timestamp 1698431365
transform 1 0 7084 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1698431365
transform 1 0 7636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 9752 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0697_
timestamp 1698431365
transform 1 0 6992 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0698_
timestamp 1698431365
transform 1 0 7820 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1698431365
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0700_
timestamp 1698431365
transform 1 0 7452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0701_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _0702_
timestamp 1698431365
transform -1 0 12052 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0703_
timestamp 1698431365
transform -1 0 9752 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0704_
timestamp 1698431365
transform 1 0 8648 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0705_
timestamp 1698431365
transform -1 0 10672 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0706_
timestamp 1698431365
transform -1 0 9844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0707_
timestamp 1698431365
transform 1 0 9844 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0708_
timestamp 1698431365
transform 1 0 13156 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0709_
timestamp 1698431365
transform -1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0710_
timestamp 1698431365
transform 1 0 10488 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0711_
timestamp 1698431365
transform 1 0 12604 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0712_
timestamp 1698431365
transform -1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0713_
timestamp 1698431365
transform -1 0 15088 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0714_
timestamp 1698431365
transform 1 0 13248 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0715_
timestamp 1698431365
transform 1 0 13064 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21068 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0717_
timestamp 1698431365
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0718_
timestamp 1698431365
transform 1 0 12052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0719_
timestamp 1698431365
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0720_
timestamp 1698431365
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0721_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 13616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0722_
timestamp 1698431365
transform -1 0 13340 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1698431365
transform -1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0724_
timestamp 1698431365
transform -1 0 11132 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1698431365
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0726_
timestamp 1698431365
transform -1 0 13984 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 18860 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _0728_
timestamp 1698431365
transform -1 0 19136 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0729_
timestamp 1698431365
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0730_
timestamp 1698431365
transform 1 0 11316 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0731_
timestamp 1698431365
transform 1 0 20884 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 10488 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0733_
timestamp 1698431365
transform 1 0 9384 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1698431365
transform 1 0 10672 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _0735_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11960 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _0736_
timestamp 1698431365
transform -1 0 11868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0737_
timestamp 1698431365
transform 1 0 9292 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1698431365
transform 1 0 8924 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 1698431365
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0740_
timestamp 1698431365
transform -1 0 8648 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _0741_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9292 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0742_
timestamp 1698431365
transform 1 0 10856 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1698431365
transform -1 0 11408 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0744_
timestamp 1698431365
transform 1 0 10488 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0745_
timestamp 1698431365
transform 1 0 9292 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0746_
timestamp 1698431365
transform -1 0 8832 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1698431365
transform -1 0 8372 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1698431365
transform -1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0749_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 7728 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0750_
timestamp 1698431365
transform 1 0 7360 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0751_
timestamp 1698431365
transform 1 0 8188 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0752_
timestamp 1698431365
transform -1 0 8188 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1698431365
transform -1 0 6164 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1698431365
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0755_
timestamp 1698431365
transform 1 0 6256 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0756_
timestamp 1698431365
transform -1 0 6808 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0757_
timestamp 1698431365
transform -1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0758_
timestamp 1698431365
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0759_
timestamp 1698431365
transform 1 0 4416 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0760_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 4968 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1698431365
transform 1 0 4232 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0762_
timestamp 1698431365
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0763_
timestamp 1698431365
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0764_
timestamp 1698431365
transform 1 0 14260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0765_
timestamp 1698431365
transform 1 0 7636 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0766_
timestamp 1698431365
transform 1 0 6900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1698431365
transform -1 0 6440 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0768_
timestamp 1698431365
transform -1 0 6164 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0769_
timestamp 1698431365
transform 1 0 5336 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0770_
timestamp 1698431365
transform 1 0 4692 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1698431365
transform -1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0772_
timestamp 1698431365
transform -1 0 8372 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0773_
timestamp 1698431365
transform -1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0774_
timestamp 1698431365
transform 1 0 5336 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0775_
timestamp 1698431365
transform 1 0 4600 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1698431365
transform -1 0 5796 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 1698431365
transform 1 0 6440 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0778_
timestamp 1698431365
transform 1 0 5980 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0779_
timestamp 1698431365
transform -1 0 10488 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _0780_
timestamp 1698431365
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0781_
timestamp 1698431365
transform 1 0 9384 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0782_
timestamp 1698431365
transform -1 0 7360 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0783_
timestamp 1698431365
transform -1 0 7636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0784_
timestamp 1698431365
transform 1 0 7636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0785_
timestamp 1698431365
transform 1 0 8280 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0786_
timestamp 1698431365
transform 1 0 7176 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0787_
timestamp 1698431365
transform 1 0 6440 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0788_
timestamp 1698431365
transform -1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0789_
timestamp 1698431365
transform 1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0790_
timestamp 1698431365
transform 1 0 6164 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0791_
timestamp 1698431365
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1698431365
transform 1 0 4784 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 1698431365
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0794_
timestamp 1698431365
transform -1 0 7912 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0795_
timestamp 1698431365
transform -1 0 8464 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 1698431365
transform 1 0 8464 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0797_
timestamp 1698431365
transform -1 0 9476 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0798_
timestamp 1698431365
transform -1 0 8188 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0799_
timestamp 1698431365
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0800_
timestamp 1698431365
transform 1 0 5520 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0801_
timestamp 1698431365
transform -1 0 6072 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1698431365
transform -1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0803_
timestamp 1698431365
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o311ai_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 10028 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1698431365
transform 1 0 8740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0806_
timestamp 1698431365
transform 1 0 7084 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1698431365
transform -1 0 13708 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0808_
timestamp 1698431365
transform -1 0 10672 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0809_
timestamp 1698431365
transform -1 0 10948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_2  _0810_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 12696 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0811_
timestamp 1698431365
transform -1 0 11684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0812_
timestamp 1698431365
transform -1 0 11408 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0813_
timestamp 1698431365
transform 1 0 9108 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1698431365
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 1698431365
transform -1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1698431365
transform -1 0 13984 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0817_
timestamp 1698431365
transform -1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0818_
timestamp 1698431365
transform -1 0 12604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0819_
timestamp 1698431365
transform 1 0 12512 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1698431365
transform 1 0 12144 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0821_
timestamp 1698431365
transform 1 0 11868 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0822_
timestamp 1698431365
transform -1 0 13984 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1698431365
transform -1 0 13708 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0824_
timestamp 1698431365
transform -1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0825_
timestamp 1698431365
transform 1 0 11776 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0826_
timestamp 1698431365
transform 1 0 12788 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0827_
timestamp 1698431365
transform 1 0 12420 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0828_
timestamp 1698431365
transform 1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0829_
timestamp 1698431365
transform -1 0 10948 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0830_
timestamp 1698431365
transform 1 0 10028 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0831_
timestamp 1698431365
transform -1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0832_
timestamp 1698431365
transform 1 0 13248 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0833_
timestamp 1698431365
transform 1 0 10304 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0834_
timestamp 1698431365
transform 1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1698431365
transform 1 0 20056 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0836_
timestamp 1698431365
transform 1 0 17020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0837_
timestamp 1698431365
transform 1 0 16836 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0838_
timestamp 1698431365
transform 1 0 16008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1698431365
transform 1 0 14720 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0840_
timestamp 1698431365
transform -1 0 16284 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1698431365
transform -1 0 15180 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0842_
timestamp 1698431365
transform -1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 16008 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1698431365
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0845_
timestamp 1698431365
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0846_
timestamp 1698431365
transform -1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0847_
timestamp 1698431365
transform -1 0 17020 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 1698431365
transform 1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0849_
timestamp 1698431365
transform 1 0 15364 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0850_
timestamp 1698431365
transform -1 0 16836 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1698431365
transform 1 0 15640 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0852_
timestamp 1698431365
transform -1 0 15640 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0853_
timestamp 1698431365
transform 1 0 18124 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0854_
timestamp 1698431365
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1698431365
transform 1 0 17664 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1698431365
transform 1 0 18400 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0857_
timestamp 1698431365
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1698431365
transform -1 0 19136 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1698431365
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0860_
timestamp 1698431365
transform -1 0 18032 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0861_
timestamp 1698431365
transform 1 0 15824 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0862_
timestamp 1698431365
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0863_
timestamp 1698431365
transform 1 0 19412 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0864_
timestamp 1698431365
transform 1 0 16100 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0865_
timestamp 1698431365
transform -1 0 20424 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0866_
timestamp 1698431365
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16836 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0868_
timestamp 1698431365
transform 1 0 15456 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1698431365
transform -1 0 18676 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0870_
timestamp 1698431365
transform -1 0 17572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0871_
timestamp 1698431365
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0872_
timestamp 1698431365
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0873_
timestamp 1698431365
transform -1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0874_
timestamp 1698431365
transform -1 0 19688 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 1698431365
transform -1 0 18952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1698431365
transform 1 0 17848 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0878_
timestamp 1698431365
transform 1 0 17296 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 22172 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0880_
timestamp 1698431365
transform -1 0 22264 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0881_
timestamp 1698431365
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1698431365
transform -1 0 20332 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0883_
timestamp 1698431365
transform -1 0 21068 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0884_
timestamp 1698431365
transform 1 0 20516 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0885_
timestamp 1698431365
transform 1 0 19872 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0886_
timestamp 1698431365
transform -1 0 20148 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0887_
timestamp 1698431365
transform 1 0 19688 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0888_
timestamp 1698431365
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0889_
timestamp 1698431365
transform 1 0 21252 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0890_
timestamp 1698431365
transform 1 0 19688 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0891_
timestamp 1698431365
transform -1 0 20608 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0892_
timestamp 1698431365
transform 1 0 21436 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1698431365
transform -1 0 23000 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1698431365
transform 1 0 22356 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0895_
timestamp 1698431365
transform -1 0 23368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1698431365
transform 1 0 24472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1698431365
transform 1 0 24932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0898_
timestamp 1698431365
transform -1 0 25392 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0899_
timestamp 1698431365
transform 1 0 24564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0900_
timestamp 1698431365
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0901_
timestamp 1698431365
transform 1 0 24840 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0902_
timestamp 1698431365
transform -1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0903_
timestamp 1698431365
transform 1 0 23276 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 25760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0905_
timestamp 1698431365
transform 1 0 24932 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1698431365
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0907_
timestamp 1698431365
transform -1 0 23276 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0908_
timestamp 1698431365
transform 1 0 25300 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1698431365
transform -1 0 22908 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1698431365
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0911_
timestamp 1698431365
transform 1 0 25668 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0912_
timestamp 1698431365
transform -1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0913_
timestamp 1698431365
transform -1 0 25760 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0914_
timestamp 1698431365
transform 1 0 21896 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0915_
timestamp 1698431365
transform 1 0 20884 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1698431365
transform 1 0 20516 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1698431365
transform -1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0918_
timestamp 1698431365
transform -1 0 25668 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0919_
timestamp 1698431365
transform 1 0 21988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1698431365
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1698431365
transform -1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1698431365
transform -1 0 26496 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0923_
timestamp 1698431365
transform 1 0 24656 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _0924_
timestamp 1698431365
transform -1 0 25852 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0925_
timestamp 1698431365
transform 1 0 24564 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1698431365
transform 1 0 20700 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0927_
timestamp 1698431365
transform 1 0 22356 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1698431365
transform 1 0 23368 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0929_
timestamp 1698431365
transform -1 0 24196 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0930_
timestamp 1698431365
transform 1 0 24748 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0931_
timestamp 1698431365
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0932_
timestamp 1698431365
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0933_
timestamp 1698431365
transform 1 0 22172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 1698431365
transform -1 0 22632 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1698431365
transform 1 0 22356 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0936_
timestamp 1698431365
transform -1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0937_
timestamp 1698431365
transform 1 0 19872 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1698431365
transform 1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0939_
timestamp 1698431365
transform 1 0 20332 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0940_
timestamp 1698431365
transform 1 0 19504 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0941_
timestamp 1698431365
transform -1 0 17020 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1698431365
transform -1 0 17572 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0943_
timestamp 1698431365
transform 1 0 17112 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0944_
timestamp 1698431365
transform -1 0 17112 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0945_
timestamp 1698431365
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1698431365
transform -1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0947_
timestamp 1698431365
transform 1 0 18400 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1698431365
transform 1 0 25668 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0949_
timestamp 1698431365
transform -1 0 23092 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1698431365
transform 1 0 19504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1698431365
transform 1 0 19964 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 19780 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1698431365
transform -1 0 21620 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0954_
timestamp 1698431365
transform -1 0 21896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21896 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0956_
timestamp 1698431365
transform 1 0 26128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0957_
timestamp 1698431365
transform -1 0 26588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0958_
timestamp 1698431365
transform 1 0 25208 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0959_
timestamp 1698431365
transform -1 0 26496 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0960_
timestamp 1698431365
transform 1 0 17756 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1698431365
transform -1 0 24656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1698431365
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0963_
timestamp 1698431365
transform 1 0 21988 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _0964_
timestamp 1698431365
transform 1 0 16468 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 23092 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0966_
timestamp 1698431365
transform 1 0 17664 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0967_
timestamp 1698431365
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0968_
timestamp 1698431365
transform 1 0 15180 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0969_
timestamp 1698431365
transform 1 0 17020 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _0970_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 16928 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0971_
timestamp 1698431365
transform 1 0 23736 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0972_
timestamp 1698431365
transform 1 0 23092 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 23276 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 24564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0975_
timestamp 1698431365
transform -1 0 18216 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0976_
timestamp 1698431365
transform 1 0 24932 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1698431365
transform -1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0978_
timestamp 1698431365
transform -1 0 18952 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1698431365
transform -1 0 26956 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0980_
timestamp 1698431365
transform -1 0 26680 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0981_
timestamp 1698431365
transform 1 0 24380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0982_
timestamp 1698431365
transform 1 0 23736 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0983_
timestamp 1698431365
transform 1 0 24380 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0984_
timestamp 1698431365
transform 1 0 23644 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0985_
timestamp 1698431365
transform 1 0 23828 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0986_
timestamp 1698431365
transform -1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0987_
timestamp 1698431365
transform -1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0988_
timestamp 1698431365
transform 1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0989_
timestamp 1698431365
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1698431365
transform -1 0 23092 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0991_
timestamp 1698431365
transform 1 0 21252 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0992_
timestamp 1698431365
transform 1 0 22080 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_1  _0993_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 21252 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _0994_
timestamp 1698431365
transform -1 0 22264 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0995_
timestamp 1698431365
transform 1 0 22632 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0996_
timestamp 1698431365
transform -1 0 22632 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1698431365
transform -1 0 21620 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1698431365
transform -1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0999_
timestamp 1698431365
transform 1 0 19780 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1000_
timestamp 1698431365
transform 1 0 20424 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1001_
timestamp 1698431365
transform 1 0 20056 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1002_
timestamp 1698431365
transform 1 0 20516 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1003_
timestamp 1698431365
transform 1 0 20516 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1698431365
transform -1 0 20884 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1698431365
transform -1 0 19964 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1006_
timestamp 1698431365
transform -1 0 18860 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1007_
timestamp 1698431365
transform -1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1008_
timestamp 1698431365
transform 1 0 18492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1009_
timestamp 1698431365
transform -1 0 19504 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1698431365
transform -1 0 18400 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1011_
timestamp 1698431365
transform 1 0 18492 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1698431365
transform 1 0 5244 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1698431365
transform 1 0 6716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1014_
timestamp 1698431365
transform 1 0 14812 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1015_
timestamp 1698431365
transform 1 0 14444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1698431365
transform -1 0 15732 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1017_
timestamp 1698431365
transform 1 0 14260 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1018_
timestamp 1698431365
transform 1 0 14444 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1698431365
transform 1 0 14996 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1698431365
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1021_
timestamp 1698431365
transform -1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1022_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1023_
timestamp 1698431365
transform -1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1024_
timestamp 1698431365
transform 1 0 15824 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1025_
timestamp 1698431365
transform 1 0 18492 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1026_
timestamp 1698431365
transform 1 0 19964 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1027_
timestamp 1698431365
transform 1 0 22356 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1028_
timestamp 1698431365
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1029_
timestamp 1698431365
transform 1 0 24472 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1030_
timestamp 1698431365
transform 1 0 12236 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1698431365
transform 1 0 12788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1032_
timestamp 1698431365
transform 1 0 13708 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1033_
timestamp 1698431365
transform 1 0 25116 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1698431365
transform 1 0 19320 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1698431365
transform 1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1698431365
transform 1 0 22816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1698431365
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1698431365
transform 1 0 25944 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1698431365
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1698431365
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1698431365
transform -1 0 24196 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1698431365
transform 1 0 27416 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1698431365
transform -1 0 23920 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1044_
timestamp 1698431365
transform 1 0 14996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1698431365
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp 1698431365
transform 1 0 26128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp 1698431365
transform -1 0 24472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp 1698431365
transform -1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1698431365
transform 1 0 19964 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1698431365
transform 1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1698431365
transform -1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1698431365
transform -1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1698431365
transform -1 0 20516 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1698431365
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1055_
timestamp 1698431365
transform -1 0 13616 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1698431365
transform 1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1698431365
transform 1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1698431365
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1698431365
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1698431365
transform -1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1698431365
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1698431365
transform -1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1698431365
transform -1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1698431365
transform -1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1698431365
transform -1 0 4416 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1066_
timestamp 1698431365
transform -1 0 14260 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1698431365
transform -1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1698431365
transform -1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1698431365
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1698431365
transform -1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1698431365
transform -1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1698431365
transform -1 0 11408 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1698431365
transform 1 0 12236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1698431365
transform -1 0 19044 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1698431365
transform 1 0 19412 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1698431365
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1698431365
transform 1 0 25668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1698431365
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1698431365
transform 1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1698431365
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1698431365
transform -1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1082_
timestamp 1698431365
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1083_
timestamp 1698431365
transform 1 0 9660 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1698431365
transform -1 0 17388 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1698431365
transform -1 0 15916 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1698431365
transform -1 0 14352 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1698431365
transform -1 0 14352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1088_
timestamp 1698431365
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1698431365
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1698431365
transform 1 0 6164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 1698431365
transform 1 0 4784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1092_
timestamp 1698431365
transform 1 0 5336 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1093_
timestamp 1698431365
transform -1 0 7728 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1698431365
transform 1 0 6348 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11500 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 12420 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _1097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 18400 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 20148 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 24196 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1100_
timestamp 1698431365
transform 1 0 24380 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1101_
timestamp 1698431365
transform 1 0 25116 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1102_
timestamp 1698431365
transform 1 0 17112 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1103_
timestamp 1698431365
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1104_
timestamp 1698431365
transform 1 0 22080 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1105_
timestamp 1698431365
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1106_
timestamp 1698431365
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1107_
timestamp 1698431365
transform 1 0 19964 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1108_
timestamp 1698431365
transform 1 0 25392 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1109_
timestamp 1698431365
transform 1 0 23092 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1110_
timestamp 1698431365
transform 1 0 21804 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1111_
timestamp 1698431365
transform 1 0 19044 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1112_
timestamp 1698431365
transform 1 0 16652 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1113_
timestamp 1698431365
transform 1 0 14076 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1114_
timestamp 1698431365
transform -1 0 16100 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1115_
timestamp 1698431365
transform 1 0 19136 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1116_
timestamp 1698431365
transform 1 0 16652 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1117_
timestamp 1698431365
transform 1 0 11776 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1118_
timestamp 1698431365
transform 1 0 9476 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1119_
timestamp 1698431365
transform 1 0 11500 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1120_
timestamp 1698431365
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1121_
timestamp 1698431365
transform 1 0 8556 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1122_
timestamp 1698431365
transform -1 0 6532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1123_
timestamp 1698431365
transform -1 0 5428 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1124_
timestamp 1698431365
transform 1 0 2944 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1125_
timestamp 1698431365
transform -1 0 5060 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1126_
timestamp 1698431365
transform -1 0 5060 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1127_
timestamp 1698431365
transform -1 0 5152 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1128_
timestamp 1698431365
transform 1 0 3312 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1129_
timestamp 1698431365
transform 1 0 6348 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1130_
timestamp 1698431365
transform 1 0 9016 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1131_
timestamp 1698431365
transform 1 0 8280 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1132_
timestamp 1698431365
transform -1 0 12052 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1133_
timestamp 1698431365
transform 1 0 11500 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1134_
timestamp 1698431365
transform 1 0 16928 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1698431365
transform 1 0 19228 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1698431365
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1698431365
transform 1 0 24564 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1698431365
transform 1 0 23000 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1139_
timestamp 1698431365
transform 1 0 16652 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1140_
timestamp 1698431365
transform 1 0 14260 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1141_
timestamp 1698431365
transform 1 0 14444 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1698431365
transform 1 0 10212 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1143_
timestamp 1698431365
transform 1 0 15916 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1144_
timestamp 1698431365
transform 1 0 14444 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1145_
timestamp 1698431365
transform 1 0 12328 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1698431365
transform 1 0 12144 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1698431365
transform 1 0 10028 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1698431365
transform 1 0 8188 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1698431365
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1698431365
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1698431365
transform 1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1698431365
transform 1 0 6716 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clock
timestamp 1698431365
transform -1 0 10672 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clock
timestamp 1698431365
transform -1 0 10764 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clock
timestamp 1698431365
transform 1 0 19228 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clock
timestamp 1698431365
transform 1 0 19596 0 -1 19584
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1698431365
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1698431365
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1698431365
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1698431365
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1698431365
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1698431365
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 1698431365
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1698431365
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1698431365
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118
timestamp 1698431365
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_126
timestamp 1698431365
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_133
timestamp 1698431365
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1698431365
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1698431365
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_154
timestamp 1698431365
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_161
timestamp 1698431365
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1698431365
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_175
timestamp 1698431365
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_182
timestamp 1698431365
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_189
timestamp 1698431365
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 1698431365
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1698431365
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_209
timestamp 1698431365
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_217
timestamp 1698431365
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1698431365
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1698431365
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1698431365
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1698431365
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1698431365
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1698431365
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1698431365
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1698431365
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1698431365
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1698431365
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_309
timestamp 1698431365
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_317
timestamp 1698431365
transform 1 0 30268 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1698431365
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1698431365
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1698431365
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1698431365
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1698431365
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1698431365
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1698431365
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1698431365
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1698431365
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1698431365
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1698431365
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1698431365
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1698431365
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1698431365
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1698431365
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1698431365
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1698431365
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1698431365
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1698431365
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1698431365
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1698431365
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1698431365
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1698431365
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1698431365
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1698431365
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1698431365
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1698431365
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1698431365
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1698431365
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1698431365
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1698431365
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1698431365
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_317
timestamp 1698431365
transform 1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1698431365
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1698431365
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1698431365
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1698431365
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1698431365
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1698431365
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1698431365
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1698431365
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1698431365
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1698431365
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1698431365
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1698431365
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1698431365
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1698431365
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1698431365
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1698431365
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1698431365
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1698431365
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1698431365
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1698431365
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1698431365
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1698431365
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1698431365
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1698431365
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1698431365
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1698431365
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1698431365
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1698431365
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1698431365
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1698431365
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1698431365
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1698431365
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1698431365
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_309
timestamp 1698431365
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_317
timestamp 1698431365
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1698431365
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1698431365
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1698431365
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1698431365
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1698431365
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1698431365
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1698431365
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1698431365
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1698431365
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1698431365
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1698431365
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1698431365
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1698431365
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1698431365
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1698431365
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1698431365
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1698431365
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1698431365
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1698431365
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1698431365
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1698431365
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1698431365
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1698431365
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1698431365
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1698431365
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1698431365
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1698431365
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1698431365
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1698431365
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1698431365
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1698431365
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1698431365
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_317
timestamp 1698431365
transform 1 0 30268 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1698431365
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1698431365
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1698431365
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1698431365
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1698431365
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1698431365
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1698431365
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1698431365
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1698431365
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1698431365
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1698431365
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1698431365
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1698431365
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1698431365
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1698431365
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1698431365
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1698431365
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1698431365
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1698431365
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1698431365
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1698431365
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1698431365
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1698431365
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1698431365
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1698431365
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1698431365
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1698431365
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1698431365
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1698431365
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1698431365
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1698431365
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1698431365
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_309
timestamp 1698431365
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_317
timestamp 1698431365
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1698431365
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1698431365
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1698431365
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1698431365
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1698431365
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1698431365
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1698431365
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1698431365
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1698431365
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1698431365
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1698431365
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1698431365
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1698431365
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1698431365
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1698431365
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1698431365
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1698431365
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1698431365
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1698431365
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1698431365
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1698431365
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1698431365
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1698431365
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1698431365
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1698431365
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1698431365
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1698431365
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1698431365
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1698431365
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1698431365
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1698431365
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1698431365
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_317
timestamp 1698431365
transform 1 0 30268 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1698431365
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1698431365
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1698431365
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1698431365
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1698431365
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1698431365
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1698431365
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1698431365
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1698431365
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1698431365
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1698431365
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1698431365
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1698431365
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1698431365
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1698431365
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1698431365
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1698431365
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1698431365
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1698431365
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1698431365
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1698431365
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1698431365
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1698431365
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1698431365
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1698431365
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1698431365
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1698431365
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1698431365
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1698431365
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1698431365
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1698431365
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1698431365
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_309
timestamp 1698431365
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_317
timestamp 1698431365
transform 1 0 30268 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1698431365
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1698431365
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1698431365
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1698431365
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1698431365
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1698431365
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1698431365
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1698431365
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1698431365
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1698431365
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1698431365
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1698431365
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1698431365
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1698431365
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1698431365
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1698431365
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1698431365
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1698431365
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1698431365
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1698431365
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1698431365
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1698431365
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1698431365
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1698431365
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1698431365
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1698431365
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1698431365
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1698431365
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1698431365
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1698431365
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1698431365
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1698431365
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_317
timestamp 1698431365
transform 1 0 30268 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1698431365
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1698431365
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1698431365
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1698431365
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1698431365
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1698431365
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1698431365
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1698431365
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1698431365
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_94
timestamp 1698431365
transform 1 0 9752 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_106
timestamp 1698431365
transform 1 0 10856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_114
timestamp 1698431365
transform 1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_120
timestamp 1698431365
transform 1 0 12144 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp 1698431365
transform 1 0 13248 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1698431365
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1698431365
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_165
timestamp 1698431365
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_173
timestamp 1698431365
transform 1 0 17020 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1698431365
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1698431365
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1698431365
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1698431365
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_208
timestamp 1698431365
transform 1 0 20240 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_220
timestamp 1698431365
transform 1 0 21344 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_232
timestamp 1698431365
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_244
timestamp 1698431365
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1698431365
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1698431365
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1698431365
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1698431365
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1698431365
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1698431365
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_309
timestamp 1698431365
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_317
timestamp 1698431365
transform 1 0 30268 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 1698431365
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1698431365
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1698431365
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_42
timestamp 1698431365
transform 1 0 4968 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_48
timestamp 1698431365
transform 1 0 5520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1698431365
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1698431365
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1698431365
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_77
timestamp 1698431365
transform 1 0 8188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1698431365
transform 1 0 10672 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_136
timestamp 1698431365
transform 1 0 13616 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_148
timestamp 1698431365
transform 1 0 14720 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_160
timestamp 1698431365
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_189
timestamp 1698431365
transform 1 0 18492 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_215
timestamp 1698431365
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1698431365
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1698431365
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1698431365
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1698431365
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1698431365
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1698431365
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1698431365
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1698431365
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1698431365
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_317
timestamp 1698431365
transform 1 0 30268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_7
timestamp 1698431365
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 1698431365
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1698431365
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1698431365
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1698431365
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_62
timestamp 1698431365
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_66
timestamp 1698431365
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1698431365
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1698431365
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1698431365
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1698431365
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_109
timestamp 1698431365
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_117
timestamp 1698431365
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_129
timestamp 1698431365
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1698431365
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1698431365
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1698431365
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_165
timestamp 1698431365
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_173
timestamp 1698431365
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_190
timestamp 1698431365
transform 1 0 18584 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1698431365
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1698431365
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_209
timestamp 1698431365
transform 1 0 20332 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_240
timestamp 1698431365
transform 1 0 23184 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1698431365
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1698431365
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1698431365
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1698431365
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1698431365
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1698431365
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_309
timestamp 1698431365
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_317
timestamp 1698431365
transform 1 0 30268 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1698431365
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1698431365
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1698431365
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_42
timestamp 1698431365
transform 1 0 4968 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_50
timestamp 1698431365
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_80
timestamp 1698431365
transform 1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_91
timestamp 1698431365
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_95
timestamp 1698431365
transform 1 0 9844 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_102
timestamp 1698431365
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1698431365
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_125
timestamp 1698431365
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_138
timestamp 1698431365
transform 1 0 13800 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_150
timestamp 1698431365
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1698431365
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1698431365
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1698431365
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_182
timestamp 1698431365
transform 1 0 17848 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_194
timestamp 1698431365
transform 1 0 18952 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1698431365
transform 1 0 19688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_207
timestamp 1698431365
transform 1 0 20148 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_213
timestamp 1698431365
transform 1 0 20700 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_245
timestamp 1698431365
transform 1 0 23644 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_254
timestamp 1698431365
transform 1 0 24472 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_266
timestamp 1698431365
transform 1 0 25576 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1698431365
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1698431365
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_305
timestamp 1698431365
transform 1 0 29164 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_313
timestamp 1698431365
transform 1 0 29900 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1698431365
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1698431365
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1698431365
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1698431365
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_40
timestamp 1698431365
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_48
timestamp 1698431365
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_56
timestamp 1698431365
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_68
timestamp 1698431365
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1698431365
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_111
timestamp 1698431365
transform 1 0 11316 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_115
timestamp 1698431365
transform 1 0 11684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_123
timestamp 1698431365
transform 1 0 12420 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1698431365
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_149
timestamp 1698431365
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_158
timestamp 1698431365
transform 1 0 15640 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_179
timestamp 1698431365
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_202
timestamp 1698431365
transform 1 0 19688 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_215
timestamp 1698431365
transform 1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_229
timestamp 1698431365
transform 1 0 22172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_234
timestamp 1698431365
transform 1 0 22632 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_240
timestamp 1698431365
transform 1 0 23184 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_248
timestamp 1698431365
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1698431365
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1698431365
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1698431365
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1698431365
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1698431365
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1698431365
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_309
timestamp 1698431365
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_315
timestamp 1698431365
transform 1 0 30084 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1698431365
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1698431365
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1698431365
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_62
timestamp 1698431365
transform 1 0 6808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_74
timestamp 1698431365
transform 1 0 7912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_86
timestamp 1698431365
transform 1 0 9016 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_98
timestamp 1698431365
transform 1 0 10120 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_102
timestamp 1698431365
transform 1 0 10488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1698431365
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1698431365
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_130
timestamp 1698431365
transform 1 0 13064 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_142
timestamp 1698431365
transform 1 0 14168 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_148
timestamp 1698431365
transform 1 0 14720 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_159
timestamp 1698431365
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1698431365
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1698431365
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_182
timestamp 1698431365
transform 1 0 17848 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_194
timestamp 1698431365
transform 1 0 18952 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_210
timestamp 1698431365
transform 1 0 20424 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1698431365
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_267
timestamp 1698431365
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1698431365
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1698431365
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1698431365
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_317
timestamp 1698431365
transform 1 0 30268 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_7
timestamp 1698431365
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1698431365
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1698431365
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1698431365
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_37
timestamp 1698431365
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_55
timestamp 1698431365
transform 1 0 6164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_61
timestamp 1698431365
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1698431365
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1698431365
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_89
timestamp 1698431365
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1698431365
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_109
timestamp 1698431365
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_113
timestamp 1698431365
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_125
timestamp 1698431365
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1698431365
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_179
timestamp 1698431365
transform 1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1698431365
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1698431365
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1698431365
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1698431365
transform 1 0 19596 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_217
timestamp 1698431365
transform 1 0 21068 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_228
timestamp 1698431365
transform 1 0 22080 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_236
timestamp 1698431365
transform 1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1698431365
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_253
timestamp 1698431365
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_269
timestamp 1698431365
transform 1 0 25852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_281
timestamp 1698431365
transform 1 0 26956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_293
timestamp 1698431365
transform 1 0 28060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_305
timestamp 1698431365
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_309
timestamp 1698431365
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_7
timestamp 1698431365
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_19
timestamp 1698431365
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_31
timestamp 1698431365
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_43
timestamp 1698431365
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1698431365
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1698431365
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_64
timestamp 1698431365
transform 1 0 6992 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_76
timestamp 1698431365
transform 1 0 8096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_82
timestamp 1698431365
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1698431365
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_126
timestamp 1698431365
transform 1 0 12696 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_130
timestamp 1698431365
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_143
timestamp 1698431365
transform 1 0 14260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_151
timestamp 1698431365
transform 1 0 14996 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1698431365
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1698431365
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1698431365
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_194
timestamp 1698431365
transform 1 0 18952 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_202
timestamp 1698431365
transform 1 0 19688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_209
timestamp 1698431365
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_230
timestamp 1698431365
transform 1 0 22264 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_247
timestamp 1698431365
transform 1 0 23828 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_261
timestamp 1698431365
transform 1 0 25116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_269
timestamp 1698431365
transform 1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1698431365
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1698431365
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1698431365
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_7
timestamp 1698431365
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_19
timestamp 1698431365
transform 1 0 2852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_29
timestamp 1698431365
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_35
timestamp 1698431365
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_47
timestamp 1698431365
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_51
timestamp 1698431365
transform 1 0 5796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_58
timestamp 1698431365
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_68
timestamp 1698431365
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_72
timestamp 1698431365
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1698431365
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1698431365
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1698431365
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_109
timestamp 1698431365
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_119
timestamp 1698431365
transform 1 0 12052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1698431365
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_170
timestamp 1698431365
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_182
timestamp 1698431365
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_186
timestamp 1698431365
transform 1 0 18216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_191
timestamp 1698431365
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1698431365
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1698431365
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_209
timestamp 1698431365
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_224
timestamp 1698431365
transform 1 0 21712 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_232
timestamp 1698431365
transform 1 0 22448 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_238
timestamp 1698431365
transform 1 0 23000 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_242
timestamp 1698431365
transform 1 0 23368 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 1698431365
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_253
timestamp 1698431365
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_257
timestamp 1698431365
transform 1 0 24748 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_263
timestamp 1698431365
transform 1 0 25300 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_284
timestamp 1698431365
transform 1 0 27232 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_296
timestamp 1698431365
transform 1 0 28336 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1698431365
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_6
timestamp 1698431365
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_18
timestamp 1698431365
transform 1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1698431365
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_64
timestamp 1698431365
transform 1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_87
timestamp 1698431365
transform 1 0 9108 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_100
timestamp 1698431365
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1698431365
transform 1 0 11776 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_128
timestamp 1698431365
transform 1 0 12880 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1698431365
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_149
timestamp 1698431365
transform 1 0 14812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_153
timestamp 1698431365
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_162
timestamp 1698431365
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1698431365
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_211
timestamp 1698431365
transform 1 0 20516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1698431365
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_241
timestamp 1698431365
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_262
timestamp 1698431365
transform 1 0 25208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_270
timestamp 1698431365
transform 1 0 25944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_289
timestamp 1698431365
transform 1 0 27692 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_301
timestamp 1698431365
transform 1 0 28796 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_313
timestamp 1698431365
transform 1 0 29900 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1698431365
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1698431365
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1698431365
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1698431365
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1698431365
transform 1 0 4876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_49
timestamp 1698431365
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_54
timestamp 1698431365
transform 1 0 6072 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_60
timestamp 1698431365
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1698431365
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1698431365
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_107
timestamp 1698431365
transform 1 0 10948 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_114
timestamp 1698431365
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_126
timestamp 1698431365
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_150
timestamp 1698431365
transform 1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_158
timestamp 1698431365
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_167
timestamp 1698431365
transform 1 0 16468 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_184
timestamp 1698431365
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_200
timestamp 1698431365
transform 1 0 19504 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_222
timestamp 1698431365
transform 1 0 21528 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_234
timestamp 1698431365
transform 1 0 22632 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 23368 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1698431365
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_253
timestamp 1698431365
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_268
timestamp 1698431365
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_280
timestamp 1698431365
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_292
timestamp 1698431365
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_304
timestamp 1698431365
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_309
timestamp 1698431365
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_317
timestamp 1698431365
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_7
timestamp 1698431365
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_19
timestamp 1698431365
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1698431365
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1698431365
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_73
timestamp 1698431365
transform 1 0 7820 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_77
timestamp 1698431365
transform 1 0 8188 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_89
timestamp 1698431365
transform 1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 1698431365
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_119
timestamp 1698431365
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_131
timestamp 1698431365
transform 1 0 13156 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_143
timestamp 1698431365
transform 1 0 14260 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_153
timestamp 1698431365
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1698431365
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1698431365
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_179
timestamp 1698431365
transform 1 0 17572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_191
timestamp 1698431365
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_200
timestamp 1698431365
transform 1 0 19504 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_208
timestamp 1698431365
transform 1 0 20240 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_214
timestamp 1698431365
transform 1 0 20792 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_225
timestamp 1698431365
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_237
timestamp 1698431365
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_241
timestamp 1698431365
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_248
timestamp 1698431365
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_264
timestamp 1698431365
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1698431365
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1698431365
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_305
timestamp 1698431365
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_313
timestamp 1698431365
transform 1 0 29900 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_7
timestamp 1698431365
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1698431365
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1698431365
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1698431365
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_36
timestamp 1698431365
transform 1 0 4416 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_42
timestamp 1698431365
transform 1 0 4968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_51
timestamp 1698431365
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_61
timestamp 1698431365
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_73
timestamp 1698431365
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1698431365
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_91
timestamp 1698431365
transform 1 0 9476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_99
timestamp 1698431365
transform 1 0 10212 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_107
timestamp 1698431365
transform 1 0 10948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_116
timestamp 1698431365
transform 1 0 11776 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_120
timestamp 1698431365
transform 1 0 12144 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1698431365
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1698431365
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_165
timestamp 1698431365
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_173
timestamp 1698431365
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_183
timestamp 1698431365
transform 1 0 17940 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_187
timestamp 1698431365
transform 1 0 18308 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1698431365
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1698431365
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_225
timestamp 1698431365
transform 1 0 21804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_239
timestamp 1698431365
transform 1 0 23092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1698431365
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1698431365
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_259
timestamp 1698431365
transform 1 0 24932 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_268
timestamp 1698431365
transform 1 0 25760 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_280
timestamp 1698431365
transform 1 0 26864 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_292
timestamp 1698431365
transform 1 0 27968 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_304
timestamp 1698431365
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_309
timestamp 1698431365
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_315
timestamp 1698431365
transform 1 0 30084 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 1698431365
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_18
timestamp 1698431365
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_22
timestamp 1698431365
transform 1 0 3128 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_43
timestamp 1698431365
transform 1 0 5060 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_47
timestamp 1698431365
transform 1 0 5428 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1698431365
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1698431365
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1698431365
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_69
timestamp 1698431365
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_73
timestamp 1698431365
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_79
timestamp 1698431365
transform 1 0 8372 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1698431365
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_133
timestamp 1698431365
transform 1 0 13340 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 13892 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_146
timestamp 1698431365
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_153
timestamp 1698431365
transform 1 0 15180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1698431365
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 1698431365
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_178
timestamp 1698431365
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_185
timestamp 1698431365
transform 1 0 18124 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_191
timestamp 1698431365
transform 1 0 18676 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_203
timestamp 1698431365
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_207
timestamp 1698431365
transform 1 0 20148 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_211
timestamp 1698431365
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 1698431365
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_225
timestamp 1698431365
transform 1 0 21804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_231
timestamp 1698431365
transform 1 0 22356 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1698431365
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_249
timestamp 1698431365
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_258
timestamp 1698431365
transform 1 0 24840 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_264
timestamp 1698431365
transform 1 0 25392 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1698431365
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1698431365
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1698431365
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_7
timestamp 1698431365
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_19
timestamp 1698431365
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1698431365
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_29
timestamp 1698431365
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_33
timestamp 1698431365
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_42
timestamp 1698431365
transform 1 0 4968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_58
timestamp 1698431365
transform 1 0 6440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_94
timestamp 1698431365
transform 1 0 9752 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_105
timestamp 1698431365
transform 1 0 10764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_117
timestamp 1698431365
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_124
timestamp 1698431365
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1698431365
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 1698431365
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_149
timestamp 1698431365
transform 1 0 14812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_184
timestamp 1698431365
transform 1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_238
timestamp 1698431365
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1698431365
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_259
timestamp 1698431365
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_272
timestamp 1698431365
transform 1 0 26128 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_284
timestamp 1698431365
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_296
timestamp 1698431365
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1698431365
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1698431365
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1698431365
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1698431365
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_27
timestamp 1698431365
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_35
timestamp 1698431365
transform 1 0 4324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_45
timestamp 1698431365
transform 1 0 5244 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1698431365
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1698431365
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_65
timestamp 1698431365
transform 1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 7728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_76
timestamp 1698431365
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_80
timestamp 1698431365
transform 1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_104
timestamp 1698431365
transform 1 0 10672 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_119
timestamp 1698431365
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_124
timestamp 1698431365
transform 1 0 12512 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1698431365
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_139
timestamp 1698431365
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_145
timestamp 1698431365
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1698431365
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1698431365
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_173
timestamp 1698431365
transform 1 0 17020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_185
timestamp 1698431365
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1698431365
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_234
timestamp 1698431365
transform 1 0 22632 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_246
timestamp 1698431365
transform 1 0 23736 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_255
timestamp 1698431365
transform 1 0 24564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_267
timestamp 1698431365
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1698431365
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1698431365
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1698431365
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_317
timestamp 1698431365
transform 1 0 30268 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_6
timestamp 1698431365
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1698431365
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1698431365
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 4508 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_59
timestamp 1698431365
transform 1 0 6532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_78
timestamp 1698431365
transform 1 0 8280 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1698431365
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_115
timestamp 1698431365
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1698431365
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_148
timestamp 1698431365
transform 1 0 14720 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_154
timestamp 1698431365
transform 1 0 15272 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_158
timestamp 1698431365
transform 1 0 15640 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1698431365
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_189
timestamp 1698431365
transform 1 0 18492 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1698431365
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 1698431365
transform 1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_221
timestamp 1698431365
transform 1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1698431365
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_253
timestamp 1698431365
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_274
timestamp 1698431365
transform 1 0 26312 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_286
timestamp 1698431365
transform 1 0 27416 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_298
timestamp 1698431365
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1698431365
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_309
timestamp 1698431365
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_315
timestamp 1698431365
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_7
timestamp 1698431365
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_19
timestamp 1698431365
transform 1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_23
timestamp 1698431365
transform 1 0 3220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1698431365
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_63
timestamp 1698431365
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_70
timestamp 1698431365
transform 1 0 7544 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_82
timestamp 1698431365
transform 1 0 8648 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_88
timestamp 1698431365
transform 1 0 9200 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_96
timestamp 1698431365
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1698431365
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_119
timestamp 1698431365
transform 1 0 12052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_127
timestamp 1698431365
transform 1 0 12788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_136
timestamp 1698431365
transform 1 0 13616 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_143
timestamp 1698431365
transform 1 0 14260 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_157
timestamp 1698431365
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1698431365
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_196
timestamp 1698431365
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_208
timestamp 1698431365
transform 1 0 20240 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_212
timestamp 1698431365
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_218
timestamp 1698431365
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_225
timestamp 1698431365
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_236
timestamp 1698431365
transform 1 0 22816 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_248
timestamp 1698431365
transform 1 0 23920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_254
timestamp 1698431365
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_260
timestamp 1698431365
transform 1 0 25024 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_268
timestamp 1698431365
transform 1 0 25760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_275
timestamp 1698431365
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1698431365
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1698431365
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_305
timestamp 1698431365
transform 1 0 29164 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_313
timestamp 1698431365
transform 1 0 29900 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_7
timestamp 1698431365
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_19
timestamp 1698431365
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1698431365
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1698431365
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_41
timestamp 1698431365
transform 1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_47
timestamp 1698431365
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_59
timestamp 1698431365
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_71
timestamp 1698431365
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_78
timestamp 1698431365
transform 1 0 8280 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1698431365
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_94
timestamp 1698431365
transform 1 0 9752 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_112
timestamp 1698431365
transform 1 0 11408 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_133
timestamp 1698431365
transform 1 0 13340 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1698431365
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_163
timestamp 1698431365
transform 1 0 16100 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_171
timestamp 1698431365
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_175
timestamp 1698431365
transform 1 0 17204 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 17572 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1698431365
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_207
timestamp 1698431365
transform 1 0 20148 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1698431365
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_253
timestamp 1698431365
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_269
timestamp 1698431365
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_282
timestamp 1698431365
transform 1 0 27048 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_294
timestamp 1698431365
transform 1 0 28152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_306
timestamp 1698431365
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_309
timestamp 1698431365
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_13
timestamp 1698431365
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_25
timestamp 1698431365
transform 1 0 3404 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_33
timestamp 1698431365
transform 1 0 4140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_43
timestamp 1698431365
transform 1 0 5060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_50
timestamp 1698431365
transform 1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_76
timestamp 1698431365
transform 1 0 8096 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_96
timestamp 1698431365
transform 1 0 9936 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1698431365
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_117
timestamp 1698431365
transform 1 0 11868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_136
timestamp 1698431365
transform 1 0 13616 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_143
timestamp 1698431365
transform 1 0 14260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_153
timestamp 1698431365
transform 1 0 15180 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_157
timestamp 1698431365
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_161
timestamp 1698431365
transform 1 0 15916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1698431365
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_173
timestamp 1698431365
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_180
timestamp 1698431365
transform 1 0 17664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_186
timestamp 1698431365
transform 1 0 18216 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1698431365
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1698431365
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_237
timestamp 1698431365
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_243
timestamp 1698431365
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_250
timestamp 1698431365
transform 1 0 24104 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_256
timestamp 1698431365
transform 1 0 24656 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_264
timestamp 1698431365
transform 1 0 25392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1698431365
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1698431365
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_305
timestamp 1698431365
transform 1 0 29164 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_313
timestamp 1698431365
transform 1 0 29900 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1698431365
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1698431365
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1698431365
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1698431365
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1698431365
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_55
timestamp 1698431365
transform 1 0 6164 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_66
timestamp 1698431365
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_70
timestamp 1698431365
transform 1 0 7544 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_74
timestamp 1698431365
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_82
timestamp 1698431365
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1698431365
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 1698431365
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1698431365
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1698431365
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1698431365
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_133
timestamp 1698431365
transform 1 0 13340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1698431365
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_166
timestamp 1698431365
transform 1 0 16376 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1698431365
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_203
timestamp 1698431365
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_210
timestamp 1698431365
transform 1 0 20424 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_222
timestamp 1698431365
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_234
timestamp 1698431365
transform 1 0 22632 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_246
timestamp 1698431365
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_253
timestamp 1698431365
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_257
timestamp 1698431365
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1698431365
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1698431365
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1698431365
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_309
timestamp 1698431365
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_317
timestamp 1698431365
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_7
timestamp 1698431365
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_19
timestamp 1698431365
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_31
timestamp 1698431365
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_43
timestamp 1698431365
transform 1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_52
timestamp 1698431365
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1698431365
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_65
timestamp 1698431365
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_82
timestamp 1698431365
transform 1 0 8648 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_88
timestamp 1698431365
transform 1 0 9200 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_120
timestamp 1698431365
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_137
timestamp 1698431365
transform 1 0 13708 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1698431365
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1698431365
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1698431365
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_173
timestamp 1698431365
transform 1 0 17020 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_179
timestamp 1698431365
transform 1 0 17572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_187
timestamp 1698431365
transform 1 0 18308 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp 1698431365
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1698431365
transform 1 0 19596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1698431365
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_237
timestamp 1698431365
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_245
timestamp 1698431365
transform 1 0 23644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_257
timestamp 1698431365
transform 1 0 24748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_270
timestamp 1698431365
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1698431365
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1698431365
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_305
timestamp 1698431365
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_313
timestamp 1698431365
transform 1 0 29900 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1698431365
transform 1 0 1656 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1698431365
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1698431365
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4048 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_43
timestamp 1698431365
transform 1 0 5060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_52
timestamp 1698431365
transform 1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1698431365
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1698431365
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1698431365
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_85
timestamp 1698431365
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_91
timestamp 1698431365
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1698431365
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_110
timestamp 1698431365
transform 1 0 11224 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_118
timestamp 1698431365
transform 1 0 11960 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_126
timestamp 1698431365
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1698431365
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1698431365
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_152
timestamp 1698431365
transform 1 0 15088 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_160
timestamp 1698431365
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_166
timestamp 1698431365
transform 1 0 16376 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_175
timestamp 1698431365
transform 1 0 17204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_186
timestamp 1698431365
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1698431365
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1698431365
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_208
timestamp 1698431365
transform 1 0 20240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_225
timestamp 1698431365
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1698431365
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_253
timestamp 1698431365
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_281
timestamp 1698431365
transform 1 0 26956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_293
timestamp 1698431365
transform 1 0 28060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_305
timestamp 1698431365
transform 1 0 29164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_309
timestamp 1698431365
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_315
timestamp 1698431365
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_6
timestamp 1698431365
transform 1 0 1656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_18
timestamp 1698431365
transform 1 0 2760 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_47
timestamp 1698431365
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1698431365
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_57
timestamp 1698431365
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1698431365
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_78
timestamp 1698431365
transform 1 0 8280 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_84
timestamp 1698431365
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1698431365
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1698431365
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_121
timestamp 1698431365
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_125
timestamp 1698431365
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_129
timestamp 1698431365
transform 1 0 12972 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_137
timestamp 1698431365
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_141
timestamp 1698431365
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1698431365
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_190
timestamp 1698431365
transform 1 0 18584 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_198
timestamp 1698431365
transform 1 0 19320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_225
timestamp 1698431365
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_235
timestamp 1698431365
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_247
timestamp 1698431365
transform 1 0 23828 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_275
timestamp 1698431365
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1698431365
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1698431365
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_305
timestamp 1698431365
transform 1 0 29164 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1698431365
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1698431365
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1698431365
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1698431365
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1698431365
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_53
timestamp 1698431365
transform 1 0 5980 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_59
timestamp 1698431365
transform 1 0 6532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_63
timestamp 1698431365
transform 1 0 6900 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_78
timestamp 1698431365
transform 1 0 8280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_94
timestamp 1698431365
transform 1 0 9752 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_98
timestamp 1698431365
transform 1 0 10120 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_123
timestamp 1698431365
transform 1 0 12420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1698431365
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_141
timestamp 1698431365
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_154
timestamp 1698431365
transform 1 0 15272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_158
timestamp 1698431365
transform 1 0 15640 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_162
timestamp 1698431365
transform 1 0 16008 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_174
timestamp 1698431365
transform 1 0 17112 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_180
timestamp 1698431365
transform 1 0 17664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_192
timestamp 1698431365
transform 1 0 18768 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_248
timestamp 1698431365
transform 1 0 23920 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1698431365
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1698431365
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1698431365
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1698431365
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1698431365
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1698431365
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_309
timestamp 1698431365
transform 1 0 29532 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_315
timestamp 1698431365
transform 1 0 30084 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1698431365
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1698431365
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1698431365
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1698431365
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1698431365
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1698431365
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_104
timestamp 1698431365
transform 1 0 10672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_108
timestamp 1698431365
transform 1 0 11040 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1698431365
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_132
timestamp 1698431365
transform 1 0 13248 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_144
timestamp 1698431365
transform 1 0 14352 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1698431365
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_180
timestamp 1698431365
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_191
timestamp 1698431365
transform 1 0 18676 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_202
timestamp 1698431365
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_212
timestamp 1698431365
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_225
timestamp 1698431365
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_275
timestamp 1698431365
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1698431365
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1698431365
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1698431365
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_317
timestamp 1698431365
transform 1 0 30268 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1698431365
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1698431365
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1698431365
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_29
timestamp 1698431365
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_58
timestamp 1698431365
transform 1 0 6440 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_70
timestamp 1698431365
transform 1 0 7544 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1698431365
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_94
timestamp 1698431365
transform 1 0 9752 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_106
timestamp 1698431365
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_118
timestamp 1698431365
transform 1 0 11960 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_124
timestamp 1698431365
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_136
timestamp 1698431365
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 1698431365
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_147
timestamp 1698431365
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_151
timestamp 1698431365
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_155
timestamp 1698431365
transform 1 0 15364 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_160
timestamp 1698431365
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1698431365
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_210
timestamp 1698431365
transform 1 0 20424 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_222
timestamp 1698431365
transform 1 0 21528 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_239
timestamp 1698431365
transform 1 0 23092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1698431365
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_268
timestamp 1698431365
transform 1 0 25760 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_281
timestamp 1698431365
transform 1 0 26956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_293
timestamp 1698431365
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1698431365
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1698431365
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_315
timestamp 1698431365
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 1698431365
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 1698431365
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_31
timestamp 1698431365
transform 1 0 3956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_37
timestamp 1698431365
transform 1 0 4508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_49
timestamp 1698431365
transform 1 0 5612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1698431365
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_60
timestamp 1698431365
transform 1 0 6624 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_100
timestamp 1698431365
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1698431365
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1698431365
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1698431365
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_181
timestamp 1698431365
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_196
timestamp 1698431365
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1698431365
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_235
timestamp 1698431365
transform 1 0 22724 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_243
timestamp 1698431365
transform 1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_251
timestamp 1698431365
transform 1 0 24196 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_261
timestamp 1698431365
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_277
timestamp 1698431365
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1698431365
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1698431365
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_305
timestamp 1698431365
transform 1 0 29164 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_7
timestamp 1698431365
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1698431365
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1698431365
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_50
timestamp 1698431365
transform 1 0 5704 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_72
timestamp 1698431365
transform 1 0 7728 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_80
timestamp 1698431365
transform 1 0 8464 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_115
timestamp 1698431365
transform 1 0 11684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_119
timestamp 1698431365
transform 1 0 12052 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_144
timestamp 1698431365
transform 1 0 14352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_178
timestamp 1698431365
transform 1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1698431365
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1698431365
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 1698431365
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_213
timestamp 1698431365
transform 1 0 20700 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_226
timestamp 1698431365
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_238
timestamp 1698431365
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_260
timestamp 1698431365
transform 1 0 25024 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_272
timestamp 1698431365
transform 1 0 26128 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_284
timestamp 1698431365
transform 1 0 27232 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_296
timestamp 1698431365
transform 1 0 28336 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_309
timestamp 1698431365
transform 1 0 29532 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_315
timestamp 1698431365
transform 1 0 30084 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_7
timestamp 1698431365
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_19
timestamp 1698431365
transform 1 0 2852 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_31
timestamp 1698431365
transform 1 0 3956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_39
timestamp 1698431365
transform 1 0 4692 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1698431365
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1698431365
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_57
timestamp 1698431365
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_80
timestamp 1698431365
transform 1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_88
timestamp 1698431365
transform 1 0 9200 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_98
timestamp 1698431365
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_110
timestamp 1698431365
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_130
timestamp 1698431365
transform 1 0 13064 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_140
timestamp 1698431365
transform 1 0 13984 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_155
timestamp 1698431365
transform 1 0 15364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1698431365
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1698431365
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_181
timestamp 1698431365
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_197
timestamp 1698431365
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_209
timestamp 1698431365
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_225
timestamp 1698431365
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_239
timestamp 1698431365
transform 1 0 23092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_251
timestamp 1698431365
transform 1 0 24196 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_259
timestamp 1698431365
transform 1 0 24932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1698431365
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1698431365
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_305
timestamp 1698431365
transform 1 0 29164 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_313
timestamp 1698431365
transform 1 0 29900 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1698431365
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1698431365
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1698431365
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1698431365
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1698431365
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1698431365
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1698431365
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1698431365
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1698431365
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1698431365
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 1698431365
transform 1 0 11500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_122
timestamp 1698431365
transform 1 0 12328 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_141
timestamp 1698431365
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_164
timestamp 1698431365
transform 1 0 16192 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_178
timestamp 1698431365
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_190
timestamp 1698431365
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_197
timestamp 1698431365
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_213
timestamp 1698431365
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_225
timestamp 1698431365
transform 1 0 21804 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_232
timestamp 1698431365
transform 1 0 22448 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_240
timestamp 1698431365
transform 1 0 23184 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_250
timestamp 1698431365
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1698431365
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_263
timestamp 1698431365
transform 1 0 25300 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_275
timestamp 1698431365
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_287
timestamp 1698431365
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_299
timestamp 1698431365
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1698431365
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_309
timestamp 1698431365
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_317
timestamp 1698431365
transform 1 0 30268 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_7
timestamp 1698431365
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_19
timestamp 1698431365
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_31
timestamp 1698431365
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_43
timestamp 1698431365
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1698431365
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1698431365
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1698431365
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1698431365
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1698431365
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1698431365
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1698431365
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_135
timestamp 1698431365
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_147
timestamp 1698431365
transform 1 0 14628 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_156
timestamp 1698431365
transform 1 0 15456 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_176
timestamp 1698431365
transform 1 0 17296 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_186
timestamp 1698431365
transform 1 0 18216 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_205
timestamp 1698431365
transform 1 0 19964 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_213
timestamp 1698431365
transform 1 0 20700 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1698431365
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1698431365
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_230
timestamp 1698431365
transform 1 0 22264 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_238
timestamp 1698431365
transform 1 0 23000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_268
timestamp 1698431365
transform 1 0 25760 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1698431365
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1698431365
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1698431365
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_305
timestamp 1698431365
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_313
timestamp 1698431365
transform 1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1698431365
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1698431365
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1698431365
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1698431365
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1698431365
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1698431365
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1698431365
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1698431365
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1698431365
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1698431365
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1698431365
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1698431365
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_121
timestamp 1698431365
transform 1 0 12236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_127
timestamp 1698431365
transform 1 0 12788 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_134
timestamp 1698431365
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_144
timestamp 1698431365
transform 1 0 14352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_156
timestamp 1698431365
transform 1 0 15456 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_165
timestamp 1698431365
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_171
timestamp 1698431365
transform 1 0 16836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_185
timestamp 1698431365
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_197
timestamp 1698431365
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_205
timestamp 1698431365
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_223
timestamp 1698431365
transform 1 0 21620 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_230
timestamp 1698431365
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_240
timestamp 1698431365
transform 1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_246
timestamp 1698431365
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_256
timestamp 1698431365
transform 1 0 24656 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_282
timestamp 1698431365
transform 1 0 27048 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_294
timestamp 1698431365
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_306
timestamp 1698431365
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_309
timestamp 1698431365
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_317
timestamp 1698431365
transform 1 0 30268 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1698431365
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1698431365
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1698431365
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1698431365
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1698431365
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1698431365
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1698431365
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1698431365
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1698431365
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1698431365
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1698431365
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1698431365
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_113
timestamp 1698431365
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_121
timestamp 1698431365
transform 1 0 12236 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1698431365
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_173
timestamp 1698431365
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_177
timestamp 1698431365
transform 1 0 17388 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_215
timestamp 1698431365
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1698431365
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_225
timestamp 1698431365
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_234
timestamp 1698431365
transform 1 0 22632 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_254
timestamp 1698431365
transform 1 0 24472 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_260
timestamp 1698431365
transform 1 0 25024 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_264
timestamp 1698431365
transform 1 0 25392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1698431365
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1698431365
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1698431365
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_317
timestamp 1698431365
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1698431365
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1698431365
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1698431365
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1698431365
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1698431365
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1698431365
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1698431365
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1698431365
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1698431365
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1698431365
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1698431365
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1698431365
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1698431365
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1698431365
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1698431365
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1698431365
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_150
timestamp 1698431365
transform 1 0 14904 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_184
timestamp 1698431365
transform 1 0 18032 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1698431365
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_197
timestamp 1698431365
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_201
timestamp 1698431365
transform 1 0 19596 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1698431365
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_276
timestamp 1698431365
transform 1 0 26496 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_288
timestamp 1698431365
transform 1 0 27600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_300
timestamp 1698431365
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1698431365
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_317
timestamp 1698431365
transform 1 0 30268 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1698431365
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1698431365
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1698431365
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1698431365
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1698431365
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1698431365
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1698431365
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1698431365
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1698431365
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1698431365
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1698431365
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1698431365
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1698431365
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1698431365
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1698431365
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1698431365
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1698431365
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1698431365
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1698431365
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1698431365
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1698431365
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1698431365
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_217
timestamp 1698431365
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1698431365
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1698431365
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1698431365
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1698431365
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1698431365
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1698431365
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1698431365
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1698431365
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1698431365
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_317
timestamp 1698431365
transform 1 0 30268 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1698431365
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1698431365
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1698431365
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1698431365
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1698431365
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1698431365
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1698431365
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1698431365
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1698431365
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1698431365
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1698431365
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1698431365
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1698431365
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1698431365
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1698431365
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1698431365
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1698431365
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1698431365
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1698431365
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1698431365
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1698431365
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1698431365
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1698431365
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1698431365
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1698431365
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1698431365
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1698431365
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1698431365
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1698431365
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1698431365
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1698431365
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1698431365
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1698431365
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_309
timestamp 1698431365
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_317
timestamp 1698431365
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1698431365
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1698431365
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1698431365
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1698431365
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1698431365
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1698431365
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1698431365
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1698431365
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1698431365
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1698431365
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1698431365
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1698431365
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1698431365
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1698431365
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1698431365
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1698431365
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1698431365
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1698431365
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1698431365
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1698431365
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1698431365
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1698431365
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1698431365
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1698431365
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1698431365
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1698431365
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1698431365
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1698431365
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1698431365
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1698431365
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1698431365
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1698431365
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1698431365
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_317
timestamp 1698431365
transform 1 0 30268 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1698431365
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1698431365
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1698431365
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1698431365
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1698431365
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1698431365
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1698431365
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1698431365
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1698431365
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1698431365
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1698431365
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1698431365
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1698431365
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1698431365
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1698431365
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1698431365
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1698431365
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1698431365
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1698431365
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1698431365
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1698431365
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1698431365
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1698431365
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1698431365
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1698431365
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1698431365
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1698431365
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1698431365
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1698431365
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1698431365
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1698431365
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1698431365
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1698431365
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_309
timestamp 1698431365
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_317
timestamp 1698431365
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1698431365
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1698431365
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1698431365
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1698431365
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1698431365
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1698431365
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1698431365
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1698431365
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1698431365
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1698431365
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1698431365
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1698431365
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1698431365
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1698431365
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1698431365
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1698431365
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1698431365
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1698431365
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1698431365
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1698431365
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1698431365
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1698431365
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1698431365
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1698431365
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1698431365
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1698431365
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1698431365
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1698431365
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1698431365
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1698431365
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1698431365
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1698431365
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_317
timestamp 1698431365
transform 1 0 30268 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1698431365
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1698431365
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1698431365
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1698431365
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1698431365
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1698431365
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1698431365
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1698431365
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1698431365
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1698431365
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1698431365
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1698431365
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1698431365
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1698431365
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1698431365
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1698431365
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1698431365
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1698431365
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1698431365
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1698431365
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1698431365
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1698431365
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1698431365
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1698431365
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1698431365
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1698431365
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1698431365
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1698431365
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1698431365
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1698431365
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1698431365
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1698431365
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1698431365
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_309
timestamp 1698431365
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_317
timestamp 1698431365
transform 1 0 30268 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1698431365
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1698431365
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_27
timestamp 1698431365
transform 1 0 3588 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_29
timestamp 1698431365
transform 1 0 3772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_41
timestamp 1698431365
transform 1 0 4876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1698431365
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1698431365
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1698431365
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_81
timestamp 1698431365
transform 1 0 8556 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_85
timestamp 1698431365
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_97
timestamp 1698431365
transform 1 0 10028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1698431365
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_113
timestamp 1698431365
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_121
timestamp 1698431365
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_128
timestamp 1698431365
transform 1 0 12880 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_132
timestamp 1698431365
transform 1 0 13248 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_141
timestamp 1698431365
transform 1 0 14076 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_149
timestamp 1698431365
transform 1 0 14812 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_154
timestamp 1698431365
transform 1 0 15272 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_163
timestamp 1698431365
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1698431365
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1698431365
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1698431365
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_193
timestamp 1698431365
transform 1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_209
timestamp 1698431365
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_219
timestamp 1698431365
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1698431365
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1698431365
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_233
timestamp 1698431365
transform 1 0 22540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_245
timestamp 1698431365
transform 1 0 23644 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_251
timestamp 1698431365
transform 1 0 24196 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_253
timestamp 1698431365
transform 1 0 24380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_265
timestamp 1698431365
transform 1 0 25484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 1698431365
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1698431365
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1698431365
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_305
timestamp 1698431365
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_309
timestamp 1698431365
transform 1 0 29532 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_317
timestamp 1698431365
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 11592 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1698431365
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1698431365
transform 1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1698431365
transform -1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1698431365
transform -1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1698431365
transform 1 0 5060 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1698431365
transform -1 0 5336 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1698431365
transform -1 0 10120 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1698431365
transform 1 0 9476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1698431365
transform -1 0 14996 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1698431365
transform -1 0 13984 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1698431365
transform -1 0 5888 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1698431365
transform -1 0 21252 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1698431365
transform 1 0 4232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1698431365
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1698431365
transform 1 0 5060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1698431365
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1698431365
transform -1 0 25668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1698431365
transform -1 0 11040 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1698431365
transform -1 0 23092 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1698431365
transform -1 0 27416 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1698431365
transform 1 0 15272 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1698431365
transform -1 0 23828 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1698431365
transform -1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1698431365
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1698431365
transform -1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1698431365
transform -1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1698431365
transform -1 0 23644 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1698431365
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1698431365
transform 1 0 25024 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1698431365
transform -1 0 21160 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1698431365
transform -1 0 26312 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1698431365
transform -1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1698431365
transform -1 0 30544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1698431365
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1698431365
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1698431365
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1698431365
transform -1 0 30544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1698431365
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1698431365
transform 1 0 14904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1698431365
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1698431365
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1698431365
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1698431365
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input12
timestamp 1698431365
transform -1 0 30544 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1698431365
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1698431365
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1698431365
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1698431365
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1698431365
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1698431365
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1698431365
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1698431365
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1698431365
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1698431365
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 30544 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1698431365
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1698431365
transform -1 0 13248 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform -1 0 30544 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1698431365
transform -1 0 30544 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1698431365
transform -1 0 30544 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1698431365
transform -1 0 30544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1698431365
transform -1 0 30544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1698431365
transform -1 0 30544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1698431365
transform 1 0 21344 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 1380 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1698431365
transform -1 0 12880 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1698431365
transform 1 0 19780 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1698431365
transform 1 0 20700 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1698431365
transform 1 0 30176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1698431365
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1698431365
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1698431365
transform 1 0 19228 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1698431365
transform -1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1698431365
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1698431365
transform -1 0 16560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1698431365
transform 1 0 30176 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1698431365
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1698431365
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1698431365
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1698431365
transform -1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1698431365
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1698431365
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1698431365
transform 1 0 30176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1698431365
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1698431365
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1698431365
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1698431365
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1698431365
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1698431365
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1698431365
transform -1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1698431365
transform -1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1698431365
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1698431365
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1698431365
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1698431365
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1698431365
transform 1 0 21988 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1698431365
transform 1 0 30176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1698431365
transform 1 0 30176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1698431365
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1698431365
transform 1 0 30176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1698431365
transform 1 0 30176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1698431365
transform 1 0 30176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1698431365
transform -1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1698431365
transform 1 0 15548 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1698431365
transform -1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_50
timestamp 1698431365
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_51
timestamp 1698431365
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 30820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_52
timestamp 1698431365
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 30820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_53
timestamp 1698431365
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 30820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_54
timestamp 1698431365
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_55
timestamp 1698431365
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 30820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_56
timestamp 1698431365
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 30820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_57
timestamp 1698431365
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 30820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_58
timestamp 1698431365
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 30820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_59
timestamp 1698431365
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_60
timestamp 1698431365
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_61
timestamp 1698431365
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 30820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_62
timestamp 1698431365
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 30820 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_63
timestamp 1698431365
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 30820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_64
timestamp 1698431365
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 30820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_65
timestamp 1698431365
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 30820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_66
timestamp 1698431365
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 30820 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_67
timestamp 1698431365
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_68
timestamp 1698431365
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 30820 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_69
timestamp 1698431365
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 30820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_70
timestamp 1698431365
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 30820 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_71
timestamp 1698431365
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 30820 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_72
timestamp 1698431365
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_73
timestamp 1698431365
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 30820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_74
timestamp 1698431365
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 30820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_75
timestamp 1698431365
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 30820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_76
timestamp 1698431365
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_77
timestamp 1698431365
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 30820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_78
timestamp 1698431365
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_79
timestamp 1698431365
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 30820 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_80
timestamp 1698431365
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 30820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_81
timestamp 1698431365
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 30820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_82
timestamp 1698431365
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 30820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_83
timestamp 1698431365
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 30820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_84
timestamp 1698431365
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 30820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_85
timestamp 1698431365
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 30820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_86
timestamp 1698431365
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_87
timestamp 1698431365
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 30820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_88
timestamp 1698431365
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 30820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_89
timestamp 1698431365
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 30820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_90
timestamp 1698431365
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 30820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_91
timestamp 1698431365
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_92
timestamp 1698431365
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_93
timestamp 1698431365
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 30820 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_94
timestamp 1698431365
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 30820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_95
timestamp 1698431365
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 30820 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_96
timestamp 1698431365
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 30820 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_97
timestamp 1698431365
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_98
timestamp 1698431365
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_99
timestamp 1698431365
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 30820 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 22908 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1698431365
transform -1 0 26956 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698431365
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1698431365
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1698431365
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1698431365
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1698431365
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1698431365
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1698431365
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1698431365
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp 1698431365
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp 1698431365
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp 1698431365
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 1698431365
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 1698431365
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_113
timestamp 1698431365
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_114
timestamp 1698431365
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_115
timestamp 1698431365
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 1698431365
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 1698431365
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_118
timestamp 1698431365
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_119
timestamp 1698431365
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_120
timestamp 1698431365
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_121
timestamp 1698431365
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 1698431365
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_123
timestamp 1698431365
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp 1698431365
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_125
timestamp 1698431365
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_126
timestamp 1698431365
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1698431365
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_128
timestamp 1698431365
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_129
timestamp 1698431365
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_130
timestamp 1698431365
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_131
timestamp 1698431365
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_132
timestamp 1698431365
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_133
timestamp 1698431365
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_134
timestamp 1698431365
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_135
timestamp 1698431365
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_136
timestamp 1698431365
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_137
timestamp 1698431365
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_138
timestamp 1698431365
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_139
timestamp 1698431365
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_140
timestamp 1698431365
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_141
timestamp 1698431365
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_142
timestamp 1698431365
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_143
timestamp 1698431365
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_144
timestamp 1698431365
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_145
timestamp 1698431365
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_146
timestamp 1698431365
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_147
timestamp 1698431365
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_148
timestamp 1698431365
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_149
timestamp 1698431365
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_150
timestamp 1698431365
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_151
timestamp 1698431365
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_152
timestamp 1698431365
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_153
timestamp 1698431365
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_154
timestamp 1698431365
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_155
timestamp 1698431365
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_156
timestamp 1698431365
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_157
timestamp 1698431365
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_158
timestamp 1698431365
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_159
timestamp 1698431365
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_160
timestamp 1698431365
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_161
timestamp 1698431365
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_162
timestamp 1698431365
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_163
timestamp 1698431365
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_164
timestamp 1698431365
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_165
timestamp 1698431365
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_166
timestamp 1698431365
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_167
timestamp 1698431365
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_168
timestamp 1698431365
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_169
timestamp 1698431365
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_170
timestamp 1698431365
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_171
timestamp 1698431365
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_172
timestamp 1698431365
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_173
timestamp 1698431365
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_174
timestamp 1698431365
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_175
timestamp 1698431365
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_176
timestamp 1698431365
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_177
timestamp 1698431365
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_178
timestamp 1698431365
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_179
timestamp 1698431365
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_180
timestamp 1698431365
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_181
timestamp 1698431365
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_182
timestamp 1698431365
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_183
timestamp 1698431365
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_184
timestamp 1698431365
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_185
timestamp 1698431365
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_186
timestamp 1698431365
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_187
timestamp 1698431365
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_188
timestamp 1698431365
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_189
timestamp 1698431365
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_190
timestamp 1698431365
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_191
timestamp 1698431365
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_192
timestamp 1698431365
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_193
timestamp 1698431365
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_194
timestamp 1698431365
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_195
timestamp 1698431365
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_196
timestamp 1698431365
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_197
timestamp 1698431365
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_198
timestamp 1698431365
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_199
timestamp 1698431365
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_200
timestamp 1698431365
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_201
timestamp 1698431365
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_202
timestamp 1698431365
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_203
timestamp 1698431365
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_204
timestamp 1698431365
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_205
timestamp 1698431365
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_206
timestamp 1698431365
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_207
timestamp 1698431365
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_208
timestamp 1698431365
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_209
timestamp 1698431365
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_210
timestamp 1698431365
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_211
timestamp 1698431365
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_212
timestamp 1698431365
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_213
timestamp 1698431365
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_214
timestamp 1698431365
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_215
timestamp 1698431365
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_216
timestamp 1698431365
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_217
timestamp 1698431365
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_218
timestamp 1698431365
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_219
timestamp 1698431365
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_220
timestamp 1698431365
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_221
timestamp 1698431365
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_222
timestamp 1698431365
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_223
timestamp 1698431365
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_224
timestamp 1698431365
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_225
timestamp 1698431365
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_226
timestamp 1698431365
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_227
timestamp 1698431365
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_228
timestamp 1698431365
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_229
timestamp 1698431365
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_230
timestamp 1698431365
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_231
timestamp 1698431365
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_232
timestamp 1698431365
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_233
timestamp 1698431365
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_234
timestamp 1698431365
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_235
timestamp 1698431365
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_236
timestamp 1698431365
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_237
timestamp 1698431365
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_238
timestamp 1698431365
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_239
timestamp 1698431365
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_240
timestamp 1698431365
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_241
timestamp 1698431365
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_242
timestamp 1698431365
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_243
timestamp 1698431365
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_244
timestamp 1698431365
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_245
timestamp 1698431365
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_246
timestamp 1698431365
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_247
timestamp 1698431365
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_248
timestamp 1698431365
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_249
timestamp 1698431365
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_250
timestamp 1698431365
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_251
timestamp 1698431365
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_252
timestamp 1698431365
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_253
timestamp 1698431365
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_254
timestamp 1698431365
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_255
timestamp 1698431365
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_256
timestamp 1698431365
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_257
timestamp 1698431365
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_258
timestamp 1698431365
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_259
timestamp 1698431365
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_260
timestamp 1698431365
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_261
timestamp 1698431365
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_262
timestamp 1698431365
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_263
timestamp 1698431365
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_264
timestamp 1698431365
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_265
timestamp 1698431365
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_266
timestamp 1698431365
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_267
timestamp 1698431365
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_268
timestamp 1698431365
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_269
timestamp 1698431365
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_270
timestamp 1698431365
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_271
timestamp 1698431365
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_272
timestamp 1698431365
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_273
timestamp 1698431365
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_274
timestamp 1698431365
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_275
timestamp 1698431365
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_276
timestamp 1698431365
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_277
timestamp 1698431365
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_278
timestamp 1698431365
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_279
timestamp 1698431365
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_280
timestamp 1698431365
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_281
timestamp 1698431365
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_282
timestamp 1698431365
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_283
timestamp 1698431365
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_284
timestamp 1698431365
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_285
timestamp 1698431365
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_286
timestamp 1698431365
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_287
timestamp 1698431365
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_288
timestamp 1698431365
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_289
timestamp 1698431365
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_290
timestamp 1698431365
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_291
timestamp 1698431365
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_292
timestamp 1698431365
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_293
timestamp 1698431365
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_294
timestamp 1698431365
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_295
timestamp 1698431365
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_296
timestamp 1698431365
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_297
timestamp 1698431365
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_298
timestamp 1698431365
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_299
timestamp 1698431365
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_300
timestamp 1698431365
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_301
timestamp 1698431365
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_302
timestamp 1698431365
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_303
timestamp 1698431365
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_304
timestamp 1698431365
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_305
timestamp 1698431365
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_306
timestamp 1698431365
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_307
timestamp 1698431365
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_308
timestamp 1698431365
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_309
timestamp 1698431365
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_310
timestamp 1698431365
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_311
timestamp 1698431365
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_312
timestamp 1698431365
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_313
timestamp 1698431365
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_314
timestamp 1698431365
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_315
timestamp 1698431365
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_316
timestamp 1698431365
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_317
timestamp 1698431365
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_318
timestamp 1698431365
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_319
timestamp 1698431365
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_320
timestamp 1698431365
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_321
timestamp 1698431365
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_322
timestamp 1698431365
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_323
timestamp 1698431365
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_324
timestamp 1698431365
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_325
timestamp 1698431365
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_326
timestamp 1698431365
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_327
timestamp 1698431365
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_328
timestamp 1698431365
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_329
timestamp 1698431365
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_330
timestamp 1698431365
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_331
timestamp 1698431365
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_332
timestamp 1698431365
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_333
timestamp 1698431365
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_334
timestamp 1698431365
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_335
timestamp 1698431365
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_336
timestamp 1698431365
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_337
timestamp 1698431365
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_338
timestamp 1698431365
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_339
timestamp 1698431365
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_340
timestamp 1698431365
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_341
timestamp 1698431365
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_342
timestamp 1698431365
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_343
timestamp 1698431365
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_344
timestamp 1698431365
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_345
timestamp 1698431365
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_346
timestamp 1698431365
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_347
timestamp 1698431365
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_348
timestamp 1698431365
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_349
timestamp 1698431365
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_350
timestamp 1698431365
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_351
timestamp 1698431365
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_352
timestamp 1698431365
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_353
timestamp 1698431365
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_354
timestamp 1698431365
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_355
timestamp 1698431365
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_356
timestamp 1698431365
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_357
timestamp 1698431365
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_358
timestamp 1698431365
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_359
timestamp 1698431365
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_360
timestamp 1698431365
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_361
timestamp 1698431365
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_362
timestamp 1698431365
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_363
timestamp 1698431365
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_364
timestamp 1698431365
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_365
timestamp 1698431365
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_366
timestamp 1698431365
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_367
timestamp 1698431365
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_368
timestamp 1698431365
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_369
timestamp 1698431365
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_370
timestamp 1698431365
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_371
timestamp 1698431365
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_372
timestamp 1698431365
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_373
timestamp 1698431365
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_374
timestamp 1698431365
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_375
timestamp 1698431365
transform 1 0 3680 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_376
timestamp 1698431365
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_377
timestamp 1698431365
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_378
timestamp 1698431365
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_379
timestamp 1698431365
transform 1 0 13984 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_380
timestamp 1698431365
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_381
timestamp 1698431365
transform 1 0 19136 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_382
timestamp 1698431365
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_383
timestamp 1698431365
transform 1 0 24288 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_384
timestamp 1698431365
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_385
timestamp 1698431365
transform 1 0 29440 0 -1 29376
box -38 -48 130 592
<< labels >>
flabel metal4 s 5318 2128 5638 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12746 2128 13066 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 20174 2128 20494 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27602 2128 27922 29424 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6076 30868 6396 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12876 30868 13196 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 19676 30868 19996 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 26476 30868 26796 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4658 2128 4978 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12086 2128 12406 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19514 2128 19834 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26942 2128 27262 29424 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5416 30868 5736 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12216 30868 12536 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 19016 30868 19336 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 25816 30868 26136 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 clock
port 2 nsew signal input
flabel metal2 s 12254 31200 12310 32000 0 FreeSans 224 90 0 0 clock_o
port 3 nsew signal tristate
flabel metal2 s 19338 31200 19394 32000 0 FreeSans 224 90 0 0 ram_addr_o[0]
port 4 nsew signal tristate
flabel metal2 s 20626 31200 20682 32000 0 FreeSans 224 90 0 0 ram_addr_o[1]
port 5 nsew signal tristate
flabel metal3 s 31200 19728 32000 19848 0 FreeSans 480 0 0 0 ram_addr_o[2]
port 6 nsew signal tristate
flabel metal3 s 31200 20408 32000 20528 0 FreeSans 480 0 0 0 ram_addr_o[3]
port 7 nsew signal tristate
flabel metal3 s 31200 21088 32000 21208 0 FreeSans 480 0 0 0 ram_addr_o[4]
port 8 nsew signal tristate
flabel metal3 s 31200 16328 32000 16448 0 FreeSans 480 0 0 0 ram_data_i[0]
port 9 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 ram_data_i[10]
port 10 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 ram_data_i[11]
port 11 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 ram_data_i[12]
port 12 nsew signal input
flabel metal3 s 31200 12248 32000 12368 0 FreeSans 480 0 0 0 ram_data_i[13]
port 13 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 ram_data_i[14]
port 14 nsew signal input
flabel metal2 s 14830 31200 14886 32000 0 FreeSans 224 90 0 0 ram_data_i[15]
port 15 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 ram_data_i[16]
port 16 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 ram_data_i[17]
port 17 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 ram_data_i[18]
port 18 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 ram_data_i[19]
port 19 nsew signal input
flabel metal3 s 31200 22448 32000 22568 0 FreeSans 480 0 0 0 ram_data_i[1]
port 20 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 ram_data_i[20]
port 21 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 ram_data_i[21]
port 22 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 ram_data_i[22]
port 23 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ram_data_i[23]
port 24 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 ram_data_i[24]
port 25 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 ram_data_i[25]
port 26 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 ram_data_i[26]
port 27 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 ram_data_i[27]
port 28 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 ram_data_i[28]
port 29 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 ram_data_i[29]
port 30 nsew signal input
flabel metal3 s 31200 19048 32000 19168 0 FreeSans 480 0 0 0 ram_data_i[2]
port 31 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 ram_data_i[30]
port 32 nsew signal input
flabel metal2 s 12898 31200 12954 32000 0 FreeSans 224 90 0 0 ram_data_i[31]
port 33 nsew signal input
flabel metal3 s 31200 21768 32000 21888 0 FreeSans 480 0 0 0 ram_data_i[3]
port 34 nsew signal input
flabel metal3 s 31200 23128 32000 23248 0 FreeSans 480 0 0 0 ram_data_i[4]
port 35 nsew signal input
flabel metal3 s 31200 13608 32000 13728 0 FreeSans 480 0 0 0 ram_data_i[5]
port 36 nsew signal input
flabel metal3 s 31200 10888 32000 11008 0 FreeSans 480 0 0 0 ram_data_i[6]
port 37 nsew signal input
flabel metal3 s 31200 10208 32000 10328 0 FreeSans 480 0 0 0 ram_data_i[7]
port 38 nsew signal input
flabel metal3 s 31200 9528 32000 9648 0 FreeSans 480 0 0 0 ram_data_i[8]
port 39 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 ram_data_i[9]
port 40 nsew signal input
flabel metal2 s 18694 31200 18750 32000 0 FreeSans 224 90 0 0 ram_data_o[0]
port 41 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 ram_data_o[10]
port 42 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 ram_data_o[11]
port 43 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 ram_data_o[12]
port 44 nsew signal tristate
flabel metal3 s 31200 14288 32000 14408 0 FreeSans 480 0 0 0 ram_data_o[13]
port 45 nsew signal tristate
flabel metal3 s 31200 15648 32000 15768 0 FreeSans 480 0 0 0 ram_data_o[14]
port 46 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 ram_data_o[15]
port 47 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 ram_data_o[16]
port 48 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 ram_data_o[17]
port 49 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 ram_data_o[18]
port 50 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 ram_data_o[19]
port 51 nsew signal tristate
flabel metal3 s 31200 17688 32000 17808 0 FreeSans 480 0 0 0 ram_data_o[1]
port 52 nsew signal tristate
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 ram_data_o[20]
port 53 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 ram_data_o[21]
port 54 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 ram_data_o[22]
port 55 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 ram_data_o[23]
port 56 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 ram_data_o[24]
port 57 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 ram_data_o[25]
port 58 nsew signal tristate
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 ram_data_o[26]
port 59 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 ram_data_o[27]
port 60 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 ram_data_o[28]
port 61 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 ram_data_o[29]
port 62 nsew signal tristate
flabel metal3 s 31200 18368 32000 18488 0 FreeSans 480 0 0 0 ram_data_o[2]
port 63 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 ram_data_o[30]
port 64 nsew signal tristate
flabel metal2 s 21914 31200 21970 32000 0 FreeSans 224 90 0 0 ram_data_o[31]
port 65 nsew signal tristate
flabel metal3 s 31200 17008 32000 17128 0 FreeSans 480 0 0 0 ram_data_o[3]
port 66 nsew signal tristate
flabel metal3 s 31200 14968 32000 15088 0 FreeSans 480 0 0 0 ram_data_o[4]
port 67 nsew signal tristate
flabel metal3 s 31200 12928 32000 13048 0 FreeSans 480 0 0 0 ram_data_o[5]
port 68 nsew signal tristate
flabel metal3 s 31200 11568 32000 11688 0 FreeSans 480 0 0 0 ram_data_o[6]
port 69 nsew signal tristate
flabel metal3 s 31200 8848 32000 8968 0 FreeSans 480 0 0 0 ram_data_o[7]
port 70 nsew signal tristate
flabel metal3 s 31200 8168 32000 8288 0 FreeSans 480 0 0 0 ram_data_o[8]
port 71 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 ram_data_o[9]
port 72 nsew signal tristate
flabel metal2 s 15474 31200 15530 32000 0 FreeSans 224 90 0 0 ram_rw_en_o
port 73 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 reset_i
port 74 nsew signal input
flabel metal2 s 14186 31200 14242 32000 0 FreeSans 224 90 0 0 stop_lamp_o
port 75 nsew signal tristate
rlabel metal1 15962 29376 15962 29376 0 VGND
rlabel metal1 15962 28832 15962 28832 0 VPWR
rlabel metal1 12742 22746 12742 22746 0 _0000_
rlabel metal2 19458 24990 19458 24990 0 _0001_
rlabel metal1 21252 25670 21252 25670 0 _0002_
rlabel metal1 22908 24922 22908 24922 0 _0003_
rlabel metal2 25254 25058 25254 25058 0 _0004_
rlabel metal2 26082 23970 26082 23970 0 _0005_
rlabel metal1 18637 17646 18637 17646 0 _0006_
rlabel metal2 19366 17000 19366 17000 0 _0007_
rlabel metal1 23506 18775 23506 18775 0 _0008_
rlabel metal1 26963 17578 26963 17578 0 _0009_
rlabel metal1 23743 15470 23743 15470 0 _0010_
rlabel metal2 21022 13464 21022 13464 0 _0011_
rlabel metal2 26266 10914 26266 10914 0 _0012_
rlabel metal1 24380 8602 24380 8602 0 _0013_
rlabel metal1 23092 8058 23092 8058 0 _0014_
rlabel metal2 20102 7208 20102 7208 0 _0015_
rlabel metal1 17664 6766 17664 6766 0 _0016_
rlabel metal1 15548 9554 15548 9554 0 _0017_
rlabel metal1 15180 10778 15180 10778 0 _0018_
rlabel metal1 20470 14042 20470 14042 0 _0019_
rlabel metal1 17243 16150 17243 16150 0 _0020_
rlabel metal1 12742 15130 12742 15130 0 _0021_
rlabel metal2 10534 14110 10534 14110 0 _0022_
rlabel metal2 12374 14110 12374 14110 0 _0023_
rlabel metal1 13255 7446 13255 7446 0 _0024_
rlabel metal1 10311 7446 10311 7446 0 _0025_
rlabel metal2 5750 7650 5750 7650 0 _0026_
rlabel metal1 4600 9146 4600 9146 0 _0027_
rlabel metal1 4232 11322 4232 11322 0 _0028_
rlabel metal1 4745 12886 4745 12886 0 _0029_
rlabel metal2 4278 13736 4278 13736 0 _0030_
rlabel metal1 4423 16150 4423 16150 0 _0031_
rlabel metal1 5067 19414 5067 19414 0 _0032_
rlabel metal1 6946 20026 6946 20026 0 _0033_
rlabel metal1 10955 15402 10955 15402 0 _0034_
rlabel metal1 9660 20774 9660 20774 0 _0035_
rlabel metal2 11270 19992 11270 19992 0 _0036_
rlabel metal2 12466 21352 12466 21352 0 _0037_
rlabel metal1 18683 20842 18683 20842 0 _0038_
rlabel metal1 19780 20230 19780 20230 0 _0039_
rlabel metal1 21712 19482 21712 19482 0 _0040_
rlabel metal1 25852 18394 25852 18394 0 _0041_
rlabel metal1 24104 20026 24104 20026 0 _0042_
rlabel metal2 17526 19652 17526 19652 0 _0043_
rlabel metal1 15364 17306 15364 17306 0 _0044_
rlabel metal2 15870 20230 15870 20230 0 _0045_
rlabel metal2 17250 25058 17250 25058 0 _0046_
rlabel metal2 15778 24990 15778 24990 0 _0047_
rlabel metal2 14214 24582 14214 24582 0 _0048_
rlabel metal1 13945 21930 13945 21930 0 _0049_
rlabel metal1 18906 24378 18906 24378 0 _0050_
rlabel metal1 20424 24922 20424 24922 0 _0051_
rlabel metal2 22586 25024 22586 25024 0 _0052_
rlabel metal1 24564 24922 24564 24922 0 _0053_
rlabel metal1 25438 24072 25438 24072 0 _0054_
rlabel metal1 17243 17578 17243 17578 0 _0055_
rlabel metal1 19090 16694 19090 16694 0 _0056_
rlabel metal2 22402 18530 22402 18530 0 _0057_
rlabel metal1 24978 17306 24978 17306 0 _0058_
rlabel metal1 22402 15402 22402 15402 0 _0059_
rlabel metal2 20562 13090 20562 13090 0 _0060_
rlabel metal2 25714 11356 25714 11356 0 _0061_
rlabel metal1 23368 9146 23368 9146 0 _0062_
rlabel metal2 22126 9214 22126 9214 0 _0063_
rlabel metal1 19412 7446 19412 7446 0 _0064_
rlabel metal1 17020 7446 17020 7446 0 _0065_
rlabel metal1 15134 9452 15134 9452 0 _0066_
rlabel metal1 15962 11050 15962 11050 0 _0067_
rlabel metal1 19412 15062 19412 15062 0 _0068_
rlabel metal1 16284 15334 16284 15334 0 _0069_
rlabel metal1 12190 15130 12190 15130 0 _0070_
rlabel metal1 10074 13498 10074 13498 0 _0071_
rlabel metal1 11868 13498 11868 13498 0 _0072_
rlabel metal1 11868 6970 11868 6970 0 _0073_
rlabel metal1 8694 7310 8694 7310 0 _0074_
rlabel metal1 6670 7922 6670 7922 0 _0075_
rlabel metal1 5796 9486 5796 9486 0 _0076_
rlabel metal1 3358 11322 3358 11322 0 _0077_
rlabel metal1 5336 12750 5336 12750 0 _0078_
rlabel metal1 4692 13974 4692 13974 0 _0079_
rlabel metal1 4600 15674 4600 15674 0 _0080_
rlabel metal1 3726 18938 3726 18938 0 _0081_
rlabel metal1 6716 18938 6716 18938 0 _0082_
rlabel via1 9331 15674 9331 15674 0 _0083_
rlabel metal2 8602 20196 8602 20196 0 _0084_
rlabel metal1 11546 18938 11546 18938 0 _0085_
rlabel metal1 11868 21454 11868 21454 0 _0086_
rlabel metal1 17342 20570 17342 20570 0 _0087_
rlabel metal1 19458 19754 19458 19754 0 _0088_
rlabel metal1 21482 18938 21482 18938 0 _0089_
rlabel metal1 25116 18938 25116 18938 0 _0090_
rlabel metal1 23506 20026 23506 20026 0 _0091_
rlabel metal2 16974 19108 16974 19108 0 _0092_
rlabel metal1 14260 17578 14260 17578 0 _0093_
rlabel metal2 14766 20638 14766 20638 0 _0094_
rlabel metal1 10304 21658 10304 21658 0 _0095_
rlabel metal1 13754 21658 13754 21658 0 _0096_
rlabel metal1 8556 21862 8556 21862 0 _0097_
rlabel metal1 5285 20842 5285 20842 0 _0098_
rlabel metal1 5382 21454 5382 21454 0 _0099_
rlabel metal2 6394 21794 6394 21794 0 _0100_
rlabel metal1 15870 22406 15870 22406 0 _0101_
rlabel metal1 13846 21420 13846 21420 0 _0102_
rlabel metal2 15502 21930 15502 21930 0 _0103_
rlabel metal1 14536 19890 14536 19890 0 _0104_
rlabel metal2 15226 20468 15226 20468 0 _0105_
rlabel metal1 14076 17306 14076 17306 0 _0106_
rlabel metal1 17296 18734 17296 18734 0 _0107_
rlabel metal1 23874 19856 23874 19856 0 _0108_
rlabel metal1 25392 18734 25392 18734 0 _0109_
rlabel metal1 21850 18734 21850 18734 0 _0110_
rlabel metal2 19458 19176 19458 19176 0 _0111_
rlabel metal1 18906 22474 18906 22474 0 _0112_
rlabel metal1 17756 20434 17756 20434 0 _0113_
rlabel metal1 16376 18734 16376 18734 0 _0114_
rlabel metal1 21160 15470 21160 15470 0 _0115_
rlabel metal1 6946 12138 6946 12138 0 _0116_
rlabel metal1 13616 14926 13616 14926 0 _0117_
rlabel metal1 17710 8058 17710 8058 0 _0118_
rlabel metal1 14674 22406 14674 22406 0 _0119_
rlabel metal1 15042 19142 15042 19142 0 _0120_
rlabel metal1 22540 16626 22540 16626 0 _0121_
rlabel metal1 22218 12920 22218 12920 0 _0122_
rlabel metal2 22034 11152 22034 11152 0 _0123_
rlabel metal2 21666 11526 21666 11526 0 _0124_
rlabel metal1 20424 10438 20424 10438 0 _0125_
rlabel metal2 18446 10948 18446 10948 0 _0126_
rlabel metal1 16238 13328 16238 13328 0 _0127_
rlabel metal1 14766 12852 14766 12852 0 _0128_
rlabel viali 13110 12207 13110 12207 0 _0129_
rlabel metal1 8372 8874 8372 8874 0 _0130_
rlabel metal1 5980 12818 5980 12818 0 _0131_
rlabel metal1 6256 13498 6256 13498 0 _0132_
rlabel via1 5658 15453 5658 15453 0 _0133_
rlabel metal1 6716 17306 6716 17306 0 _0134_
rlabel metal1 13018 17306 13018 17306 0 _0135_
rlabel metal1 13662 19278 13662 19278 0 _0136_
rlabel metal1 13340 18666 13340 18666 0 _0137_
rlabel metal1 9522 16592 9522 16592 0 _0138_
rlabel metal1 25990 15538 25990 15538 0 _0139_
rlabel metal1 24978 16592 24978 16592 0 _0140_
rlabel metal1 22862 18224 22862 18224 0 _0141_
rlabel metal1 21160 18394 21160 18394 0 _0142_
rlabel metal1 21022 18258 21022 18258 0 _0143_
rlabel metal1 21206 18224 21206 18224 0 _0144_
rlabel metal1 22218 18292 22218 18292 0 _0145_
rlabel metal2 22862 17476 22862 17476 0 _0146_
rlabel metal1 24702 13328 24702 13328 0 _0147_
rlabel metal1 24426 12818 24426 12818 0 _0148_
rlabel metal1 25714 13294 25714 13294 0 _0149_
rlabel metal2 24794 14348 24794 14348 0 _0150_
rlabel metal1 24518 13906 24518 13906 0 _0151_
rlabel metal1 24978 13702 24978 13702 0 _0152_
rlabel metal1 25806 14586 25806 14586 0 _0153_
rlabel metal1 25898 16694 25898 16694 0 _0154_
rlabel metal2 24978 14144 24978 14144 0 _0155_
rlabel metal1 24058 11730 24058 11730 0 _0156_
rlabel metal1 24610 10608 24610 10608 0 _0157_
rlabel metal1 23736 10234 23736 10234 0 _0158_
rlabel metal1 23966 11866 23966 11866 0 _0159_
rlabel metal1 24334 12342 24334 12342 0 _0160_
rlabel metal1 21482 12240 21482 12240 0 _0161_
rlabel metal1 24334 11798 24334 11798 0 _0162_
rlabel metal1 21206 12172 21206 12172 0 _0163_
rlabel metal1 16606 9010 16606 9010 0 _0164_
rlabel metal1 18676 8874 18676 8874 0 _0165_
rlabel metal2 18354 9316 18354 9316 0 _0166_
rlabel metal1 21022 8398 21022 8398 0 _0167_
rlabel metal1 21482 7990 21482 7990 0 _0168_
rlabel metal1 20930 9350 20930 9350 0 _0169_
rlabel metal1 21482 8466 21482 8466 0 _0170_
rlabel metal1 22586 9010 22586 9010 0 _0171_
rlabel metal1 21022 9962 21022 9962 0 _0172_
rlabel metal1 20010 11798 20010 11798 0 _0173_
rlabel metal1 16790 15028 16790 15028 0 _0174_
rlabel metal1 14812 14994 14812 14994 0 _0175_
rlabel metal1 17802 11730 17802 11730 0 _0176_
rlabel metal1 18078 11696 18078 11696 0 _0177_
rlabel metal1 17342 12206 17342 12206 0 _0178_
rlabel metal1 19136 13906 19136 13906 0 _0179_
rlabel metal1 18584 14246 18584 14246 0 _0180_
rlabel metal1 18906 13294 18906 13294 0 _0181_
rlabel metal1 17158 12784 17158 12784 0 _0182_
rlabel metal1 21027 12200 21027 12200 0 _0183_
rlabel metal1 13570 12240 13570 12240 0 _0184_
rlabel metal1 15180 9690 15180 9690 0 _0185_
rlabel metal2 18998 9180 18998 9180 0 _0186_
rlabel metal1 17526 8534 17526 8534 0 _0187_
rlabel metal1 17020 9146 17020 9146 0 _0188_
rlabel metal2 17802 11016 17802 11016 0 _0189_
rlabel metal1 17986 13974 17986 13974 0 _0190_
rlabel metal1 17388 14314 17388 14314 0 _0191_
rlabel metal1 17342 12852 17342 12852 0 _0192_
rlabel metal1 14490 14586 14490 14586 0 _0193_
rlabel metal1 15226 14450 15226 14450 0 _0194_
rlabel metal1 14214 13974 14214 13974 0 _0195_
rlabel metal1 17480 12818 17480 12818 0 _0196_
rlabel metal1 15226 12716 15226 12716 0 _0197_
rlabel metal1 5566 11152 5566 11152 0 _0198_
rlabel metal2 6118 11322 6118 11322 0 _0199_
rlabel metal1 6854 11152 6854 11152 0 _0200_
rlabel metal1 8694 12886 8694 12886 0 _0201_
rlabel metal1 8740 12614 8740 12614 0 _0202_
rlabel metal1 8004 11662 8004 11662 0 _0203_
rlabel metal1 8326 11186 8326 11186 0 _0204_
rlabel metal1 8372 8466 8372 8466 0 _0205_
rlabel metal1 7820 7990 7820 7990 0 _0206_
rlabel metal2 8418 9384 8418 9384 0 _0207_
rlabel metal2 6394 9282 6394 9282 0 _0208_
rlabel metal1 7406 9690 7406 9690 0 _0209_
rlabel metal1 6670 10676 6670 10676 0 _0210_
rlabel metal1 8188 10098 8188 10098 0 _0211_
rlabel metal1 8510 11764 8510 11764 0 _0212_
rlabel metal1 12466 12172 12466 12172 0 _0213_
rlabel metal1 11592 11730 11592 11730 0 _0214_
rlabel metal1 10902 11662 10902 11662 0 _0215_
rlabel metal1 13754 10438 13754 10438 0 _0216_
rlabel metal1 13754 10676 13754 10676 0 _0217_
rlabel metal1 13294 10540 13294 10540 0 _0218_
rlabel metal2 10718 8772 10718 8772 0 _0219_
rlabel metal2 10258 10642 10258 10642 0 _0220_
rlabel metal1 12834 9520 12834 9520 0 _0221_
rlabel metal1 12926 8602 12926 8602 0 _0222_
rlabel metal2 11638 9826 11638 9826 0 _0223_
rlabel metal2 10626 10591 10626 10591 0 _0224_
rlabel metal2 9890 12036 9890 12036 0 _0225_
rlabel metal1 9154 14246 9154 14246 0 _0226_
rlabel metal1 11776 10030 11776 10030 0 _0227_
rlabel metal1 10258 10710 10258 10710 0 _0228_
rlabel metal1 10074 10472 10074 10472 0 _0229_
rlabel metal1 6992 11118 6992 11118 0 _0230_
rlabel metal1 8556 11322 8556 11322 0 _0231_
rlabel metal2 9062 12648 9062 12648 0 _0232_
rlabel metal2 8970 13940 8970 13940 0 _0233_
rlabel metal1 7544 18190 7544 18190 0 _0234_
rlabel metal2 7038 18462 7038 18462 0 _0235_
rlabel metal1 6762 18734 6762 18734 0 _0236_
rlabel metal1 7038 17646 7038 17646 0 _0237_
rlabel metal1 8556 16626 8556 16626 0 _0238_
rlabel metal1 6946 15402 6946 15402 0 _0239_
rlabel metal1 7038 15878 7038 15878 0 _0240_
rlabel metal2 8050 15266 8050 15266 0 _0241_
rlabel metal1 7866 14450 7866 14450 0 _0242_
rlabel metal1 7636 14382 7636 14382 0 _0243_
rlabel metal1 8418 14314 8418 14314 0 _0244_
rlabel metal2 9706 15844 9706 15844 0 _0245_
rlabel metal1 7682 16558 7682 16558 0 _0246_
rlabel metal2 8970 16932 8970 16932 0 _0247_
rlabel metal2 8142 19652 8142 19652 0 _0248_
rlabel metal1 7728 19482 7728 19482 0 _0249_
rlabel metal1 8832 17170 8832 17170 0 _0250_
rlabel metal1 11546 16048 11546 16048 0 _0251_
rlabel metal1 9522 17170 9522 17170 0 _0252_
rlabel metal1 9614 17680 9614 17680 0 _0253_
rlabel metal1 9982 18734 9982 18734 0 _0254_
rlabel metal1 10718 18768 10718 18768 0 _0255_
rlabel metal2 10442 17952 10442 17952 0 _0256_
rlabel metal1 12788 18258 12788 18258 0 _0257_
rlabel metal1 11500 18258 11500 18258 0 _0258_
rlabel metal2 11822 18564 11822 18564 0 _0259_
rlabel metal1 13248 18734 13248 18734 0 _0260_
rlabel metal1 13248 19346 13248 19346 0 _0261_
rlabel metal1 14122 18870 14122 18870 0 _0262_
rlabel metal1 13340 18938 13340 18938 0 _0263_
rlabel metal1 12788 19278 12788 19278 0 _0264_
rlabel metal1 16100 17170 16100 17170 0 _0265_
rlabel metal2 12098 19618 12098 19618 0 _0266_
rlabel metal1 15870 17306 15870 17306 0 _0267_
rlabel metal1 13524 16490 13524 16490 0 _0268_
rlabel metal1 13148 16490 13148 16490 0 _0269_
rlabel metal1 12788 16762 12788 16762 0 _0270_
rlabel metal1 20424 13158 20424 13158 0 _0271_
rlabel metal1 11178 18224 11178 18224 0 _0272_
rlabel metal1 11500 18190 11500 18190 0 _0273_
rlabel metal1 13202 16422 13202 16422 0 _0274_
rlabel metal1 19044 16082 19044 16082 0 _0275_
rlabel metal1 14490 9554 14490 9554 0 _0276_
rlabel metal1 11592 18394 11592 18394 0 _0277_
rlabel metal1 16422 14348 16422 14348 0 _0278_
rlabel metal1 9614 18156 9614 18156 0 _0279_
rlabel metal1 9476 17850 9476 17850 0 _0280_
rlabel metal1 11316 17170 11316 17170 0 _0281_
rlabel metal1 12466 16728 12466 16728 0 _0282_
rlabel metal1 10994 17034 10994 17034 0 _0283_
rlabel metal1 9384 18394 9384 18394 0 _0284_
rlabel metal1 8878 19822 8878 19822 0 _0285_
rlabel metal1 9430 17068 9430 17068 0 _0286_
rlabel metal1 9522 16150 9522 16150 0 _0287_
rlabel metal2 5842 14382 5842 14382 0 _0288_
rlabel metal1 10672 16626 10672 16626 0 _0289_
rlabel metal1 9614 16116 9614 16116 0 _0290_
rlabel metal1 8372 14586 8372 14586 0 _0291_
rlabel metal1 8050 14246 8050 14246 0 _0292_
rlabel metal2 7038 17374 7038 17374 0 _0293_
rlabel metal1 7406 18054 7406 18054 0 _0294_
rlabel metal1 7958 18088 7958 18088 0 _0295_
rlabel metal1 8272 18394 8272 18394 0 _0296_
rlabel metal1 7176 18394 7176 18394 0 _0297_
rlabel metal1 5520 17714 5520 17714 0 _0298_
rlabel metal1 6348 17306 6348 17306 0 _0299_
rlabel metal1 6394 17850 6394 17850 0 _0300_
rlabel metal1 5336 17306 5336 17306 0 _0301_
rlabel metal1 5428 17102 5428 17102 0 _0302_
rlabel metal2 5014 17408 5014 17408 0 _0303_
rlabel metal2 5014 18224 5014 18224 0 _0304_
rlabel metal1 4140 18734 4140 18734 0 _0305_
rlabel metal1 7268 14858 7268 14858 0 _0306_
rlabel metal2 20102 18632 20102 18632 0 _0307_
rlabel metal1 6946 15504 6946 15504 0 _0308_
rlabel metal1 4922 15402 4922 15402 0 _0309_
rlabel metal1 6072 14586 6072 14586 0 _0310_
rlabel metal1 5566 15606 5566 15606 0 _0311_
rlabel metal1 5014 15436 5014 15436 0 _0312_
rlabel metal1 8180 14042 8180 14042 0 _0313_
rlabel metal1 7176 14042 7176 14042 0 _0314_
rlabel metal1 5704 14042 5704 14042 0 _0315_
rlabel metal1 5244 14518 5244 14518 0 _0316_
rlabel metal1 5750 12954 5750 12954 0 _0317_
rlabel metal1 6410 13226 6410 13226 0 _0318_
rlabel metal1 7406 12852 7406 12852 0 _0319_
rlabel metal2 12650 11424 12650 11424 0 _0320_
rlabel metal1 9614 10608 9614 10608 0 _0321_
rlabel metal1 9062 10676 9062 10676 0 _0322_
rlabel metal1 7314 11662 7314 11662 0 _0323_
rlabel metal1 7540 11866 7540 11866 0 _0324_
rlabel metal1 8050 11866 8050 11866 0 _0325_
rlabel metal1 7498 12784 7498 12784 0 _0326_
rlabel metal1 6440 10778 6440 10778 0 _0327_
rlabel metal1 6440 11662 6440 11662 0 _0328_
rlabel metal1 6218 12070 6218 12070 0 _0329_
rlabel metal2 6854 11900 6854 11900 0 _0330_
rlabel metal1 5842 11866 5842 11866 0 _0331_
rlabel metal1 3634 11152 3634 11152 0 _0332_
rlabel metal1 8280 9418 8280 9418 0 _0333_
rlabel metal1 8464 10030 8464 10030 0 _0334_
rlabel metal1 5842 9588 5842 9588 0 _0335_
rlabel metal1 7958 8534 7958 8534 0 _0336_
rlabel metal1 6348 8262 6348 8262 0 _0337_
rlabel metal1 6026 9146 6026 9146 0 _0338_
rlabel metal2 5750 9724 5750 9724 0 _0339_
rlabel metal1 6624 8058 6624 8058 0 _0340_
rlabel metal1 6762 8466 6762 8466 0 _0341_
rlabel metal1 9200 10234 9200 10234 0 _0342_
rlabel metal1 7452 8466 7452 8466 0 _0343_
rlabel metal1 12627 8874 12627 8874 0 _0344_
rlabel metal1 9706 9044 9706 9044 0 _0345_
rlabel metal1 11178 8500 11178 8500 0 _0346_
rlabel metal1 12236 10030 12236 10030 0 _0347_
rlabel metal1 11178 8398 11178 8398 0 _0348_
rlabel metal1 10810 8364 10810 8364 0 _0349_
rlabel metal1 9292 6834 9292 6834 0 _0350_
rlabel metal1 8648 6970 8648 6970 0 _0351_
rlabel metal1 12742 8976 12742 8976 0 _0352_
rlabel metal1 12558 9996 12558 9996 0 _0353_
rlabel metal1 12985 8874 12985 8874 0 _0354_
rlabel metal1 12604 7922 12604 7922 0 _0355_
rlabel metal1 12052 6766 12052 6766 0 _0356_
rlabel metal1 13616 11730 13616 11730 0 _0357_
rlabel metal1 13294 11866 13294 11866 0 _0358_
rlabel metal1 12328 12274 12328 12274 0 _0359_
rlabel metal1 13294 12104 13294 12104 0 _0360_
rlabel metal1 13018 13158 13018 13158 0 _0361_
rlabel metal1 12466 13226 12466 13226 0 _0362_
rlabel metal1 10304 12410 10304 12410 0 _0363_
rlabel metal1 10580 12954 10580 12954 0 _0364_
rlabel metal1 13478 12852 13478 12852 0 _0365_
rlabel metal1 10626 13260 10626 13260 0 _0366_
rlabel metal1 20424 9486 20424 9486 0 _0367_
rlabel metal1 18162 12070 18162 12070 0 _0368_
rlabel metal1 17618 13294 17618 13294 0 _0369_
rlabel metal1 16422 14450 16422 14450 0 _0370_
rlabel metal1 15042 14994 15042 14994 0 _0371_
rlabel metal1 15594 14926 15594 14926 0 _0372_
rlabel metal1 15548 13498 15548 13498 0 _0373_
rlabel metal1 15410 14042 15410 14042 0 _0374_
rlabel metal1 15548 12954 15548 12954 0 _0375_
rlabel metal1 14490 15130 14490 15130 0 _0376_
rlabel metal1 12466 15028 12466 15028 0 _0377_
rlabel metal1 17480 14586 17480 14586 0 _0378_
rlabel metal1 16744 14450 16744 14450 0 _0379_
rlabel metal1 15464 13158 15464 13158 0 _0380_
rlabel metal1 16054 13498 16054 13498 0 _0381_
rlabel metal1 16698 14586 16698 14586 0 _0382_
rlabel metal1 15548 15470 15548 15470 0 _0383_
rlabel metal1 19734 11628 19734 11628 0 _0384_
rlabel metal1 19182 12750 19182 12750 0 _0385_
rlabel metal1 18170 13362 18170 13362 0 _0386_
rlabel metal1 19149 12886 19149 12886 0 _0387_
rlabel metal1 18722 12954 18722 12954 0 _0388_
rlabel metal1 18998 15130 18998 15130 0 _0389_
rlabel metal1 16744 12342 16744 12342 0 _0390_
rlabel metal2 16330 11594 16330 11594 0 _0391_
rlabel metal1 18814 11322 18814 11322 0 _0392_
rlabel metal1 16422 11084 16422 11084 0 _0393_
rlabel via1 19450 8806 19450 8806 0 _0394_
rlabel metal1 17710 9078 17710 9078 0 _0395_
rlabel metal1 16330 8398 16330 8398 0 _0396_
rlabel metal1 16192 8602 16192 8602 0 _0397_
rlabel metal1 18078 10030 18078 10030 0 _0398_
rlabel metal1 16882 9996 16882 9996 0 _0399_
rlabel metal1 16422 9996 16422 9996 0 _0400_
rlabel metal1 15548 9622 15548 9622 0 _0401_
rlabel metal1 18262 8976 18262 8976 0 _0402_
rlabel metal1 17526 7820 17526 7820 0 _0403_
rlabel metal1 18446 10098 18446 10098 0 _0404_
rlabel metal1 17664 7854 17664 7854 0 _0405_
rlabel metal1 21896 10438 21896 10438 0 _0406_
rlabel metal1 21482 10472 21482 10472 0 _0407_
rlabel metal1 20370 10778 20370 10778 0 _0408_
rlabel metal2 19918 8177 19918 8177 0 _0409_
rlabel metal1 20470 10030 20470 10030 0 _0410_
rlabel metal1 20332 8466 20332 8466 0 _0411_
rlabel metal1 19964 8466 19964 8466 0 _0412_
rlabel metal2 20010 8058 20010 8058 0 _0413_
rlabel metal1 21352 10778 21352 10778 0 _0414_
rlabel metal2 21666 10234 21666 10234 0 _0415_
rlabel metal1 20286 10098 20286 10098 0 _0416_
rlabel metal1 21758 9996 21758 9996 0 _0417_
rlabel metal1 22770 11322 22770 11322 0 _0418_
rlabel metal1 22862 10676 22862 10676 0 _0419_
rlabel metal2 23506 9724 23506 9724 0 _0420_
rlabel metal1 25484 10030 25484 10030 0 _0421_
rlabel metal1 25438 12818 25438 12818 0 _0422_
rlabel metal1 25208 12614 25208 12614 0 _0423_
rlabel metal2 25162 10234 25162 10234 0 _0424_
rlabel metal1 24886 10030 24886 10030 0 _0425_
rlabel metal1 24794 10098 24794 10098 0 _0426_
rlabel metal1 23644 8942 23644 8942 0 _0427_
rlabel metal1 25316 12138 25316 12138 0 _0428_
rlabel metal1 25438 11730 25438 11730 0 _0429_
rlabel metal1 23092 11662 23092 11662 0 _0430_
rlabel metal1 25714 11730 25714 11730 0 _0431_
rlabel metal2 22494 13260 22494 13260 0 _0432_
rlabel metal1 22678 12886 22678 12886 0 _0433_
rlabel metal1 25438 14450 25438 14450 0 _0434_
rlabel metal1 25300 13362 25300 13362 0 _0435_
rlabel metal1 22609 13226 22609 13226 0 _0436_
rlabel metal1 21620 12954 21620 12954 0 _0437_
rlabel metal1 20838 12818 20838 12818 0 _0438_
rlabel metal1 22218 14416 22218 14416 0 _0439_
rlabel metal1 23805 14314 23805 14314 0 _0440_
rlabel metal2 22126 14756 22126 14756 0 _0441_
rlabel metal1 21942 15130 21942 15130 0 _0442_
rlabel metal1 25806 16592 25806 16592 0 _0443_
rlabel metal1 24748 15878 24748 15878 0 _0444_
rlabel metal1 25221 16218 25221 16218 0 _0445_
rlabel metal2 24978 16558 24978 16558 0 _0446_
rlabel metal1 20930 15878 20930 15878 0 _0447_
rlabel metal1 22632 16218 22632 16218 0 _0448_
rlabel metal1 23782 16218 23782 16218 0 _0449_
rlabel metal2 24150 16966 24150 16966 0 _0450_
rlabel metal2 22402 16762 22402 16762 0 _0451_
rlabel via1 22691 16558 22691 16558 0 _0452_
rlabel metal2 22218 16796 22218 16796 0 _0453_
rlabel metal2 22586 17782 22586 17782 0 _0454_
rlabel metal1 20102 17714 20102 17714 0 _0455_
rlabel metal1 19734 16660 19734 16660 0 _0456_
rlabel metal2 20562 16388 20562 16388 0 _0457_
rlabel metal1 19826 16626 19826 16626 0 _0458_
rlabel metal2 16882 17748 16882 17748 0 _0459_
rlabel metal2 17526 17612 17526 17612 0 _0460_
rlabel metal1 16882 17306 16882 17306 0 _0461_
rlabel metal1 17204 23494 17204 23494 0 _0462_
rlabel metal1 17158 22202 17158 22202 0 _0463_
rlabel metal2 18814 22372 18814 22372 0 _0464_
rlabel metal2 26174 21046 26174 21046 0 _0465_
rlabel metal1 22678 21556 22678 21556 0 _0466_
rlabel metal1 19872 21590 19872 21590 0 _0467_
rlabel metal1 20332 21522 20332 21522 0 _0468_
rlabel metal1 20286 21658 20286 21658 0 _0469_
rlabel viali 22051 21522 22051 21522 0 _0470_
rlabel metal1 21942 21046 21942 21046 0 _0471_
rlabel metal1 25776 20978 25776 20978 0 _0472_
rlabel metal1 26726 20876 26726 20876 0 _0473_
rlabel metal1 26082 21658 26082 21658 0 _0474_
rlabel metal1 25990 22474 25990 22474 0 _0475_
rlabel metal2 25898 22916 25898 22916 0 _0476_
rlabel metal1 19182 22576 19182 22576 0 _0477_
rlabel metal1 24288 23086 24288 23086 0 _0478_
rlabel metal1 23276 23630 23276 23630 0 _0479_
rlabel metal1 23184 23222 23184 23222 0 _0480_
rlabel metal1 18998 23630 18998 23630 0 _0481_
rlabel metal1 23828 22066 23828 22066 0 _0482_
rlabel metal1 18630 23766 18630 23766 0 _0483_
rlabel metal1 23736 23290 23736 23290 0 _0484_
rlabel metal1 16054 22100 16054 22100 0 _0485_
rlabel metal1 18906 25466 18906 25466 0 _0486_
rlabel metal1 17664 23698 17664 23698 0 _0487_
rlabel metal1 23690 23630 23690 23630 0 _0488_
rlabel metal1 23552 23086 23552 23086 0 _0489_
rlabel metal1 24610 23120 24610 23120 0 _0490_
rlabel metal1 25346 23290 25346 23290 0 _0491_
rlabel metal1 20838 24752 20838 24752 0 _0492_
rlabel metal2 24978 24004 24978 24004 0 _0493_
rlabel metal1 20470 24752 20470 24752 0 _0494_
rlabel metal1 26450 20944 26450 20944 0 _0495_
rlabel metal1 25024 21114 25024 21114 0 _0496_
rlabel metal1 24288 23494 24288 23494 0 _0497_
rlabel metal1 24380 21658 24380 21658 0 _0498_
rlabel metal1 24610 21862 24610 21862 0 _0499_
rlabel metal1 23736 22202 23736 22202 0 _0500_
rlabel metal1 18354 22576 18354 22576 0 _0501_
rlabel metal1 22540 24242 22540 24242 0 _0502_
rlabel metal1 21390 22542 21390 22542 0 _0503_
rlabel metal1 21574 21658 21574 21658 0 _0504_
rlabel metal1 22678 22678 22678 22678 0 _0505_
rlabel metal1 21804 22066 21804 22066 0 _0506_
rlabel metal1 21718 22616 21718 22616 0 _0507_
rlabel metal1 21666 22746 21666 22746 0 _0508_
rlabel metal2 21850 24582 21850 24582 0 _0509_
rlabel metal1 22540 24378 22540 24378 0 _0510_
rlabel metal1 20746 24310 20746 24310 0 _0511_
rlabel metal1 19688 23154 19688 23154 0 _0512_
rlabel metal1 20838 22712 20838 22712 0 _0513_
rlabel metal2 21022 21760 21022 21760 0 _0514_
rlabel metal1 20608 22202 20608 22202 0 _0515_
rlabel metal1 21252 22746 21252 22746 0 _0516_
rlabel metal1 20608 24378 20608 24378 0 _0517_
rlabel metal1 19412 23630 19412 23630 0 _0518_
rlabel metal1 18446 22746 18446 22746 0 _0519_
rlabel metal1 18860 22746 18860 22746 0 _0520_
rlabel metal1 18998 23732 18998 23732 0 _0521_
rlabel metal1 19182 23834 19182 23834 0 _0522_
rlabel metal1 18722 24208 18722 24208 0 _0523_
rlabel metal2 6762 22406 6762 22406 0 _0524_
rlabel metal2 15410 23970 15410 23970 0 _0525_
rlabel metal1 15226 21862 15226 21862 0 _0526_
rlabel metal1 14904 24106 14904 24106 0 _0527_
rlabel metal1 13386 24208 13386 24208 0 _0528_
rlabel metal1 13064 23834 13064 23834 0 _0529_
rlabel metal1 17802 22950 17802 22950 0 _0530_
rlabel metal1 20148 20434 20148 20434 0 _0531_
rlabel metal1 13018 22576 13018 22576 0 _0532_
rlabel metal1 14306 24106 14306 24106 0 _0533_
rlabel metal1 19734 25262 19734 25262 0 _0534_
rlabel metal1 16146 16558 16146 16558 0 _0535_
rlabel metal1 12742 14960 12742 14960 0 _0536_
rlabel metal1 18722 20910 18722 20910 0 _0537_
rlabel metal1 9476 22066 9476 22066 0 _0538_
rlabel metal1 9108 20774 9108 20774 0 _0539_
rlabel metal1 5014 22406 5014 22406 0 _0540_
rlabel metal1 6578 21590 6578 21590 0 _0541_
rlabel metal2 15594 18122 15594 18122 0 clknet_0_clock
rlabel metal1 14122 10166 14122 10166 0 clknet_2_0__leaf_clock
rlabel metal1 12236 23086 12236 23086 0 clknet_2_1__leaf_clock
rlabel metal1 21252 14586 21252 14586 0 clknet_2_2__leaf_clock
rlabel metal2 18446 25024 18446 25024 0 clknet_2_3__leaf_clock
rlabel metal3 2062 25228 2062 25228 0 clock
rlabel metal1 12420 29274 12420 29274 0 clock_o
rlabel metal1 5290 21114 5290 21114 0 manchester_baby_instance.BASE_0.s_countReg\[0\]
rlabel metal2 5198 22372 5198 22372 0 manchester_baby_instance.BASE_0.s_countReg\[1\]
rlabel metal1 7222 21896 7222 21896 0 manchester_baby_instance.BASE_0.s_countReg\[2\]
rlabel metal1 7222 22542 7222 22542 0 manchester_baby_instance.BASE_0.s_tickNext
rlabel metal1 8970 21046 8970 21046 0 manchester_baby_instance.BASE_0.s_tickReg
rlabel metal1 11546 23154 11546 23154 0 manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
rlabel metal1 9706 21658 9706 21658 0 manchester_baby_instance.BASE_1.s_counterValue
rlabel metal2 11638 22372 11638 22372 0 manchester_baby_instance.BASE_1.s_derivedClock
rlabel metal1 20240 24174 20240 24174 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
rlabel metal2 21390 24616 21390 24616 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
rlabel metal1 23000 20842 23000 20842 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
rlabel metal2 24196 24786 24196 24786 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
rlabel metal1 25070 21590 25070 21590 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
rlabel metal2 17986 23494 17986 23494 0 manchester_baby_instance.CIRCUIT_0.Acc.tick
rlabel metal1 15226 24718 15226 24718 0 manchester_baby_instance.CIRCUIT_0.GATES_13.result
rlabel metal1 19274 20978 19274 20978 0 manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
rlabel metal2 15686 19074 15686 19074 0 manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
rlabel metal2 16330 22100 16330 22100 0 manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
rlabel metal1 17066 21998 17066 21998 0 manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
rlabel metal2 21022 20128 21022 20128 0 manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
rlabel metal1 22632 20026 22632 20026 0 manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
rlabel metal1 26312 19482 26312 19482 0 manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
rlabel metal1 24656 20366 24656 20366 0 manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
rlabel metal1 17802 24174 17802 24174 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
rlabel metal1 17342 24208 17342 24208 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
rlabel metal1 17158 24174 17158 24174 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
rlabel metal1 16192 24378 16192 24378 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
rlabel metal1 14812 25330 14812 25330 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
rlabel metal1 12926 24378 12926 24378 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
rlabel metal1 30314 16456 30314 16456 0 net1
rlabel metal1 13156 8466 13156 8466 0 net10
rlabel metal1 18768 20570 18768 20570 0 net100
rlabel metal1 26450 11730 26450 11730 0 net101
rlabel metal1 6210 18700 6210 18700 0 net102
rlabel metal1 22632 19482 22632 19482 0 net103
rlabel metal2 11914 18938 11914 18938 0 net104
rlabel metal1 25484 20570 25484 20570 0 net105
rlabel metal1 20148 18666 20148 18666 0 net106
rlabel metal1 25254 18666 25254 18666 0 net107
rlabel metal1 20148 16558 20148 16558 0 net108
rlabel metal1 10074 9078 10074 9078 0 net11
rlabel metal1 21022 22678 21022 22678 0 net12
rlabel metal1 1610 7480 1610 7480 0 net13
rlabel metal1 5980 8942 5980 8942 0 net14
rlabel metal1 6670 12818 6670 12818 0 net15
rlabel metal2 7038 13056 7038 13056 0 net16
rlabel metal1 5566 13974 5566 13974 0 net17
rlabel metal1 5750 15402 5750 15402 0 net18
rlabel metal1 2990 19482 2990 19482 0 net19
rlabel metal1 17802 2618 17802 2618 0 net2
rlabel metal1 4324 23562 4324 23562 0 net20
rlabel metal1 6762 18836 6762 18836 0 net21
rlabel metal1 2231 19754 2231 19754 0 net22
rlabel metal1 21666 20876 21666 20876 0 net23
rlabel metal1 12650 18054 12650 18054 0 net24
rlabel metal1 12788 29002 12788 29002 0 net25
rlabel metal1 26358 20468 26358 20468 0 net26
rlabel metal1 25484 20502 25484 20502 0 net27
rlabel metal1 26358 13430 26358 13430 0 net28
rlabel metal1 23506 11084 23506 11084 0 net29
rlabel metal1 17112 2618 17112 2618 0 net3
rlabel metal1 27048 10710 27048 10710 0 net30
rlabel metal1 21896 9554 21896 9554 0 net31
rlabel metal1 21528 2618 21528 2618 0 net32
rlabel metal2 1702 16932 1702 16932 0 net33
rlabel metal1 13248 23562 13248 23562 0 net34
rlabel metal1 19504 21658 19504 21658 0 net35
rlabel metal1 20700 20570 20700 20570 0 net36
rlabel metal1 27462 19822 27462 19822 0 net37
rlabel metal1 30222 20978 30222 20978 0 net38
rlabel metal2 25070 21828 25070 21828 0 net39
rlabel metal2 18998 2689 18998 2689 0 net4
rlabel metal2 19366 23494 19366 23494 0 net40
rlabel metal1 18308 7854 18308 7854 0 net41
rlabel metal1 15548 8942 15548 8942 0 net42
rlabel metal2 16514 2587 16514 2587 0 net43
rlabel metal1 19090 14416 19090 14416 0 net44
rlabel metal1 17066 15572 17066 15572 0 net45
rlabel metal1 1702 14348 1702 14348 0 net46
rlabel metal1 1702 11084 1702 11084 0 net47
rlabel metal1 13064 13294 13064 13294 0 net48
rlabel metal1 12604 7718 12604 7718 0 net49
rlabel metal1 18400 14518 18400 14518 0 net5
rlabel metal1 10396 7174 10396 7174 0 net50
rlabel metal1 20010 18156 20010 18156 0 net51
rlabel metal1 1702 7888 1702 7888 0 net52
rlabel metal1 4968 10030 4968 10030 0 net53
rlabel metal1 4646 11526 4646 11526 0 net54
rlabel metal1 2231 12818 2231 12818 0 net55
rlabel metal1 2484 13702 2484 13702 0 net56
rlabel metal1 1702 16048 1702 16048 0 net57
rlabel metal1 3082 22610 3082 22610 0 net58
rlabel metal2 1702 21658 1702 21658 0 net59
rlabel metal1 15686 2550 15686 2550 0 net6
rlabel metal1 10074 16014 10074 16014 0 net60
rlabel metal1 1702 20842 1702 20842 0 net61
rlabel metal1 24242 18598 24242 18598 0 net62
rlabel metal1 1702 21454 1702 21454 0 net63
rlabel metal1 19734 23800 19734 23800 0 net64
rlabel metal2 27370 17408 27370 17408 0 net65
rlabel metal1 30222 15402 30222 15402 0 net66
rlabel metal2 21298 13192 21298 13192 0 net67
rlabel metal1 27416 11322 27416 11322 0 net68
rlabel metal2 25622 9214 25622 9214 0 net69
rlabel metal1 14950 19890 14950 19890 0 net7
rlabel metal1 26910 8398 26910 8398 0 net70
rlabel metal1 20930 7174 20930 7174 0 net71
rlabel metal2 15686 25398 15686 25398 0 net72
rlabel metal1 14076 23766 14076 23766 0 net73
rlabel metal1 23874 16660 23874 16660 0 net74
rlabel metal2 26450 17612 26450 17612 0 net75
rlabel metal1 12052 23290 12052 23290 0 net76
rlabel metal1 10104 23018 10104 23018 0 net77
rlabel metal1 5566 22610 5566 22610 0 net78
rlabel metal1 7360 22610 7360 22610 0 net79
rlabel metal1 11500 2618 11500 2618 0 net8
rlabel via1 7033 21522 7033 21522 0 net80
rlabel metal1 5566 22406 5566 22406 0 net81
rlabel metal2 4646 21794 4646 21794 0 net82
rlabel metal1 9338 22202 9338 22202 0 net83
rlabel metal1 9890 21454 9890 21454 0 net84
rlabel metal1 14214 21454 14214 21454 0 net85
rlabel metal1 12643 22202 12643 22202 0 net86
rlabel via1 5290 15453 5290 15453 0 net87
rlabel metal1 20424 7854 20424 7854 0 net88
rlabel metal1 5198 14892 5198 14892 0 net89
rlabel metal1 13938 2618 13938 2618 0 net9
rlabel via1 7673 8466 7673 8466 0 net90
rlabel metal1 7774 12886 7774 12886 0 net91
rlabel metal1 5474 9588 5474 9588 0 net92
rlabel metal1 24426 8942 24426 8942 0 net93
rlabel metal1 10120 16082 10120 16082 0 net94
rlabel metal2 22402 9860 22402 9860 0 net95
rlabel metal1 26036 17170 26036 17170 0 net96
rlabel metal1 16606 11118 16606 11118 0 net97
rlabel metal1 22586 24752 22586 24752 0 net98
rlabel metal1 10994 13294 10994 13294 0 net99
rlabel metal1 19826 29274 19826 29274 0 ram_addr_o[0]
rlabel metal1 20792 29274 20792 29274 0 ram_addr_o[1]
rlabel metal2 30406 19873 30406 19873 0 ram_addr_o[2]
rlabel metal1 30360 20774 30360 20774 0 ram_addr_o[3]
rlabel metal2 30406 21505 30406 21505 0 ram_addr_o[4]
rlabel metal1 30728 16558 30728 16558 0 ram_data_i[0]
rlabel metal2 17434 959 17434 959 0 ram_data_i[10]
rlabel metal2 16790 959 16790 959 0 ram_data_i[11]
rlabel metal2 18722 1588 18722 1588 0 ram_data_i[12]
rlabel metal1 30360 12818 30360 12818 0 ram_data_i[13]
rlabel metal2 14858 1554 14858 1554 0 ram_data_i[14]
rlabel metal1 14950 29206 14950 29206 0 ram_data_i[15]
rlabel metal2 11638 1027 11638 1027 0 ram_data_i[16]
rlabel metal2 13570 1027 13570 1027 0 ram_data_i[17]
rlabel metal2 9062 1027 9062 1027 0 ram_data_i[18]
rlabel metal2 9706 1027 9706 1027 0 ram_data_i[19]
rlabel metal1 30728 22610 30728 22610 0 ram_data_i[1]
rlabel metal3 1050 6868 1050 6868 0 ram_data_i[20]
rlabel metal3 1050 8228 1050 8228 0 ram_data_i[21]
rlabel metal3 820 8908 820 8908 0 ram_data_i[22]
rlabel metal3 820 11628 820 11628 0 ram_data_i[23]
rlabel metal3 1050 13668 1050 13668 0 ram_data_i[24]
rlabel metal3 1050 15028 1050 15028 0 ram_data_i[25]
rlabel metal3 751 19108 751 19108 0 ram_data_i[26]
rlabel metal3 751 23188 751 23188 0 ram_data_i[27]
rlabel metal3 751 17748 751 17748 0 ram_data_i[28]
rlabel metal3 820 19788 820 19788 0 ram_data_i[29]
rlabel metal1 30360 19346 30360 19346 0 ram_data_i[2]
rlabel metal3 820 18428 820 18428 0 ram_data_i[30]
rlabel metal1 13156 29138 13156 29138 0 ram_data_i[31]
rlabel metal2 30498 21675 30498 21675 0 ram_data_i[3]
rlabel metal1 30360 23698 30360 23698 0 ram_data_i[4]
rlabel metal1 30498 13872 30498 13872 0 ram_data_i[5]
rlabel metal1 30406 11118 30406 11118 0 ram_data_i[6]
rlabel metal1 30728 10642 30728 10642 0 ram_data_i[7]
rlabel metal1 30406 10030 30406 10030 0 ram_data_i[8]
rlabel metal2 21298 1588 21298 1588 0 ram_data_i[9]
rlabel metal1 19090 29274 19090 29274 0 ram_data_o[0]
rlabel metal2 18078 1520 18078 1520 0 ram_data_o[10]
rlabel metal2 15502 959 15502 959 0 ram_data_o[11]
rlabel metal2 16146 959 16146 959 0 ram_data_o[12]
rlabel metal2 30406 14433 30406 14433 0 ram_data_o[13]
rlabel metal2 30406 15793 30406 15793 0 ram_data_o[14]
rlabel metal3 820 14348 820 14348 0 ram_data_o[15]
rlabel metal3 1096 10948 1096 10948 0 ram_data_o[16]
rlabel metal2 12926 959 12926 959 0 ram_data_o[17]
rlabel metal2 12282 1520 12282 1520 0 ram_data_o[18]
rlabel metal2 10350 1520 10350 1520 0 ram_data_o[19]
rlabel metal1 30360 18054 30360 18054 0 ram_data_o[1]
rlabel metal3 820 7548 820 7548 0 ram_data_o[20]
rlabel metal3 1096 9588 1096 9588 0 ram_data_o[21]
rlabel metal3 820 10268 820 10268 0 ram_data_o[22]
rlabel metal3 1096 12308 1096 12308 0 ram_data_o[23]
rlabel metal3 820 12988 820 12988 0 ram_data_o[24]
rlabel metal3 820 15708 820 15708 0 ram_data_o[25]
rlabel metal3 820 22508 820 22508 0 ram_data_o[26]
rlabel metal3 820 21828 820 21828 0 ram_data_o[27]
rlabel metal1 1242 16422 1242 16422 0 ram_data_o[28]
rlabel metal3 751 20468 751 20468 0 ram_data_o[29]
rlabel metal2 30406 18513 30406 18513 0 ram_data_o[2]
rlabel metal3 820 21148 820 21148 0 ram_data_o[30]
rlabel metal2 21942 30304 21942 30304 0 ram_data_o[31]
rlabel via2 30406 17051 30406 17051 0 ram_data_o[3]
rlabel metal1 30360 15334 30360 15334 0 ram_data_o[4]
rlabel metal2 30406 13073 30406 13073 0 ram_data_o[5]
rlabel via2 30406 11611 30406 11611 0 ram_data_o[6]
rlabel metal2 30406 9027 30406 9027 0 ram_data_o[7]
rlabel metal1 30360 8330 30360 8330 0 ram_data_o[8]
rlabel metal2 20654 1520 20654 1520 0 ram_data_o[9]
rlabel metal2 15778 30311 15778 30311 0 ram_rw_en_o
rlabel metal3 820 17068 820 17068 0 reset_i
rlabel metal1 14352 29274 14352 29274 0 stop_lamp_o
<< properties >>
string FIXED_BBOX 0 0 32000 32000
<< end >>
