magic
tech sky130A
magscale 1 2
timestamp 1700142110
<< viali >>
rect 15761 37417 15795 37451
rect 17693 37417 17727 37451
rect 19625 37417 19659 37451
rect 22109 37417 22143 37451
rect 15669 37145 15703 37179
rect 17601 37145 17635 37179
rect 19533 37145 19567 37179
rect 22385 37145 22419 37179
rect 7573 31229 7607 31263
rect 8217 31093 8251 31127
rect 7297 30889 7331 30923
rect 6837 30753 6871 30787
rect 7389 30753 7423 30787
rect 8125 30753 8159 30787
rect 6745 30685 6779 30719
rect 7113 30685 7147 30719
rect 7205 30685 7239 30719
rect 7481 30685 7515 30719
rect 8217 30685 8251 30719
rect 8401 30685 8435 30719
rect 10609 30685 10643 30719
rect 11805 30685 11839 30719
rect 12265 30685 12299 30719
rect 16957 30685 16991 30719
rect 6377 30549 6411 30583
rect 8401 30549 8435 30583
rect 10793 30549 10827 30583
rect 11253 30549 11287 30583
rect 12909 30549 12943 30583
rect 17601 30549 17635 30583
rect 7481 30345 7515 30379
rect 10793 30345 10827 30379
rect 11345 30345 11379 30379
rect 8594 30277 8628 30311
rect 10333 30277 10367 30311
rect 6561 30209 6595 30243
rect 8861 30209 8895 30243
rect 10885 30209 10919 30243
rect 13165 30209 13199 30243
rect 15761 30209 15795 30243
rect 19605 30209 19639 30243
rect 12449 30141 12483 30175
rect 12909 30141 12943 30175
rect 19349 30141 19383 30175
rect 20913 30141 20947 30175
rect 10701 30073 10735 30107
rect 14289 30073 14323 30107
rect 20729 30073 20763 30107
rect 7205 30005 7239 30039
rect 11161 30005 11195 30039
rect 11897 30005 11931 30039
rect 15669 30005 15703 30039
rect 21557 30005 21591 30039
rect 11989 29801 12023 29835
rect 12633 29801 12667 29835
rect 7849 29733 7883 29767
rect 20269 29733 20303 29767
rect 7665 29665 7699 29699
rect 12265 29665 12299 29699
rect 14473 29665 14507 29699
rect 16589 29665 16623 29699
rect 20177 29665 20211 29699
rect 20637 29665 20671 29699
rect 5825 29597 5859 29631
rect 6009 29597 6043 29631
rect 6193 29597 6227 29631
rect 7398 29597 7432 29631
rect 7757 29597 7791 29631
rect 8033 29597 8067 29631
rect 8953 29597 8987 29631
rect 9137 29597 9171 29631
rect 10609 29597 10643 29631
rect 10876 29597 10910 29631
rect 12357 29597 12391 29631
rect 13277 29597 13311 29631
rect 19901 29597 19935 29631
rect 20821 29597 20855 29631
rect 21088 29597 21122 29631
rect 8493 29529 8527 29563
rect 14749 29529 14783 29563
rect 16497 29529 16531 29563
rect 16865 29529 16899 29563
rect 18613 29529 18647 29563
rect 5273 29461 5307 29495
rect 6009 29461 6043 29495
rect 6285 29461 6319 29495
rect 9045 29461 9079 29495
rect 13369 29461 13403 29495
rect 20085 29461 20119 29495
rect 22201 29461 22235 29495
rect 4813 29257 4847 29291
rect 9689 29257 9723 29291
rect 11161 29257 11195 29291
rect 15025 29257 15059 29291
rect 16773 29257 16807 29291
rect 17693 29257 17727 29291
rect 15393 29189 15427 29223
rect 5937 29121 5971 29155
rect 6193 29121 6227 29155
rect 7113 29121 7147 29155
rect 8309 29121 8343 29155
rect 8576 29121 8610 29155
rect 9781 29121 9815 29155
rect 10048 29121 10082 29155
rect 15209 29121 15243 29155
rect 15301 29121 15335 29155
rect 15577 29121 15611 29155
rect 16957 29121 16991 29155
rect 17049 29121 17083 29155
rect 17141 29121 17175 29155
rect 17325 29121 17359 29155
rect 17601 29121 17635 29155
rect 18245 29121 18279 29155
rect 6377 29053 6411 29087
rect 6929 29053 6963 29087
rect 7389 29053 7423 29087
rect 8033 29053 8067 29087
rect 12357 29053 12391 29087
rect 12633 29053 12667 29087
rect 14105 29053 14139 29087
rect 14841 29053 14875 29087
rect 20269 29053 20303 29087
rect 7205 28985 7239 29019
rect 7297 28917 7331 28951
rect 7481 28917 7515 28951
rect 14289 28917 14323 28951
rect 18502 28917 18536 28951
rect 5365 28713 5399 28747
rect 7757 28713 7791 28747
rect 8953 28713 8987 28747
rect 12817 28713 12851 28747
rect 18245 28713 18279 28747
rect 19349 28713 19383 28747
rect 5825 28645 5859 28679
rect 8677 28645 8711 28679
rect 5135 28577 5169 28611
rect 5696 28577 5730 28611
rect 5917 28577 5951 28611
rect 6101 28577 6135 28611
rect 6377 28577 6411 28611
rect 9505 28577 9539 28611
rect 12357 28577 12391 28611
rect 16405 28577 16439 28611
rect 16681 28577 16715 28611
rect 4997 28509 5031 28543
rect 5273 28509 5307 28543
rect 5457 28509 5491 28543
rect 8585 28509 8619 28543
rect 8769 28509 8803 28543
rect 9689 28509 9723 28543
rect 9873 28509 9907 28543
rect 12633 28509 12667 28543
rect 13001 28509 13035 28543
rect 13093 28509 13127 28543
rect 13369 28509 13403 28543
rect 16313 28509 16347 28543
rect 18429 28509 18463 28543
rect 18797 28509 18831 28543
rect 19257 28509 19291 28543
rect 20361 28509 20395 28543
rect 20617 28509 20651 28543
rect 5549 28441 5583 28475
rect 6644 28441 6678 28475
rect 10333 28441 10367 28475
rect 12081 28441 12115 28475
rect 13185 28441 13219 28475
rect 18521 28441 18555 28475
rect 18613 28441 18647 28475
rect 9965 28373 9999 28407
rect 12541 28373 12575 28407
rect 21741 28373 21775 28407
rect 6745 28169 6779 28203
rect 7021 28169 7055 28203
rect 9413 28169 9447 28203
rect 12909 28169 12943 28203
rect 13829 28169 13863 28203
rect 18889 28169 18923 28203
rect 19165 28169 19199 28203
rect 19809 28169 19843 28203
rect 20545 28169 20579 28203
rect 6837 28101 6871 28135
rect 13185 28101 13219 28135
rect 13277 28101 13311 28135
rect 16297 28101 16331 28135
rect 16497 28101 16531 28135
rect 18521 28101 18555 28135
rect 23029 28101 23063 28135
rect 6377 28033 6411 28067
rect 7113 28033 7147 28067
rect 8401 28033 8435 28067
rect 8585 28033 8619 28067
rect 9229 28033 9263 28067
rect 9413 28033 9447 28067
rect 9965 28033 9999 28067
rect 10241 28033 10275 28067
rect 13093 28033 13127 28067
rect 13461 28033 13495 28067
rect 14013 28033 14047 28067
rect 14197 28033 14231 28067
rect 15761 28033 15795 28067
rect 15945 28033 15979 28067
rect 16037 28033 16071 28067
rect 18429 28033 18463 28067
rect 18705 28033 18739 28067
rect 20729 28033 20763 28067
rect 20913 28033 20947 28067
rect 22569 28033 22603 28067
rect 22845 28033 22879 28067
rect 6469 27965 6503 27999
rect 9781 27965 9815 27999
rect 15025 27965 15059 27999
rect 19349 27965 19383 27999
rect 19441 27965 19475 27999
rect 21005 27965 21039 27999
rect 22017 27965 22051 27999
rect 23213 27965 23247 27999
rect 6837 27897 6871 27931
rect 14749 27897 14783 27931
rect 16129 27897 16163 27931
rect 22293 27897 22327 27931
rect 22753 27897 22787 27931
rect 6377 27829 6411 27863
rect 8493 27829 8527 27863
rect 10149 27829 10183 27863
rect 10425 27829 10459 27863
rect 14197 27829 14231 27863
rect 14565 27829 14599 27863
rect 15577 27829 15611 27863
rect 16313 27829 16347 27863
rect 22477 27829 22511 27863
rect 6377 27625 6411 27659
rect 8953 27625 8987 27659
rect 12725 27625 12759 27659
rect 12909 27625 12943 27659
rect 18705 27625 18739 27659
rect 22569 27625 22603 27659
rect 5181 27557 5215 27591
rect 12265 27557 12299 27591
rect 14105 27557 14139 27591
rect 15025 27557 15059 27591
rect 17233 27557 17267 27591
rect 5825 27489 5859 27523
rect 13277 27489 13311 27523
rect 13645 27489 13679 27523
rect 14473 27489 14507 27523
rect 19257 27489 19291 27523
rect 3801 27421 3835 27455
rect 6009 27421 6043 27455
rect 7389 27421 7423 27455
rect 7573 27421 7607 27455
rect 8401 27421 8435 27455
rect 9597 27421 9631 27455
rect 10802 27421 10836 27455
rect 11069 27421 11103 27455
rect 11989 27421 12023 27455
rect 12357 27421 12391 27455
rect 12633 27421 12667 27455
rect 13921 27421 13955 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 14565 27421 14599 27455
rect 15163 27421 15197 27455
rect 15301 27421 15335 27455
rect 15393 27421 15427 27455
rect 15521 27421 15555 27455
rect 15669 27421 15703 27455
rect 16589 27421 16623 27455
rect 16682 27421 16716 27455
rect 17054 27421 17088 27455
rect 18153 27421 18187 27455
rect 18521 27421 18555 27455
rect 18981 27421 19015 27455
rect 19441 27421 19475 27455
rect 19625 27421 19659 27455
rect 19717 27421 19751 27455
rect 20269 27421 20303 27455
rect 22293 27421 22327 27455
rect 22385 27421 22419 27455
rect 23774 27421 23808 27455
rect 24041 27421 24075 27455
rect 4068 27353 4102 27387
rect 6193 27353 6227 27387
rect 7757 27353 7791 27387
rect 12265 27353 12299 27387
rect 13160 27353 13194 27387
rect 16865 27353 16899 27387
rect 16977 27353 17011 27387
rect 18337 27353 18371 27387
rect 18429 27353 18463 27387
rect 18889 27353 18923 27387
rect 20545 27353 20579 27387
rect 5273 27285 5307 27319
rect 7389 27285 7423 27319
rect 9689 27285 9723 27319
rect 12081 27285 12115 27319
rect 13001 27285 13035 27319
rect 13369 27285 13403 27319
rect 13829 27285 13863 27319
rect 22017 27285 22051 27319
rect 22661 27285 22695 27319
rect 4169 27081 4203 27115
rect 10977 27081 11011 27115
rect 12541 27081 12575 27115
rect 13461 27081 13495 27115
rect 14105 27081 14139 27115
rect 15577 27081 15611 27115
rect 17049 27081 17083 27115
rect 17233 27081 17267 27115
rect 17969 27081 18003 27115
rect 18337 27081 18371 27115
rect 18429 27081 18463 27115
rect 20453 27081 20487 27115
rect 21373 27081 21407 27115
rect 22661 27081 22695 27115
rect 23213 27081 23247 27115
rect 15301 27013 15335 27047
rect 16707 27013 16741 27047
rect 18705 27013 18739 27047
rect 18797 27013 18831 27047
rect 19625 27013 19659 27047
rect 21005 27013 21039 27047
rect 16911 26979 16945 27013
rect 5273 26945 5307 26979
rect 5733 26945 5767 26979
rect 6009 26945 6043 26979
rect 6193 26945 6227 26979
rect 6929 26945 6963 26979
rect 7113 26945 7147 26979
rect 7297 26945 7331 26979
rect 8217 26945 8251 26979
rect 8401 26945 8435 26979
rect 8668 26945 8702 26979
rect 10609 26945 10643 26979
rect 10793 26945 10827 26979
rect 11253 26945 11287 26979
rect 11345 26945 11379 26979
rect 11805 26945 11839 26979
rect 11989 26945 12023 26979
rect 12357 26945 12391 26979
rect 12817 26945 12851 26979
rect 13645 26945 13679 26979
rect 13829 26945 13863 26979
rect 14289 26945 14323 26979
rect 15025 26945 15059 26979
rect 15209 26945 15243 26979
rect 15393 26945 15427 26979
rect 15669 26945 15703 26979
rect 15761 26945 15795 26979
rect 16129 26945 16163 26979
rect 17141 26945 17175 26979
rect 17417 26945 17451 26979
rect 17509 26945 17543 26979
rect 17693 26945 17727 26979
rect 17880 26945 17914 26979
rect 18153 26945 18187 26979
rect 18613 26945 18647 26979
rect 18981 26945 19015 26979
rect 19165 26945 19199 26979
rect 19257 26945 19291 26979
rect 20867 26945 20901 26979
rect 21281 26945 21315 26979
rect 22385 26945 22419 26979
rect 22661 26945 22695 26979
rect 22845 26945 22879 26979
rect 23029 26945 23063 26979
rect 3341 26877 3375 26911
rect 4813 26877 4847 26911
rect 4905 26877 4939 26911
rect 5365 26877 5399 26911
rect 5917 26877 5951 26911
rect 6377 26877 6411 26911
rect 7849 26877 7883 26911
rect 10425 26877 10459 26911
rect 11069 26877 11103 26911
rect 12081 26877 12115 26911
rect 12633 26877 12667 26911
rect 13001 26877 13035 26911
rect 13737 26877 13771 26911
rect 13921 26877 13955 26911
rect 14565 26877 14599 26911
rect 15945 26877 15979 26911
rect 20637 26877 20671 26911
rect 20729 26877 20763 26911
rect 21097 26877 21131 26911
rect 6009 26809 6043 26843
rect 9781 26809 9815 26843
rect 14473 26809 14507 26843
rect 17417 26809 17451 26843
rect 17509 26809 17543 26843
rect 19441 26809 19475 26843
rect 19993 26809 20027 26843
rect 21833 26809 21867 26843
rect 3985 26741 4019 26775
rect 5549 26741 5583 26775
rect 7205 26741 7239 26775
rect 9873 26741 9907 26775
rect 11161 26741 11195 26775
rect 11989 26741 12023 26775
rect 12173 26741 12207 26775
rect 16865 26741 16899 26775
rect 19625 26741 19659 26775
rect 2237 26537 2271 26571
rect 6009 26537 6043 26571
rect 8401 26537 8435 26571
rect 9413 26537 9447 26571
rect 11161 26537 11195 26571
rect 15209 26537 15243 26571
rect 16313 26537 16347 26571
rect 19257 26537 19291 26571
rect 19441 26537 19475 26571
rect 20177 26537 20211 26571
rect 21649 26537 21683 26571
rect 21833 26537 21867 26571
rect 9321 26469 9355 26503
rect 19993 26469 20027 26503
rect 22201 26469 22235 26503
rect 3617 26401 3651 26435
rect 6561 26401 6595 26435
rect 9505 26401 9539 26435
rect 10517 26401 10551 26435
rect 4445 26333 4479 26367
rect 4629 26333 4663 26367
rect 6828 26333 6862 26367
rect 8033 26333 8067 26367
rect 8953 26333 8987 26367
rect 9965 26333 9999 26367
rect 15577 26333 15611 26367
rect 16497 26333 16531 26367
rect 16957 26333 16991 26367
rect 19809 26333 19843 26367
rect 22477 26333 22511 26367
rect 23121 26333 23155 26367
rect 23305 26333 23339 26367
rect 23397 26333 23431 26367
rect 23581 26333 23615 26367
rect 28181 26333 28215 26367
rect 28457 26333 28491 26367
rect 3372 26265 3406 26299
rect 4896 26265 4930 26299
rect 8217 26265 8251 26299
rect 12633 26265 12667 26299
rect 15393 26265 15427 26299
rect 16589 26265 16623 26299
rect 16681 26265 16715 26299
rect 16819 26265 16853 26299
rect 19441 26265 19475 26299
rect 20177 26265 20211 26299
rect 20361 26265 20395 26299
rect 21833 26265 21867 26299
rect 3893 26197 3927 26231
rect 7941 26197 7975 26231
rect 9781 26197 9815 26231
rect 22385 26197 22419 26231
rect 23121 26197 23155 26231
rect 23581 26197 23615 26231
rect 29193 26197 29227 26231
rect 4353 25993 4387 26027
rect 5089 25993 5123 26027
rect 9781 25993 9815 26027
rect 11253 25993 11287 26027
rect 13829 25993 13863 26027
rect 16865 25993 16899 26027
rect 17509 25993 17543 26027
rect 18429 25993 18463 26027
rect 20637 25993 20671 26027
rect 22201 25993 22235 26027
rect 25513 25993 25547 26027
rect 12173 25925 12207 25959
rect 17785 25925 17819 25959
rect 21373 25925 21407 25959
rect 24378 25925 24412 25959
rect 2798 25857 2832 25891
rect 3525 25857 3559 25891
rect 4629 25857 4663 25891
rect 5273 25857 5307 25891
rect 5457 25857 5491 25891
rect 7297 25857 7331 25891
rect 9321 25857 9355 25891
rect 9413 25857 9447 25891
rect 9597 25857 9631 25891
rect 9873 25857 9907 25891
rect 11069 25857 11103 25891
rect 11345 25857 11379 25891
rect 11713 25857 11747 25891
rect 12357 25857 12391 25891
rect 13277 25857 13311 25891
rect 13461 25857 13495 25891
rect 13553 25857 13587 25891
rect 13645 25857 13679 25891
rect 16313 25857 16347 25891
rect 16497 25857 16531 25891
rect 17141 25857 17175 25891
rect 18153 25857 18187 25891
rect 18337 25857 18371 25891
rect 18521 25857 18555 25891
rect 18705 25857 18739 25891
rect 20545 25857 20579 25891
rect 20729 25857 20763 25891
rect 20913 25857 20947 25891
rect 21281 25857 21315 25891
rect 21465 25857 21499 25891
rect 21833 25857 21867 25891
rect 23774 25857 23808 25891
rect 24041 25857 24075 25891
rect 24133 25857 24167 25891
rect 28273 25857 28307 25891
rect 29101 25857 29135 25891
rect 29469 25857 29503 25891
rect 3065 25789 3099 25823
rect 4077 25789 4111 25823
rect 4353 25789 4387 25823
rect 5549 25789 5583 25823
rect 8677 25789 8711 25823
rect 10885 25789 10919 25823
rect 11805 25789 11839 25823
rect 12633 25789 12667 25823
rect 17049 25789 17083 25823
rect 29377 25789 29411 25823
rect 29745 25789 29779 25823
rect 7297 25721 7331 25755
rect 22661 25721 22695 25755
rect 1685 25653 1719 25687
rect 4537 25653 4571 25687
rect 9413 25653 9447 25687
rect 11989 25653 12023 25687
rect 12541 25653 12575 25687
rect 16129 25653 16163 25687
rect 17601 25653 17635 25687
rect 17785 25653 17819 25687
rect 19993 25653 20027 25687
rect 21097 25653 21131 25687
rect 22201 25653 22235 25687
rect 22385 25653 22419 25687
rect 31217 25653 31251 25687
rect 2605 25449 2639 25483
rect 3046 25449 3080 25483
rect 3525 25449 3559 25483
rect 3893 25449 3927 25483
rect 8033 25449 8067 25483
rect 10517 25449 10551 25483
rect 12817 25449 12851 25483
rect 15117 25449 15151 25483
rect 15577 25449 15611 25483
rect 16773 25449 16807 25483
rect 17325 25449 17359 25483
rect 17509 25449 17543 25483
rect 20913 25449 20947 25483
rect 22569 25449 22603 25483
rect 23397 25449 23431 25483
rect 29745 25449 29779 25483
rect 30573 25449 30607 25483
rect 3157 25381 3191 25415
rect 14381 25381 14415 25415
rect 21005 25381 21039 25415
rect 28273 25381 28307 25415
rect 3249 25313 3283 25347
rect 7849 25313 7883 25347
rect 11897 25313 11931 25347
rect 12633 25313 12667 25347
rect 14197 25313 14231 25347
rect 14841 25313 14875 25347
rect 16037 25313 16071 25347
rect 21373 25313 21407 25347
rect 22385 25313 22419 25347
rect 1869 25245 1903 25279
rect 1961 25245 1995 25279
rect 3801 25245 3835 25279
rect 3985 25245 4019 25279
rect 5273 25245 5307 25279
rect 5457 25245 5491 25279
rect 5549 25245 5583 25279
rect 7757 25245 7791 25279
rect 9137 25245 9171 25279
rect 10793 25245 10827 25279
rect 11805 25245 11839 25279
rect 12541 25245 12575 25279
rect 14473 25245 14507 25279
rect 14749 25245 14783 25279
rect 15669 25245 15703 25279
rect 15853 25245 15887 25279
rect 15945 25245 15979 25279
rect 16129 25245 16163 25279
rect 16681 25245 16715 25279
rect 16865 25245 16899 25279
rect 17141 25245 17175 25279
rect 17601 25245 17635 25279
rect 19809 25245 19843 25279
rect 20177 25245 20211 25279
rect 20269 25245 20303 25279
rect 20545 25245 20579 25279
rect 21189 25245 21223 25279
rect 22109 25245 22143 25279
rect 22477 25245 22511 25279
rect 22753 25245 22787 25279
rect 22937 25245 22971 25279
rect 23213 25245 23247 25279
rect 25421 25245 25455 25279
rect 27261 25245 27295 25279
rect 27537 25245 27571 25279
rect 29561 25245 29595 25279
rect 30481 25245 30515 25279
rect 2881 25177 2915 25211
rect 9404 25177 9438 25211
rect 14197 25177 14231 25211
rect 15209 25177 15243 25211
rect 15393 25177 15427 25211
rect 16957 25177 16991 25211
rect 19901 25177 19935 25211
rect 19993 25177 20027 25211
rect 20754 25177 20788 25211
rect 22845 25177 22879 25211
rect 23029 25177 23063 25211
rect 25697 25177 25731 25211
rect 1685 25109 1719 25143
rect 5089 25109 5123 25143
rect 11345 25109 11379 25143
rect 12173 25109 12207 25143
rect 15761 25109 15795 25143
rect 19625 25109 19659 25143
rect 20637 25109 20671 25143
rect 27169 25109 27203 25143
rect 1961 24905 1995 24939
rect 2421 24905 2455 24939
rect 6009 24905 6043 24939
rect 10793 24905 10827 24939
rect 13369 24905 13403 24939
rect 14841 24905 14875 24939
rect 20177 24905 20211 24939
rect 22201 24905 22235 24939
rect 25973 24905 26007 24939
rect 26433 24905 26467 24939
rect 27261 24905 27295 24939
rect 29653 24905 29687 24939
rect 4712 24837 4746 24871
rect 9965 24837 9999 24871
rect 13645 24837 13679 24871
rect 14289 24837 14323 24871
rect 15209 24837 15243 24871
rect 16957 24837 16991 24871
rect 17049 24837 17083 24871
rect 22109 24837 22143 24871
rect 30021 24837 30055 24871
rect 32505 24837 32539 24871
rect 1593 24769 1627 24803
rect 2329 24769 2363 24803
rect 2605 24769 2639 24803
rect 2789 24769 2823 24803
rect 4445 24769 4479 24803
rect 5917 24769 5951 24803
rect 6101 24769 6135 24803
rect 6561 24769 6595 24803
rect 7665 24769 7699 24803
rect 7757 24769 7791 24803
rect 7941 24769 7975 24803
rect 8309 24769 8343 24803
rect 10793 24769 10827 24803
rect 11253 24769 11287 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 11805 24769 11839 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 13921 24769 13955 24803
rect 14197 24769 14231 24803
rect 14381 24769 14415 24803
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 14933 24769 14967 24803
rect 15025 24769 15059 24803
rect 15301 24769 15335 24803
rect 15393 24769 15427 24803
rect 16773 24769 16807 24803
rect 17141 24769 17175 24803
rect 18889 24769 18923 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 19257 24769 19291 24803
rect 20085 24769 20119 24803
rect 20269 24769 20303 24803
rect 20913 24769 20947 24803
rect 21281 24769 21315 24803
rect 21373 24769 21407 24803
rect 22017 24769 22051 24803
rect 23213 24769 23247 24803
rect 25053 24769 25087 24803
rect 25421 24769 25455 24803
rect 26157 24769 26191 24803
rect 26341 24769 26375 24803
rect 27997 24769 28031 24803
rect 28273 24769 28307 24803
rect 28365 24769 28399 24803
rect 30113 24769 30147 24803
rect 31493 24769 31527 24803
rect 31585 24769 31619 24803
rect 32597 24769 32631 24803
rect 1501 24701 1535 24735
rect 4261 24701 4295 24735
rect 6653 24701 6687 24735
rect 7021 24701 7055 24735
rect 10057 24701 10091 24735
rect 30297 24701 30331 24735
rect 32689 24701 32723 24735
rect 6929 24633 6963 24667
rect 14013 24633 14047 24667
rect 22385 24633 22419 24667
rect 32137 24633 32171 24667
rect 2145 24565 2179 24599
rect 3709 24565 3743 24599
rect 5825 24565 5859 24599
rect 7757 24565 7791 24599
rect 10701 24565 10735 24599
rect 10977 24565 11011 24599
rect 11115 24565 11149 24599
rect 11529 24565 11563 24599
rect 15577 24565 15611 24599
rect 17325 24565 17359 24599
rect 19441 24565 19475 24599
rect 21373 24565 21407 24599
rect 21557 24565 21591 24599
rect 21833 24565 21867 24599
rect 24501 24565 24535 24599
rect 25237 24565 25271 24599
rect 25513 24565 25547 24599
rect 28457 24565 28491 24599
rect 28825 24565 28859 24599
rect 31309 24565 31343 24599
rect 31677 24565 31711 24599
rect 3065 24361 3099 24395
rect 5273 24361 5307 24395
rect 5733 24361 5767 24395
rect 9597 24361 9631 24395
rect 19073 24361 19107 24395
rect 23029 24361 23063 24395
rect 26617 24361 26651 24395
rect 27629 24361 27663 24395
rect 33609 24361 33643 24395
rect 12817 24293 12851 24327
rect 3801 24225 3835 24259
rect 13553 24225 13587 24259
rect 17601 24225 17635 24259
rect 19809 24225 19843 24259
rect 27077 24225 27111 24259
rect 27261 24225 27295 24259
rect 28574 24225 28608 24259
rect 29837 24225 29871 24259
rect 30757 24225 30791 24259
rect 31033 24225 31067 24259
rect 1685 24157 1719 24191
rect 3157 24157 3191 24191
rect 3341 24157 3375 24191
rect 3433 24157 3467 24191
rect 3617 24157 3651 24191
rect 5457 24157 5491 24191
rect 5549 24157 5583 24191
rect 6857 24157 6891 24191
rect 7113 24157 7147 24191
rect 7205 24157 7239 24191
rect 10977 24157 11011 24191
rect 11069 24157 11103 24191
rect 17325 24157 17359 24191
rect 21465 24157 21499 24191
rect 22937 24157 22971 24191
rect 24409 24157 24443 24191
rect 27537 24157 27571 24191
rect 28089 24157 28123 24191
rect 29009 24157 29043 24191
rect 29929 24157 29963 24191
rect 32597 24157 32631 24191
rect 32873 24157 32907 24191
rect 1952 24089 1986 24123
rect 3525 24089 3559 24123
rect 4046 24089 4080 24123
rect 7472 24089 7506 24123
rect 10732 24089 10766 24123
rect 11345 24089 11379 24123
rect 13369 24089 13403 24123
rect 22661 24089 22695 24123
rect 24685 24089 24719 24123
rect 26985 24089 27019 24123
rect 28457 24089 28491 24123
rect 3249 24021 3283 24055
rect 5181 24021 5215 24055
rect 8585 24021 8619 24055
rect 12909 24021 12943 24055
rect 13277 24021 13311 24055
rect 19257 24021 19291 24055
rect 21281 24021 21315 24055
rect 22569 24021 22603 24055
rect 26157 24021 26191 24055
rect 27997 24021 28031 24055
rect 28365 24021 28399 24055
rect 28733 24021 28767 24055
rect 28917 24021 28951 24055
rect 30297 24021 30331 24055
rect 32505 24021 32539 24055
rect 2053 23817 2087 23851
rect 3893 23817 3927 23851
rect 4445 23817 4479 23851
rect 7665 23817 7699 23851
rect 8861 23817 8895 23851
rect 11621 23817 11655 23851
rect 12357 23817 12391 23851
rect 13093 23817 13127 23851
rect 14197 23817 14231 23851
rect 16681 23817 16715 23851
rect 17141 23817 17175 23851
rect 18613 23817 18647 23851
rect 23489 23817 23523 23851
rect 24685 23817 24719 23851
rect 26065 23817 26099 23851
rect 28641 23817 28675 23851
rect 5181 23749 5215 23783
rect 21465 23749 21499 23783
rect 32321 23749 32355 23783
rect 2053 23681 2087 23715
rect 2237 23681 2271 23715
rect 2789 23681 2823 23715
rect 3341 23681 3375 23715
rect 3801 23681 3835 23715
rect 4261 23681 4295 23715
rect 4942 23681 4976 23715
rect 5089 23681 5123 23715
rect 5733 23681 5767 23715
rect 7849 23681 7883 23715
rect 8125 23681 8159 23715
rect 8493 23681 8527 23715
rect 9505 23681 9539 23715
rect 9597 23681 9631 23715
rect 9781 23681 9815 23715
rect 11805 23681 11839 23715
rect 12449 23681 12483 23715
rect 13737 23681 13771 23715
rect 14105 23681 14139 23715
rect 14565 23681 14599 23715
rect 15025 23681 15059 23715
rect 15577 23681 15611 23715
rect 16037 23681 16071 23715
rect 17049 23681 17083 23715
rect 17509 23681 17543 23715
rect 19165 23681 19199 23715
rect 19257 23681 19291 23715
rect 19625 23681 19659 23715
rect 22753 23681 22787 23715
rect 23581 23681 23615 23715
rect 23857 23681 23891 23715
rect 24869 23681 24903 23715
rect 24961 23681 24995 23715
rect 25237 23681 25271 23715
rect 26433 23681 26467 23715
rect 28273 23681 28307 23715
rect 28644 23681 28678 23715
rect 30481 23681 30515 23715
rect 30665 23681 30699 23715
rect 30757 23681 30791 23715
rect 30941 23681 30975 23715
rect 33609 23681 33643 23715
rect 33977 23681 34011 23715
rect 34161 23681 34195 23715
rect 4721 23613 4755 23647
rect 8677 23613 8711 23647
rect 9139 23613 9173 23647
rect 14657 23613 14691 23647
rect 14841 23613 14875 23647
rect 17325 23613 17359 23647
rect 18061 23613 18095 23647
rect 18705 23613 18739 23647
rect 18889 23613 18923 23647
rect 22477 23613 22511 23647
rect 26525 23613 26559 23647
rect 26709 23613 26743 23647
rect 28181 23613 28215 23647
rect 33885 23613 33919 23647
rect 4123 23545 4157 23579
rect 4813 23545 4847 23579
rect 9358 23545 9392 23579
rect 9597 23545 9631 23579
rect 32689 23545 32723 23579
rect 32781 23545 32815 23579
rect 3985 23477 4019 23511
rect 8033 23477 8067 23511
rect 8309 23477 8343 23511
rect 9229 23477 9263 23511
rect 13921 23477 13955 23511
rect 15853 23477 15887 23511
rect 18245 23477 18279 23511
rect 19809 23477 19843 23511
rect 21189 23477 21223 23511
rect 24593 23477 24627 23511
rect 25973 23477 26007 23511
rect 28825 23477 28859 23511
rect 30665 23477 30699 23511
rect 30849 23477 30883 23511
rect 32873 23477 32907 23511
rect 33977 23477 34011 23511
rect 17141 23273 17175 23307
rect 18245 23273 18279 23307
rect 21189 23273 21223 23307
rect 27905 23273 27939 23307
rect 28273 23273 28307 23307
rect 12173 23205 12207 23239
rect 33149 23205 33183 23239
rect 33333 23205 33367 23239
rect 2973 23137 3007 23171
rect 3893 23137 3927 23171
rect 12817 23137 12851 23171
rect 13645 23137 13679 23171
rect 15393 23137 15427 23171
rect 19441 23137 19475 23171
rect 19717 23137 19751 23171
rect 28181 23137 28215 23171
rect 28917 23137 28951 23171
rect 32873 23137 32907 23171
rect 2881 23069 2915 23103
rect 4537 23069 4571 23103
rect 6377 23069 6411 23103
rect 9045 23069 9079 23103
rect 9689 23069 9723 23103
rect 9781 23069 9815 23103
rect 9965 23069 9999 23103
rect 11897 23069 11931 23103
rect 14381 23069 14415 23103
rect 17417 23069 17451 23103
rect 18153 23069 18187 23103
rect 18429 23069 18463 23103
rect 18521 23069 18555 23103
rect 21465 23069 21499 23103
rect 21557 23069 21591 23103
rect 25053 23069 25087 23103
rect 25513 23069 25547 23103
rect 25789 23069 25823 23103
rect 27353 23069 27387 23103
rect 27629 23069 27663 23103
rect 28365 23069 28399 23103
rect 28457 23069 28491 23103
rect 28733 23069 28767 23103
rect 29009 23069 29043 23103
rect 30665 23069 30699 23103
rect 12541 23001 12575 23035
rect 13001 23001 13035 23035
rect 15669 23001 15703 23035
rect 17325 23001 17359 23035
rect 21373 23001 21407 23035
rect 21833 23001 21867 23035
rect 23581 23001 23615 23035
rect 28089 23001 28123 23035
rect 28549 23001 28583 23035
rect 3249 22933 3283 22967
rect 6929 22933 6963 22967
rect 9873 22933 9907 22967
rect 11713 22933 11747 22967
rect 12633 22933 12667 22967
rect 14473 22933 14507 22967
rect 17969 22933 18003 22967
rect 18613 22933 18647 22967
rect 25237 22933 25271 22967
rect 26525 22933 26559 22967
rect 27451 22933 27485 22967
rect 27537 22933 27571 22967
rect 27721 22933 27755 22967
rect 27889 22933 27923 22967
rect 29101 22933 29135 22967
rect 30757 22933 30791 22967
rect 2789 22729 2823 22763
rect 4721 22729 4755 22763
rect 6377 22729 6411 22763
rect 9137 22729 9171 22763
rect 13277 22729 13311 22763
rect 15209 22729 15243 22763
rect 19441 22729 19475 22763
rect 19809 22729 19843 22763
rect 20453 22729 20487 22763
rect 21557 22729 21591 22763
rect 22937 22729 22971 22763
rect 25513 22729 25547 22763
rect 27997 22729 28031 22763
rect 28273 22729 28307 22763
rect 29015 22729 29049 22763
rect 29101 22729 29135 22763
rect 29837 22729 29871 22763
rect 30573 22729 30607 22763
rect 32873 22729 32907 22763
rect 13737 22661 13771 22695
rect 17877 22661 17911 22695
rect 25605 22661 25639 22695
rect 30067 22661 30101 22695
rect 33241 22661 33275 22695
rect 33517 22661 33551 22695
rect 33011 22627 33045 22661
rect 3341 22593 3375 22627
rect 3608 22593 3642 22627
rect 4997 22593 5031 22627
rect 6377 22593 6411 22627
rect 6561 22593 6595 22627
rect 7481 22593 7515 22627
rect 7665 22593 7699 22627
rect 7757 22593 7791 22627
rect 8493 22593 8527 22627
rect 9505 22593 9539 22627
rect 11529 22593 11563 22627
rect 20361 22593 20395 22627
rect 20545 22593 20579 22627
rect 21097 22593 21131 22627
rect 21465 22593 21499 22627
rect 21833 22593 21867 22627
rect 22845 22593 22879 22627
rect 23489 22593 23523 22627
rect 24133 22593 24167 22627
rect 25329 22593 25363 22627
rect 25513 22593 25547 22627
rect 25881 22593 25915 22627
rect 26249 22593 26283 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 27721 22593 27755 22627
rect 27813 22593 27847 22627
rect 28457 22593 28491 22627
rect 28641 22593 28675 22627
rect 28917 22593 28951 22627
rect 29193 22593 29227 22627
rect 29469 22593 29503 22627
rect 30205 22593 30239 22627
rect 30297 22593 30331 22627
rect 30389 22593 30423 22627
rect 30665 22593 30699 22627
rect 30849 22593 30883 22627
rect 32781 22593 32815 22627
rect 33333 22593 33367 22627
rect 33609 22593 33643 22627
rect 3249 22525 3283 22559
rect 5089 22525 5123 22559
rect 5457 22525 5491 22559
rect 7297 22525 7331 22559
rect 8401 22525 8435 22559
rect 8861 22525 8895 22559
rect 10149 22525 10183 22559
rect 11805 22525 11839 22559
rect 13461 22525 13495 22559
rect 17601 22525 17635 22559
rect 19901 22525 19935 22559
rect 20085 22525 20119 22559
rect 20913 22525 20947 22559
rect 22109 22525 22143 22559
rect 23029 22525 23063 22559
rect 23581 22525 23615 22559
rect 25605 22525 25639 22559
rect 25973 22525 26007 22559
rect 27997 22525 28031 22559
rect 28549 22525 28583 22559
rect 28733 22525 28767 22559
rect 29377 22525 29411 22559
rect 29929 22525 29963 22559
rect 32505 22525 32539 22559
rect 5365 22457 5399 22491
rect 32689 22457 32723 22491
rect 33333 22457 33367 22491
rect 4997 22389 5031 22423
rect 6101 22389 6135 22423
rect 6745 22389 6779 22423
rect 7573 22389 7607 22423
rect 8658 22389 8692 22423
rect 8769 22389 8803 22423
rect 10057 22389 10091 22423
rect 10793 22389 10827 22423
rect 19349 22389 19383 22423
rect 22477 22389 22511 22423
rect 23765 22389 23799 22423
rect 24041 22389 24075 22423
rect 25789 22389 25823 22423
rect 27169 22389 27203 22423
rect 30757 22389 30791 22423
rect 32597 22389 32631 22423
rect 33057 22389 33091 22423
rect 5825 22185 5859 22219
rect 12449 22185 12483 22219
rect 13921 22185 13955 22219
rect 18061 22185 18095 22219
rect 20913 22185 20947 22219
rect 22109 22185 22143 22219
rect 26065 22185 26099 22219
rect 30021 22185 30055 22219
rect 30573 22185 30607 22219
rect 33701 22185 33735 22219
rect 17693 22117 17727 22151
rect 20545 22117 20579 22151
rect 3617 22049 3651 22083
rect 4353 22049 4387 22083
rect 12909 22049 12943 22083
rect 14105 22049 14139 22083
rect 18705 22049 18739 22083
rect 23673 22049 23707 22083
rect 28917 22049 28951 22083
rect 29009 22049 29043 22083
rect 32045 22049 32079 22083
rect 3985 21981 4019 22015
rect 6938 21981 6972 22015
rect 7205 21981 7239 22015
rect 7297 21981 7331 22015
rect 9505 21981 9539 22015
rect 10802 21981 10836 22015
rect 11069 21981 11103 22015
rect 12541 21981 12575 22015
rect 13185 21981 13219 22015
rect 14381 21981 14415 22015
rect 16405 21981 16439 22015
rect 16681 21981 16715 22015
rect 17509 21981 17543 22015
rect 18429 21981 18463 22015
rect 22293 21981 22327 22015
rect 23581 21981 23615 22015
rect 26249 21981 26283 22015
rect 26433 21981 26467 22015
rect 28733 21981 28767 22015
rect 29101 21981 29135 22015
rect 29285 21981 29319 22015
rect 29745 21981 29779 22015
rect 29929 21981 29963 22015
rect 30205 21981 30239 22015
rect 30481 21981 30515 22015
rect 30573 21981 30607 22015
rect 31769 21981 31803 22015
rect 31861 21981 31895 22015
rect 32505 21981 32539 22015
rect 32781 21981 32815 22015
rect 33149 21981 33183 22015
rect 33425 21981 33459 22015
rect 3372 21913 3406 21947
rect 3893 21913 3927 21947
rect 4620 21913 4654 21947
rect 7564 21913 7598 21947
rect 15209 21913 15243 21947
rect 15485 21913 15519 21947
rect 30684 21913 30718 21947
rect 30849 21913 30883 21947
rect 32321 21913 32355 21947
rect 33885 21913 33919 21947
rect 2237 21845 2271 21879
rect 5733 21845 5767 21879
rect 8677 21845 8711 21879
rect 8953 21845 8987 21879
rect 9689 21845 9723 21879
rect 15117 21845 15151 21879
rect 15393 21845 15427 21879
rect 15577 21845 15611 21879
rect 15761 21845 15795 21879
rect 17417 21845 17451 21879
rect 18521 21845 18555 21879
rect 20913 21845 20947 21879
rect 21097 21845 21131 21879
rect 23949 21845 23983 21879
rect 28549 21845 28583 21879
rect 29561 21845 29595 21879
rect 30389 21845 30423 21879
rect 32045 21845 32079 21879
rect 32689 21845 32723 21879
rect 32965 21845 32999 21879
rect 33333 21845 33367 21879
rect 33517 21845 33551 21879
rect 33680 21845 33714 21879
rect 4813 21641 4847 21675
rect 5549 21641 5583 21675
rect 7297 21641 7331 21675
rect 8033 21641 8067 21675
rect 8861 21641 8895 21675
rect 14565 21641 14599 21675
rect 15469 21641 15503 21675
rect 16681 21641 16715 21675
rect 23305 21641 23339 21675
rect 24691 21641 24725 21675
rect 31775 21641 31809 21675
rect 32137 21641 32171 21675
rect 6377 21573 6411 21607
rect 7113 21573 7147 21607
rect 10066 21573 10100 21607
rect 14749 21573 14783 21607
rect 15669 21573 15703 21607
rect 15945 21573 15979 21607
rect 21925 21573 21959 21607
rect 32965 21573 32999 21607
rect 3249 21505 3283 21539
rect 6101 21505 6135 21539
rect 6524 21505 6558 21539
rect 7205 21505 7239 21539
rect 7389 21505 7423 21539
rect 7849 21505 7883 21539
rect 8033 21505 8067 21539
rect 8125 21505 8159 21539
rect 8309 21505 8343 21539
rect 8493 21505 8527 21539
rect 8585 21505 8619 21539
rect 10333 21505 10367 21539
rect 11529 21505 11563 21539
rect 14381 21505 14415 21539
rect 14657 21505 14691 21539
rect 15117 21505 15151 21539
rect 17417 21505 17451 21539
rect 17693 21505 17727 21539
rect 17969 21505 18003 21539
rect 20085 21505 20119 21539
rect 20821 21505 20855 21539
rect 21097 21505 21131 21539
rect 23581 21505 23615 21539
rect 24133 21505 24167 21539
rect 24225 21505 24259 21539
rect 24593 21505 24627 21539
rect 24777 21505 24811 21539
rect 24869 21505 24903 21539
rect 25973 21505 26007 21539
rect 26249 21505 26283 21539
rect 31677 21505 31711 21539
rect 31861 21505 31895 21539
rect 31953 21505 31987 21539
rect 32321 21505 32355 21539
rect 32505 21505 32539 21539
rect 32873 21505 32907 21539
rect 33149 21505 33183 21539
rect 33333 21505 33367 21539
rect 5457 21437 5491 21471
rect 6745 21437 6779 21471
rect 8861 21437 8895 21471
rect 11805 21437 11839 21471
rect 20177 21437 20211 21471
rect 20269 21437 20303 21471
rect 21557 21437 21591 21471
rect 23305 21437 23339 21471
rect 24317 21437 24351 21471
rect 24409 21437 24443 21471
rect 26341 21437 26375 21471
rect 32413 21437 32447 21471
rect 32597 21437 32631 21471
rect 33241 21437 33275 21471
rect 6653 21369 6687 21403
rect 8953 21369 8987 21403
rect 14381 21369 14415 21403
rect 15301 21369 15335 21403
rect 15761 21369 15795 21403
rect 20821 21369 20855 21403
rect 3801 21301 3835 21335
rect 8677 21301 8711 21335
rect 13277 21301 13311 21335
rect 15485 21301 15519 21335
rect 17877 21301 17911 21335
rect 19717 21301 19751 21335
rect 22201 21301 22235 21335
rect 23489 21301 23523 21335
rect 23949 21301 23983 21335
rect 25881 21301 25915 21335
rect 26617 21301 26651 21335
rect 5181 21097 5215 21131
rect 5273 21097 5307 21131
rect 5549 21097 5583 21131
rect 9413 21097 9447 21131
rect 11805 21097 11839 21131
rect 12081 21097 12115 21131
rect 18613 21097 18647 21131
rect 25973 21097 26007 21131
rect 27905 21097 27939 21131
rect 30481 21097 30515 21131
rect 33149 21097 33183 21131
rect 14841 21029 14875 21063
rect 15025 21029 15059 21063
rect 15117 21029 15151 21063
rect 22569 21029 22603 21063
rect 28733 21029 28767 21063
rect 5365 20961 5399 20995
rect 9045 20961 9079 20995
rect 15209 20961 15243 20995
rect 20821 20961 20855 20995
rect 26065 20961 26099 20995
rect 27445 20961 27479 20995
rect 29193 20961 29227 20995
rect 5089 20893 5123 20927
rect 5457 20893 5491 20927
rect 5641 20893 5675 20927
rect 9137 20893 9171 20927
rect 11621 20893 11655 20927
rect 11989 20893 12023 20927
rect 14657 20893 14691 20927
rect 14841 20893 14875 20927
rect 14934 20893 14968 20927
rect 15577 20893 15611 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 19717 20893 19751 20927
rect 19993 20893 20027 20927
rect 22661 20893 22695 20927
rect 25973 20893 26007 20927
rect 27629 20893 27663 20927
rect 28089 20893 28123 20927
rect 28457 20893 28491 20927
rect 28549 20893 28583 20927
rect 28641 20893 28675 20927
rect 29009 20893 29043 20927
rect 30113 20893 30147 20927
rect 31309 20893 31343 20927
rect 31493 20893 31527 20927
rect 33057 20893 33091 20927
rect 15393 20825 15427 20859
rect 16957 20825 16991 20859
rect 18705 20825 18739 20859
rect 21097 20825 21131 20859
rect 22753 20825 22787 20859
rect 25605 20825 25639 20859
rect 25789 20825 25823 20859
rect 28181 20825 28215 20859
rect 28273 20825 28307 20859
rect 30297 20825 30331 20859
rect 31677 20825 31711 20859
rect 15761 20757 15795 20791
rect 16589 20757 16623 20791
rect 18429 20757 18463 20791
rect 19533 20757 19567 20791
rect 20085 20757 20119 20791
rect 25421 20757 25455 20791
rect 26341 20757 26375 20791
rect 27813 20757 27847 20791
rect 16957 20553 16991 20587
rect 20729 20553 20763 20587
rect 21373 20553 21407 20587
rect 21833 20553 21867 20587
rect 22201 20553 22235 20587
rect 24409 20553 24443 20587
rect 25881 20553 25915 20587
rect 28365 20553 28399 20587
rect 28641 20553 28675 20587
rect 31769 20553 31803 20587
rect 32597 20553 32631 20587
rect 13395 20485 13429 20519
rect 19257 20485 19291 20519
rect 24133 20485 24167 20519
rect 27813 20485 27847 20519
rect 27997 20485 28031 20519
rect 28181 20485 28215 20519
rect 30941 20485 30975 20519
rect 31171 20485 31205 20519
rect 9689 20417 9723 20451
rect 9781 20417 9815 20451
rect 11621 20417 11655 20451
rect 12541 20417 12575 20451
rect 13520 20417 13554 20451
rect 14749 20417 14783 20451
rect 17325 20417 17359 20451
rect 18061 20417 18095 20451
rect 18889 20417 18923 20451
rect 18981 20417 19015 20451
rect 21557 20417 21591 20451
rect 22845 20417 22879 20451
rect 23489 20417 23523 20451
rect 23673 20417 23707 20451
rect 23765 20417 23799 20451
rect 23903 20417 23937 20451
rect 24041 20417 24075 20451
rect 24224 20439 24258 20473
rect 24685 20417 24719 20451
rect 24869 20417 24903 20451
rect 24961 20417 24995 20451
rect 25145 20417 25179 20451
rect 25329 20417 25363 20451
rect 25421 20417 25455 20451
rect 25605 20417 25639 20451
rect 25789 20417 25823 20451
rect 26065 20417 26099 20451
rect 26341 20417 26375 20451
rect 27721 20417 27755 20451
rect 27905 20417 27939 20451
rect 28825 20417 28859 20451
rect 28917 20417 28951 20451
rect 29009 20417 29043 20451
rect 29193 20417 29227 20451
rect 29285 20417 29319 20451
rect 29929 20417 29963 20451
rect 30849 20417 30883 20451
rect 31033 20417 31067 20451
rect 31309 20417 31343 20451
rect 31401 20417 31435 20451
rect 31585 20417 31619 20451
rect 32965 20417 32999 20451
rect 12081 20349 12115 20383
rect 12633 20349 12667 20383
rect 12817 20349 12851 20383
rect 13001 20349 13035 20383
rect 14473 20349 14507 20383
rect 17417 20349 17451 20383
rect 17509 20349 17543 20383
rect 17785 20349 17819 20383
rect 22293 20349 22327 20383
rect 22477 20349 22511 20383
rect 23305 20349 23339 20383
rect 27445 20349 27479 20383
rect 33057 20349 33091 20383
rect 12173 20281 12207 20315
rect 13645 20281 13679 20315
rect 23121 20281 23155 20315
rect 23489 20281 23523 20315
rect 26157 20281 26191 20315
rect 26249 20281 26283 20315
rect 27077 20281 27111 20315
rect 9505 20213 9539 20247
rect 9873 20213 9907 20247
rect 11897 20213 11931 20247
rect 13093 20213 13127 20247
rect 14565 20213 14599 20247
rect 14657 20213 14691 20247
rect 24501 20213 24535 20247
rect 25053 20213 25087 20247
rect 26985 20213 27019 20247
rect 29745 20213 29779 20247
rect 30665 20213 30699 20247
rect 14565 20009 14599 20043
rect 17969 20009 18003 20043
rect 23305 20009 23339 20043
rect 29745 20009 29779 20043
rect 30113 20009 30147 20043
rect 31125 20009 31159 20043
rect 11989 19941 12023 19975
rect 15393 19941 15427 19975
rect 23121 19941 23155 19975
rect 9229 19873 9263 19907
rect 12541 19873 12575 19907
rect 13093 19873 13127 19907
rect 14381 19873 14415 19907
rect 14841 19873 14875 19907
rect 18981 19873 19015 19907
rect 22845 19873 22879 19907
rect 24777 19873 24811 19907
rect 30665 19873 30699 19907
rect 32413 19873 32447 19907
rect 32781 19873 32815 19907
rect 33977 19873 34011 19907
rect 8953 19805 8987 19839
rect 10793 19805 10827 19839
rect 11069 19805 11103 19839
rect 11897 19805 11931 19839
rect 14289 19805 14323 19839
rect 14749 19805 14783 19839
rect 14933 19805 14967 19839
rect 15577 19805 15611 19839
rect 15761 19805 15795 19839
rect 15879 19805 15913 19839
rect 16037 19805 16071 19839
rect 18705 19805 18739 19839
rect 24961 19805 24995 19839
rect 25145 19805 25179 19839
rect 25789 19805 25823 19839
rect 26341 19805 26375 19839
rect 26801 19805 26835 19839
rect 26893 19805 26927 19839
rect 27445 19805 27479 19839
rect 27629 19805 27663 19839
rect 27807 19805 27841 19839
rect 30481 19805 30515 19839
rect 31033 19805 31067 19839
rect 31217 19805 31251 19839
rect 31861 19805 31895 19839
rect 32045 19805 32079 19839
rect 32321 19805 32355 19839
rect 33057 19805 33091 19839
rect 33885 19805 33919 19839
rect 12357 19737 12391 19771
rect 13921 19737 13955 19771
rect 15669 19737 15703 19771
rect 25697 19737 25731 19771
rect 29561 19737 29595 19771
rect 10701 19669 10735 19703
rect 12449 19669 12483 19703
rect 27721 19669 27755 19703
rect 29761 19669 29795 19703
rect 29929 19669 29963 19703
rect 30573 19669 30607 19703
rect 31861 19669 31895 19703
rect 32689 19669 32723 19703
rect 33793 19669 33827 19703
rect 9873 19465 9907 19499
rect 14749 19465 14783 19499
rect 15117 19465 15151 19499
rect 15761 19465 15795 19499
rect 16313 19465 16347 19499
rect 24225 19465 24259 19499
rect 25697 19465 25731 19499
rect 31033 19465 31067 19499
rect 32505 19465 32539 19499
rect 32965 19465 32999 19499
rect 34345 19465 34379 19499
rect 16681 19397 16715 19431
rect 20821 19397 20855 19431
rect 24317 19397 24351 19431
rect 29561 19397 29595 19431
rect 32873 19397 32907 19431
rect 10609 19329 10643 19363
rect 10885 19329 10919 19363
rect 11897 19329 11931 19363
rect 13829 19329 13863 19363
rect 14933 19329 14967 19363
rect 15206 19329 15240 19363
rect 15945 19329 15979 19363
rect 16129 19329 16163 19363
rect 16221 19329 16255 19363
rect 16405 19329 16439 19363
rect 18521 19329 18555 19363
rect 19625 19329 19659 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 21833 19329 21867 19363
rect 22109 19329 22143 19363
rect 23581 19329 23615 19363
rect 23765 19329 23799 19363
rect 24133 19329 24167 19363
rect 25329 19329 25363 19363
rect 25513 19329 25547 19363
rect 27261 19329 27295 19363
rect 29285 19329 29319 19363
rect 32689 19329 32723 19363
rect 32965 19329 32999 19363
rect 33149 19329 33183 19363
rect 33609 19329 33643 19363
rect 14105 19261 14139 19295
rect 14197 19261 14231 19295
rect 23489 19261 23523 19295
rect 23673 19261 23707 19295
rect 24501 19261 24535 19295
rect 27353 19261 27387 19295
rect 33333 19261 33367 19295
rect 17969 19193 18003 19227
rect 13369 19125 13403 19159
rect 18613 19125 18647 19159
rect 20085 19125 20119 19159
rect 20913 19125 20947 19159
rect 22845 19125 22879 19159
rect 23305 19125 23339 19159
rect 23949 19125 23983 19159
rect 27537 19125 27571 19159
rect 13553 18921 13587 18955
rect 17969 18921 18003 18955
rect 18153 18921 18187 18955
rect 21465 18921 21499 18955
rect 22937 18921 22971 18955
rect 23765 18921 23799 18955
rect 24961 18921 24995 18955
rect 28733 18921 28767 18955
rect 30297 18921 30331 18955
rect 12633 18853 12667 18887
rect 23949 18853 23983 18887
rect 25053 18853 25087 18887
rect 10517 18785 10551 18819
rect 12173 18785 12207 18819
rect 12725 18785 12759 18819
rect 13093 18785 13127 18819
rect 13210 18785 13244 18819
rect 15209 18785 15243 18819
rect 15301 18785 15335 18819
rect 16957 18785 16991 18819
rect 18613 18785 18647 18819
rect 18705 18785 18739 18819
rect 21005 18785 21039 18819
rect 21925 18785 21959 18819
rect 23489 18785 23523 18819
rect 10793 18717 10827 18751
rect 11621 18717 11655 18751
rect 12265 18717 12299 18751
rect 13645 18717 13679 18751
rect 14381 18717 14415 18751
rect 14657 18717 14691 18751
rect 14933 18717 14967 18751
rect 15945 18717 15979 18751
rect 16313 18717 16347 18751
rect 16865 18717 16899 18751
rect 17325 18717 17359 18751
rect 17601 18717 17635 18751
rect 17785 18717 17819 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 18889 18717 18923 18751
rect 21649 18717 21683 18751
rect 22201 18717 22235 18751
rect 23397 18717 23431 18751
rect 23857 18717 23891 18751
rect 24041 18717 24075 18751
rect 26985 18717 27019 18751
rect 27261 18717 27295 18751
rect 27353 18717 27387 18751
rect 28641 18717 28675 18751
rect 30205 18717 30239 18751
rect 30757 18717 30791 18751
rect 13001 18649 13035 18683
rect 17463 18649 17497 18683
rect 17693 18649 17727 18683
rect 18981 18649 19015 18683
rect 20729 18649 20763 18683
rect 21189 18649 21223 18683
rect 25421 18649 25455 18683
rect 27169 18649 27203 18683
rect 13369 18581 13403 18615
rect 14657 18581 14691 18615
rect 17233 18581 17267 18615
rect 19257 18581 19291 18615
rect 21741 18581 21775 18615
rect 27537 18581 27571 18615
rect 30849 18581 30883 18615
rect 15209 18377 15243 18411
rect 16681 18377 16715 18411
rect 17877 18377 17911 18411
rect 19073 18377 19107 18411
rect 23857 18377 23891 18411
rect 25421 18377 25455 18411
rect 26157 18377 26191 18411
rect 27077 18377 27111 18411
rect 27445 18377 27479 18411
rect 29745 18377 29779 18411
rect 17325 18309 17359 18343
rect 18337 18309 18371 18343
rect 20085 18309 20119 18343
rect 20453 18309 20487 18343
rect 20913 18309 20947 18343
rect 24961 18309 24995 18343
rect 30113 18309 30147 18343
rect 15393 18241 15427 18275
rect 15945 18241 15979 18275
rect 18061 18241 18095 18275
rect 19165 18241 19199 18275
rect 20177 18241 20211 18275
rect 20361 18241 20395 18275
rect 20545 18241 20579 18275
rect 23305 18241 23339 18275
rect 25789 18241 25823 18275
rect 26801 18241 26835 18275
rect 29561 18241 29595 18275
rect 32505 18241 32539 18275
rect 33609 18241 33643 18275
rect 8493 18173 8527 18207
rect 8769 18173 8803 18207
rect 12541 18173 12575 18207
rect 13369 18173 13403 18207
rect 15669 18173 15703 18207
rect 15853 18173 15887 18207
rect 17141 18173 17175 18207
rect 17785 18173 17819 18207
rect 18153 18173 18187 18207
rect 19533 18173 19567 18207
rect 23581 18173 23615 18207
rect 25881 18173 25915 18207
rect 27537 18173 27571 18207
rect 27629 18173 27663 18207
rect 29837 18173 29871 18207
rect 32229 18173 32263 18207
rect 33333 18173 33367 18207
rect 15577 18105 15611 18139
rect 16773 18105 16807 18139
rect 17601 18105 17635 18139
rect 21097 18105 21131 18139
rect 25329 18105 25363 18139
rect 33241 18105 33275 18139
rect 10241 18037 10275 18071
rect 18337 18037 18371 18071
rect 20729 18037 20763 18071
rect 23673 18037 23707 18071
rect 26617 18037 26651 18071
rect 31585 18037 31619 18071
rect 34345 18037 34379 18071
rect 9045 17833 9079 17867
rect 9505 17833 9539 17867
rect 9873 17833 9907 17867
rect 20821 17833 20855 17867
rect 28089 17833 28123 17867
rect 30297 17833 30331 17867
rect 32781 17833 32815 17867
rect 33149 17833 33183 17867
rect 33517 17833 33551 17867
rect 20085 17765 20119 17799
rect 25605 17765 25639 17799
rect 10885 17697 10919 17731
rect 11529 17697 11563 17731
rect 14749 17697 14783 17731
rect 15025 17697 15059 17731
rect 22017 17697 22051 17731
rect 23765 17697 23799 17731
rect 24593 17697 24627 17731
rect 29653 17697 29687 17731
rect 30849 17697 30883 17731
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 10609 17629 10643 17663
rect 12357 17629 12391 17663
rect 12633 17629 12667 17663
rect 12817 17629 12851 17663
rect 14289 17629 14323 17663
rect 14473 17629 14507 17663
rect 14657 17629 14691 17663
rect 15117 17629 15151 17663
rect 18613 17629 18647 17663
rect 18889 17629 18923 17663
rect 20269 17629 20303 17663
rect 20361 17629 20395 17663
rect 22293 17629 22327 17663
rect 23305 17629 23339 17663
rect 24041 17629 24075 17663
rect 24869 17629 24903 17663
rect 26341 17629 26375 17663
rect 28365 17629 28399 17663
rect 28641 17629 28675 17663
rect 29745 17629 29779 17663
rect 32689 17629 32723 17663
rect 33241 17629 33275 17663
rect 14381 17561 14415 17595
rect 16681 17561 16715 17595
rect 20085 17561 20119 17595
rect 21097 17561 21131 17595
rect 21557 17561 21591 17595
rect 26617 17561 26651 17595
rect 28273 17561 28307 17595
rect 12725 17493 12759 17527
rect 14105 17493 14139 17527
rect 16405 17493 16439 17527
rect 21833 17493 21867 17527
rect 23029 17493 23063 17527
rect 23213 17493 23247 17527
rect 28733 17493 28767 17527
rect 30113 17493 30147 17527
rect 30665 17493 30699 17527
rect 30757 17493 30791 17527
rect 33701 17493 33735 17527
rect 13829 17289 13863 17323
rect 14657 17289 14691 17323
rect 19625 17289 19659 17323
rect 21649 17289 21683 17323
rect 23581 17289 23615 17323
rect 30849 17289 30883 17323
rect 32889 17289 32923 17323
rect 38301 17289 38335 17323
rect 10425 17221 10459 17255
rect 22109 17221 22143 17255
rect 32413 17221 32447 17255
rect 32597 17221 32631 17255
rect 32689 17221 32723 17255
rect 33149 17221 33183 17255
rect 11529 17153 11563 17187
rect 14197 17153 14231 17187
rect 14289 17153 14323 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 17325 17153 17359 17187
rect 17785 17153 17819 17187
rect 18613 17153 18647 17187
rect 18889 17153 18923 17187
rect 21465 17153 21499 17187
rect 24317 17153 24351 17187
rect 24409 17153 24443 17187
rect 25699 17153 25733 17187
rect 25973 17153 26007 17187
rect 29837 17153 29871 17187
rect 31125 17153 31159 17187
rect 32321 17153 32355 17187
rect 33425 17153 33459 17187
rect 38485 17153 38519 17187
rect 17417 17085 17451 17119
rect 21833 17085 21867 17119
rect 24041 17085 24075 17119
rect 24685 17085 24719 17119
rect 27629 17085 27663 17119
rect 27905 17085 27939 17119
rect 29377 17085 29411 17119
rect 29929 17085 29963 17119
rect 30113 17085 30147 17119
rect 30849 17085 30883 17119
rect 33149 17085 33183 17119
rect 16957 17017 16991 17051
rect 24961 17017 24995 17051
rect 29469 17017 29503 17051
rect 32597 17017 32631 17051
rect 33333 17017 33367 17051
rect 8953 16949 8987 16983
rect 11621 16949 11655 16983
rect 14473 16949 14507 16983
rect 17693 16949 17727 16983
rect 31033 16949 31067 16983
rect 32873 16949 32907 16983
rect 33057 16949 33091 16983
rect 9597 16745 9631 16779
rect 11897 16745 11931 16779
rect 12449 16745 12483 16779
rect 13553 16745 13587 16779
rect 21649 16745 21683 16779
rect 28181 16745 28215 16779
rect 29653 16745 29687 16779
rect 30757 16745 30791 16779
rect 31677 16745 31711 16779
rect 33701 16745 33735 16779
rect 13645 16677 13679 16711
rect 18797 16677 18831 16711
rect 33241 16677 33275 16711
rect 9229 16609 9263 16643
rect 10057 16609 10091 16643
rect 10241 16609 10275 16643
rect 10977 16609 11011 16643
rect 11345 16609 11379 16643
rect 11805 16609 11839 16643
rect 12633 16609 12667 16643
rect 13369 16609 13403 16643
rect 14381 16609 14415 16643
rect 15761 16609 15795 16643
rect 17785 16609 17819 16643
rect 20177 16609 20211 16643
rect 22109 16609 22143 16643
rect 22201 16609 22235 16643
rect 23673 16609 23707 16643
rect 31034 16609 31068 16643
rect 31217 16575 31251 16609
rect 10885 16541 10919 16575
rect 11437 16541 11471 16575
rect 11897 16541 11931 16575
rect 11989 16541 12023 16575
rect 12357 16541 12391 16575
rect 13277 16541 13311 16575
rect 13645 16541 13679 16575
rect 13921 16541 13955 16575
rect 14289 16541 14323 16575
rect 18061 16541 18095 16575
rect 19441 16541 19475 16575
rect 19625 16541 19659 16575
rect 20085 16541 20119 16575
rect 22569 16541 22603 16575
rect 23397 16541 23431 16575
rect 24685 16541 24719 16575
rect 28365 16541 28399 16575
rect 29837 16541 29871 16575
rect 29929 16541 29963 16575
rect 30139 16541 30173 16575
rect 30297 16541 30331 16575
rect 30941 16541 30975 16575
rect 31125 16541 31159 16575
rect 31401 16541 31435 16575
rect 32597 16541 32631 16575
rect 32781 16541 32815 16575
rect 32873 16541 32907 16575
rect 9413 16473 9447 16507
rect 12633 16473 12667 16507
rect 13737 16473 13771 16507
rect 16037 16473 16071 16507
rect 20361 16473 20395 16507
rect 20545 16473 20579 16507
rect 26065 16473 26099 16507
rect 30021 16473 30055 16507
rect 31677 16473 31711 16507
rect 32965 16473 32999 16507
rect 33885 16473 33919 16507
rect 9965 16405 9999 16439
rect 10425 16405 10459 16439
rect 10793 16405 10827 16439
rect 12265 16405 12299 16439
rect 12909 16405 12943 16439
rect 14657 16405 14691 16439
rect 17509 16405 17543 16439
rect 19625 16405 19659 16439
rect 19717 16405 19751 16439
rect 20729 16405 20763 16439
rect 22017 16405 22051 16439
rect 24501 16405 24535 16439
rect 26157 16405 26191 16439
rect 31493 16405 31527 16439
rect 32413 16405 32447 16439
rect 33425 16405 33459 16439
rect 33517 16405 33551 16439
rect 33685 16405 33719 16439
rect 13553 16201 13587 16235
rect 14381 16201 14415 16235
rect 16313 16201 16347 16235
rect 18981 16201 19015 16235
rect 32137 16201 32171 16235
rect 33793 16201 33827 16235
rect 9689 16133 9723 16167
rect 11069 16133 11103 16167
rect 12449 16133 12483 16167
rect 17325 16133 17359 16167
rect 18521 16133 18555 16167
rect 20913 16133 20947 16167
rect 23673 16133 23707 16167
rect 30757 16133 30791 16167
rect 31033 16133 31067 16167
rect 9781 16065 9815 16099
rect 10149 16065 10183 16099
rect 11253 16065 11287 16099
rect 11345 16065 11379 16099
rect 11621 16065 11655 16099
rect 11805 16065 11839 16099
rect 12265 16065 12299 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 14565 16065 14599 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 14933 16065 14967 16099
rect 16497 16065 16531 16099
rect 17233 16065 17267 16099
rect 19993 16065 20027 16099
rect 20177 16065 20211 16099
rect 24133 16065 24167 16099
rect 27261 16065 27295 16099
rect 28917 16065 28951 16099
rect 30573 16065 30607 16099
rect 30941 16065 30975 16099
rect 31217 16065 31251 16099
rect 31585 16065 31619 16099
rect 31769 16065 31803 16099
rect 32575 16065 32609 16099
rect 32965 16095 32999 16129
rect 34529 16065 34563 16099
rect 7757 15997 7791 16031
rect 8033 15997 8067 16031
rect 9873 15997 9907 16031
rect 12633 15997 12667 16031
rect 17417 15997 17451 16031
rect 23857 15997 23891 16031
rect 25053 15997 25087 16031
rect 25329 15997 25363 16031
rect 26801 15997 26835 16031
rect 26985 15997 27019 16031
rect 29009 15997 29043 16031
rect 31401 15997 31435 16031
rect 31493 15997 31527 16031
rect 32689 15997 32723 16031
rect 34805 15997 34839 16031
rect 10885 15929 10919 15963
rect 11069 15929 11103 15963
rect 16865 15929 16899 15963
rect 18797 15929 18831 15963
rect 21189 15929 21223 15963
rect 27997 15929 28031 15963
rect 33701 15929 33735 15963
rect 9505 15861 9539 15895
rect 11989 15861 12023 15895
rect 20085 15861 20119 15895
rect 21373 15861 21407 15895
rect 23581 15861 23615 15895
rect 24869 15861 24903 15895
rect 29193 15861 29227 15895
rect 32505 15861 32539 15895
rect 8401 15657 8435 15691
rect 13737 15657 13771 15691
rect 14749 15657 14783 15691
rect 27169 15657 27203 15691
rect 11069 15589 11103 15623
rect 20269 15589 20303 15623
rect 23305 15589 23339 15623
rect 28549 15589 28583 15623
rect 30481 15589 30515 15623
rect 31033 15589 31067 15623
rect 10701 15521 10735 15555
rect 14565 15521 14599 15555
rect 16865 15521 16899 15555
rect 20453 15521 20487 15555
rect 23765 15521 23799 15555
rect 8585 15453 8619 15487
rect 9873 15453 9907 15487
rect 10149 15453 10183 15487
rect 11897 15453 11931 15487
rect 12081 15453 12115 15487
rect 13461 15453 13495 15487
rect 13599 15453 13633 15487
rect 13921 15453 13955 15487
rect 14473 15453 14507 15487
rect 14749 15453 14783 15487
rect 16773 15453 16807 15487
rect 20177 15453 20211 15487
rect 20729 15453 20763 15487
rect 20913 15453 20947 15487
rect 21005 15453 21039 15487
rect 23673 15453 23707 15487
rect 27905 15453 27939 15487
rect 28181 15453 28215 15487
rect 29745 15453 29779 15487
rect 30021 15453 30055 15487
rect 30205 15453 30239 15487
rect 30665 15453 30699 15487
rect 30941 15453 30975 15487
rect 31033 15453 31067 15487
rect 25237 15385 25271 15419
rect 26985 15385 27019 15419
rect 28273 15385 28307 15419
rect 29561 15385 29595 15419
rect 31125 15385 31159 15419
rect 31309 15385 31343 15419
rect 9137 15317 9171 15351
rect 11161 15317 11195 15351
rect 12265 15317 12299 15351
rect 13921 15317 13955 15351
rect 14933 15317 14967 15351
rect 17141 15317 17175 15351
rect 20453 15317 20487 15351
rect 20545 15317 20579 15351
rect 28733 15317 28767 15351
rect 29929 15317 29963 15351
rect 30113 15317 30147 15351
rect 30849 15317 30883 15351
rect 14749 15113 14783 15147
rect 18521 15113 18555 15147
rect 22201 15113 22235 15147
rect 25881 15113 25915 15147
rect 26433 15113 26467 15147
rect 26985 15113 27019 15147
rect 27445 15113 27479 15147
rect 11713 15045 11747 15079
rect 17325 15045 17359 15079
rect 21189 15045 21223 15079
rect 21373 15045 21407 15079
rect 23673 15045 23707 15079
rect 25697 15045 25731 15079
rect 27997 15045 28031 15079
rect 11529 14977 11563 15011
rect 14105 14977 14139 15011
rect 14381 14977 14415 15011
rect 14565 14977 14599 15011
rect 17049 14977 17083 15011
rect 18245 14977 18279 15011
rect 19993 14977 20027 15011
rect 20085 14977 20119 15011
rect 20177 14977 20211 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 20729 14977 20763 15011
rect 21557 14977 21591 15011
rect 25513 14977 25547 15011
rect 25789 14977 25823 15011
rect 26065 14977 26099 15011
rect 26525 14977 26559 15011
rect 27353 14977 27387 15011
rect 28825 14977 28859 15011
rect 29009 14977 29043 15011
rect 29929 14977 29963 15011
rect 30113 14977 30147 15011
rect 14013 14909 14047 14943
rect 16681 14909 16715 14943
rect 17141 14909 17175 14943
rect 17693 14909 17727 14943
rect 17785 14909 17819 14943
rect 17877 14909 17911 14943
rect 17969 14909 18003 14943
rect 18521 14909 18555 14943
rect 20821 14909 20855 14943
rect 25237 14909 25271 14943
rect 27537 14909 27571 14943
rect 28457 14909 28491 14943
rect 30021 14909 30055 14943
rect 13737 14841 13771 14875
rect 28273 14841 28307 14875
rect 11897 14773 11931 14807
rect 18153 14773 18187 14807
rect 18337 14773 18371 14807
rect 19809 14773 19843 14807
rect 21097 14773 21131 14807
rect 23765 14773 23799 14807
rect 28825 14773 28859 14807
rect 14197 14569 14231 14603
rect 16773 14569 16807 14603
rect 17601 14569 17635 14603
rect 18061 14569 18095 14603
rect 20085 14569 20119 14603
rect 22477 14569 22511 14603
rect 27261 14569 27295 14603
rect 29009 14569 29043 14603
rect 31125 14569 31159 14603
rect 31585 14569 31619 14603
rect 19625 14501 19659 14535
rect 21833 14501 21867 14535
rect 27445 14501 27479 14535
rect 32689 14501 32723 14535
rect 9597 14433 9631 14467
rect 11529 14433 11563 14467
rect 12265 14433 12299 14467
rect 16957 14433 16991 14467
rect 19901 14433 19935 14467
rect 22109 14433 22143 14467
rect 23857 14433 23891 14467
rect 30941 14433 30975 14467
rect 32229 14433 32263 14467
rect 32505 14433 32539 14467
rect 8585 14365 8619 14399
rect 11437 14365 11471 14399
rect 12817 14365 12851 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 14105 14365 14139 14399
rect 15117 14365 15151 14399
rect 15209 14365 15243 14399
rect 15393 14365 15427 14399
rect 15853 14365 15887 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 16221 14365 16255 14399
rect 17049 14365 17083 14399
rect 17417 14365 17451 14399
rect 17785 14365 17819 14399
rect 17877 14365 17911 14399
rect 18245 14365 18279 14399
rect 18521 14365 18555 14399
rect 18613 14365 18647 14399
rect 19073 14365 19107 14399
rect 19257 14365 19291 14399
rect 19441 14365 19475 14399
rect 20177 14365 20211 14399
rect 22201 14365 22235 14399
rect 22661 14365 22695 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 24409 14365 24443 14399
rect 25237 14365 25271 14399
rect 25513 14365 25547 14399
rect 26801 14365 26835 14399
rect 26893 14365 26927 14399
rect 27077 14365 27111 14399
rect 27629 14365 27663 14399
rect 27721 14365 27755 14399
rect 27905 14365 27939 14399
rect 27997 14365 28031 14399
rect 30205 14365 30239 14399
rect 31401 14365 31435 14399
rect 31493 14365 31527 14399
rect 31677 14365 31711 14399
rect 32137 14365 32171 14399
rect 32597 14365 32631 14399
rect 32873 14365 32907 14399
rect 12909 14297 12943 14331
rect 15577 14297 15611 14331
rect 17325 14297 17359 14331
rect 17601 14297 17635 14331
rect 18981 14297 19015 14331
rect 19349 14297 19383 14331
rect 22753 14297 22787 14331
rect 28641 14297 28675 14331
rect 28825 14297 28859 14331
rect 8401 14229 8435 14263
rect 8953 14229 8987 14263
rect 9321 14229 9355 14263
rect 9413 14229 9447 14263
rect 12633 14229 12667 14263
rect 14565 14229 14599 14263
rect 15669 14229 15703 14263
rect 18429 14229 18463 14263
rect 18889 14229 18923 14263
rect 23305 14229 23339 14263
rect 23673 14229 23707 14263
rect 23765 14229 23799 14263
rect 30297 14229 30331 14263
rect 33057 14229 33091 14263
rect 9505 14025 9539 14059
rect 11345 14025 11379 14059
rect 12357 14025 12391 14059
rect 17785 14025 17819 14059
rect 18705 14025 18739 14059
rect 20821 14025 20855 14059
rect 23581 14025 23615 14059
rect 27077 14025 27111 14059
rect 31493 14025 31527 14059
rect 31861 14025 31895 14059
rect 8033 13957 8067 13991
rect 30021 13957 30055 13991
rect 30113 13957 30147 13991
rect 7757 13889 7791 13923
rect 9689 13889 9723 13923
rect 9965 13889 9999 13923
rect 10977 13889 11011 13923
rect 11989 13889 12023 13923
rect 13829 13889 13863 13923
rect 14013 13889 14047 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 14289 13889 14323 13923
rect 14933 13889 14967 13923
rect 15025 13889 15059 13923
rect 15209 13889 15243 13923
rect 15393 13889 15427 13923
rect 17601 13889 17635 13923
rect 17785 13889 17819 13923
rect 18613 13889 18647 13923
rect 18797 13889 18831 13923
rect 19625 13889 19659 13923
rect 21097 13889 21131 13923
rect 22201 13889 22235 13923
rect 22845 13889 22879 13923
rect 22937 13889 22971 13923
rect 23121 13889 23155 13923
rect 23397 13889 23431 13923
rect 24869 13889 24903 13923
rect 25421 13889 25455 13923
rect 25605 13889 25639 13923
rect 27261 13889 27295 13923
rect 27629 13889 27663 13923
rect 27813 13889 27847 13923
rect 29883 13889 29917 13923
rect 30205 13889 30239 13923
rect 31217 13889 31251 13923
rect 31401 13889 31435 13923
rect 31677 13889 31711 13923
rect 31953 13889 31987 13923
rect 32505 13889 32539 13923
rect 11069 13821 11103 13855
rect 12081 13821 12115 13855
rect 14749 13821 14783 13855
rect 14841 13821 14875 13855
rect 19349 13821 19383 13855
rect 19441 13821 19475 13855
rect 20821 13821 20855 13855
rect 22109 13821 22143 13855
rect 23305 13821 23339 13855
rect 27537 13821 27571 13855
rect 29745 13821 29779 13855
rect 31309 13821 31343 13855
rect 32413 13821 32447 13855
rect 10701 13753 10735 13787
rect 14473 13753 14507 13787
rect 19809 13753 19843 13787
rect 22569 13753 22603 13787
rect 32137 13753 32171 13787
rect 14565 13685 14599 13719
rect 15301 13685 15335 13719
rect 21005 13685 21039 13719
rect 24961 13685 24995 13719
rect 25513 13685 25547 13719
rect 27445 13685 27479 13719
rect 27997 13685 28031 13719
rect 30389 13685 30423 13719
rect 8677 13481 8711 13515
rect 13921 13481 13955 13515
rect 14197 13481 14231 13515
rect 18245 13481 18279 13515
rect 23305 13481 23339 13515
rect 27537 13481 27571 13515
rect 28089 13481 28123 13515
rect 28181 13481 28215 13515
rect 31493 13481 31527 13515
rect 31861 13481 31895 13515
rect 9045 13413 9079 13447
rect 11253 13413 11287 13447
rect 13369 13413 13403 13447
rect 15117 13413 15151 13447
rect 22017 13413 22051 13447
rect 11345 13345 11379 13379
rect 14565 13345 14599 13379
rect 18061 13345 18095 13379
rect 21557 13345 21591 13379
rect 24685 13345 24719 13379
rect 28273 13345 28307 13379
rect 32229 13345 32263 13379
rect 8769 13277 8803 13311
rect 9781 13277 9815 13311
rect 10057 13277 10091 13311
rect 13093 13277 13127 13311
rect 13464 13255 13498 13289
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 14473 13277 14507 13311
rect 14933 13277 14967 13311
rect 17969 13277 18003 13311
rect 21649 13277 21683 13311
rect 22845 13277 22879 13311
rect 22937 13277 22971 13311
rect 23121 13277 23155 13311
rect 24777 13277 24811 13311
rect 25237 13277 25271 13311
rect 25329 13277 25363 13311
rect 25513 13277 25547 13311
rect 27537 13277 27571 13311
rect 27813 13277 27847 13311
rect 27997 13277 28031 13311
rect 29561 13277 29595 13311
rect 31401 13277 31435 13311
rect 31585 13277 31619 13311
rect 32045 13277 32079 13311
rect 10885 13209 10919 13243
rect 12265 13209 12299 13243
rect 12449 13209 12483 13243
rect 13185 13209 13219 13243
rect 13369 13209 13403 13243
rect 14749 13209 14783 13243
rect 29837 13209 29871 13243
rect 25145 13141 25179 13175
rect 25697 13141 25731 13175
rect 27721 13141 27755 13175
rect 31309 13141 31343 13175
rect 12633 12937 12667 12971
rect 12909 12937 12943 12971
rect 13093 12937 13127 12971
rect 17325 12937 17359 12971
rect 21195 12937 21229 12971
rect 22746 12937 22780 12971
rect 24777 12937 24811 12971
rect 27629 12937 27663 12971
rect 27721 12937 27755 12971
rect 28365 12937 28399 12971
rect 29285 12937 29319 12971
rect 29561 12937 29595 12971
rect 30021 12937 30055 12971
rect 9781 12869 9815 12903
rect 21097 12869 21131 12903
rect 22661 12869 22695 12903
rect 22845 12869 22879 12903
rect 25697 12869 25731 12903
rect 27353 12869 27387 12903
rect 30113 12869 30147 12903
rect 30665 12869 30699 12903
rect 12541 12801 12575 12835
rect 12725 12801 12759 12835
rect 13277 12801 13311 12835
rect 13369 12801 13403 12835
rect 15669 12801 15703 12835
rect 16865 12801 16899 12835
rect 17785 12801 17819 12835
rect 18797 12801 18831 12835
rect 20637 12801 20671 12835
rect 20821 12801 20855 12835
rect 21281 12801 21315 12835
rect 21373 12801 21407 12835
rect 22569 12801 22603 12835
rect 24777 12801 24811 12835
rect 24961 12801 24995 12835
rect 25329 12801 25363 12835
rect 26249 12801 26283 12835
rect 27537 12801 27571 12835
rect 27997 12801 28031 12835
rect 28181 12801 28215 12835
rect 28917 12801 28951 12835
rect 29377 12801 29411 12835
rect 30849 12801 30883 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 9873 12733 9907 12767
rect 10057 12733 10091 12767
rect 11805 12733 11839 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 13645 12733 13679 12767
rect 13737 12733 13771 12767
rect 16957 12733 16991 12767
rect 18889 12733 18923 12767
rect 25237 12733 25271 12767
rect 26157 12733 26191 12767
rect 28825 12733 28859 12767
rect 30205 12733 30239 12767
rect 30481 12733 30515 12767
rect 12357 12665 12391 12699
rect 17233 12665 17267 12699
rect 17417 12665 17451 12699
rect 19165 12665 19199 12699
rect 25881 12665 25915 12699
rect 27905 12665 27939 12699
rect 29653 12665 29687 12699
rect 9413 12597 9447 12631
rect 12265 12597 12299 12631
rect 15485 12597 15519 12631
rect 21005 12597 21039 12631
rect 25053 12597 25087 12631
rect 32505 12597 32539 12631
rect 12633 12393 12667 12427
rect 13001 12393 13035 12427
rect 16773 12393 16807 12427
rect 19073 12393 19107 12427
rect 31309 12393 31343 12427
rect 31953 12393 31987 12427
rect 12357 12325 12391 12359
rect 20361 12325 20395 12359
rect 23213 12325 23247 12359
rect 31769 12325 31803 12359
rect 33057 12325 33091 12359
rect 11897 12257 11931 12291
rect 15301 12257 15335 12291
rect 16957 12257 16991 12291
rect 18061 12257 18095 12291
rect 20177 12257 20211 12291
rect 22937 12257 22971 12291
rect 25053 12257 25087 12291
rect 25329 12257 25363 12291
rect 31493 12257 31527 12291
rect 8585 12189 8619 12223
rect 8953 12189 8987 12223
rect 11989 12189 12023 12223
rect 12541 12189 12575 12223
rect 15025 12189 15059 12223
rect 17233 12189 17267 12223
rect 18337 12189 18371 12223
rect 20085 12189 20119 12223
rect 20545 12189 20579 12223
rect 20729 12189 20763 12223
rect 20913 12189 20947 12223
rect 21281 12189 21315 12223
rect 21833 12189 21867 12223
rect 22017 12189 22051 12223
rect 22845 12189 22879 12223
rect 23489 12189 23523 12223
rect 23857 12189 23891 12223
rect 24961 12189 24995 12223
rect 25973 12189 26007 12223
rect 26157 12189 26191 12223
rect 27629 12189 27663 12223
rect 31217 12189 31251 12223
rect 31401 12189 31435 12223
rect 32045 12189 32079 12223
rect 32321 12189 32355 12223
rect 33885 12189 33919 12223
rect 34161 12189 34195 12223
rect 9229 12121 9263 12155
rect 20637 12121 20671 12155
rect 21005 12121 21039 12155
rect 21373 12121 21407 12155
rect 21649 12121 21683 12155
rect 23581 12121 23615 12155
rect 23673 12121 23707 12155
rect 26065 12121 26099 12155
rect 27813 12121 27847 12155
rect 8769 12053 8803 12087
rect 10701 12053 10735 12087
rect 17969 12053 18003 12087
rect 19717 12053 19751 12087
rect 21189 12053 21223 12087
rect 21557 12053 21591 12087
rect 23305 12053 23339 12087
rect 27445 12053 27479 12087
rect 33149 12053 33183 12087
rect 9045 11849 9079 11883
rect 11345 11849 11379 11883
rect 16313 11849 16347 11883
rect 16681 11849 16715 11883
rect 17049 11849 17083 11883
rect 19441 11849 19475 11883
rect 20361 11849 20395 11883
rect 21021 11849 21055 11883
rect 21189 11849 21223 11883
rect 25513 11849 25547 11883
rect 26249 11849 26283 11883
rect 27261 11849 27295 11883
rect 32597 11849 32631 11883
rect 17141 11781 17175 11815
rect 19717 11781 19751 11815
rect 19809 11781 19843 11815
rect 20821 11781 20855 11815
rect 25605 11781 25639 11815
rect 25789 11781 25823 11815
rect 27629 11781 27663 11815
rect 27829 11781 27863 11815
rect 32137 11781 32171 11815
rect 8953 11713 8987 11747
rect 9965 11713 9999 11747
rect 10609 11713 10643 11747
rect 16405 11713 16439 11747
rect 19625 11713 19659 11747
rect 19993 11713 20027 11747
rect 20545 11713 20579 11747
rect 20729 11713 20763 11747
rect 25237 11713 25271 11747
rect 25421 11713 25455 11747
rect 26065 11713 26099 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 28825 11713 28859 11747
rect 29009 11713 29043 11747
rect 31493 11713 31527 11747
rect 10241 11645 10275 11679
rect 10333 11645 10367 11679
rect 17325 11645 17359 11679
rect 25881 11645 25915 11679
rect 31401 11645 31435 11679
rect 9229 11577 9263 11611
rect 26985 11577 27019 11611
rect 27537 11577 27571 11611
rect 31861 11577 31895 11611
rect 32413 11577 32447 11611
rect 21005 11509 21039 11543
rect 27813 11509 27847 11543
rect 27997 11509 28031 11543
rect 28917 11509 28951 11543
rect 15945 11305 15979 11339
rect 16129 11305 16163 11339
rect 24409 11305 24443 11339
rect 25881 11305 25915 11339
rect 28733 11305 28767 11339
rect 12081 11237 12115 11271
rect 23673 11237 23707 11271
rect 13645 11169 13679 11203
rect 14105 11169 14139 11203
rect 14289 11169 14323 11203
rect 14381 11169 14415 11203
rect 22937 11169 22971 11203
rect 23857 11169 23891 11203
rect 24777 11169 24811 11203
rect 25145 11169 25179 11203
rect 25237 11169 25271 11203
rect 25421 11169 25455 11203
rect 27813 11169 27847 11203
rect 28273 11169 28307 11203
rect 11345 11101 11379 11135
rect 11621 11101 11655 11135
rect 11713 11101 11747 11135
rect 11897 11101 11931 11135
rect 12173 11101 12207 11135
rect 12449 11101 12483 11135
rect 13553 11101 13587 11135
rect 15025 11101 15059 11135
rect 15117 11101 15151 11135
rect 15209 11101 15243 11135
rect 15485 11101 15519 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 17693 11101 17727 11135
rect 17785 11101 17819 11135
rect 17969 11101 18003 11135
rect 18061 11101 18095 11135
rect 22661 11101 22695 11135
rect 24409 11101 24443 11135
rect 24593 11101 24627 11135
rect 25697 11101 25731 11135
rect 27905 11101 27939 11135
rect 27997 11101 28031 11135
rect 28181 11101 28215 11135
rect 28365 11101 28399 11135
rect 28549 11101 28583 11135
rect 29101 11101 29135 11135
rect 29377 11101 29411 11135
rect 30481 11101 30515 11135
rect 11437 11033 11471 11067
rect 12265 11033 12299 11067
rect 12633 11033 12667 11067
rect 23397 11033 23431 11067
rect 25513 11033 25547 11067
rect 13921 10965 13955 10999
rect 14749 10965 14783 10999
rect 15393 10965 15427 10999
rect 18245 10965 18279 10999
rect 22293 10965 22327 10999
rect 22753 10965 22787 10999
rect 28917 10965 28951 10999
rect 29285 10965 29319 10999
rect 30389 10965 30423 10999
rect 11713 10761 11747 10795
rect 14381 10761 14415 10795
rect 16053 10761 16087 10795
rect 16221 10761 16255 10795
rect 18245 10761 18279 10795
rect 24041 10761 24075 10795
rect 24777 10761 24811 10795
rect 28365 10761 28399 10795
rect 29929 10761 29963 10795
rect 31309 10761 31343 10795
rect 32137 10761 32171 10795
rect 15853 10693 15887 10727
rect 27077 10693 27111 10727
rect 28615 10693 28649 10727
rect 28825 10693 28859 10727
rect 29193 10693 29227 10727
rect 30633 10693 30667 10727
rect 30849 10693 30883 10727
rect 30941 10693 30975 10727
rect 10057 10625 10091 10659
rect 10149 10625 10183 10659
rect 10701 10625 10735 10659
rect 11621 10625 11655 10659
rect 11805 10625 11839 10659
rect 12265 10625 12299 10659
rect 14105 10625 14139 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 14657 10625 14691 10659
rect 15485 10625 15519 10659
rect 15577 10625 15611 10659
rect 15761 10625 15795 10659
rect 16313 10625 16347 10659
rect 16497 10625 16531 10659
rect 16957 10625 16991 10659
rect 17233 10625 17267 10659
rect 17417 10625 17451 10659
rect 17509 10625 17543 10659
rect 17693 10625 17727 10659
rect 17969 10625 18003 10659
rect 18429 10625 18463 10659
rect 18613 10625 18647 10659
rect 18981 10625 19015 10659
rect 22017 10625 22051 10659
rect 24685 10625 24719 10659
rect 24869 10625 24903 10659
rect 25421 10625 25455 10659
rect 25513 10625 25547 10659
rect 25789 10625 25823 10659
rect 25973 10625 26007 10659
rect 27261 10625 27295 10659
rect 27353 10625 27387 10659
rect 27445 10625 27479 10659
rect 27537 10625 27571 10659
rect 27721 10625 27755 10659
rect 27997 10625 28031 10659
rect 28181 10625 28215 10659
rect 28457 10625 28491 10659
rect 28733 10625 28767 10659
rect 28917 10625 28951 10659
rect 29377 10625 29411 10659
rect 29469 10625 29503 10659
rect 29653 10625 29687 10659
rect 29745 10625 29779 10659
rect 30205 10625 30239 10659
rect 31125 10625 31159 10659
rect 32873 10625 32907 10659
rect 10241 10557 10275 10591
rect 12357 10557 12391 10591
rect 13737 10557 13771 10591
rect 16773 10557 16807 10591
rect 18889 10557 18923 10591
rect 23581 10557 23615 10591
rect 29837 10557 29871 10591
rect 30389 10557 30423 10591
rect 33149 10557 33183 10591
rect 15761 10489 15795 10523
rect 17785 10489 17819 10523
rect 17877 10489 17911 10523
rect 18153 10489 18187 10523
rect 23949 10489 23983 10523
rect 9689 10421 9723 10455
rect 10609 10421 10643 10455
rect 12633 10421 12667 10455
rect 14565 10421 14599 10455
rect 16037 10421 16071 10455
rect 16313 10421 16347 10455
rect 19349 10421 19383 10455
rect 21833 10421 21867 10455
rect 25697 10421 25731 10455
rect 25881 10421 25915 10455
rect 27353 10421 27387 10455
rect 27905 10421 27939 10455
rect 28089 10421 28123 10455
rect 29101 10421 29135 10455
rect 30481 10421 30515 10455
rect 30665 10421 30699 10455
rect 10701 10217 10735 10251
rect 12541 10217 12575 10251
rect 13829 10217 13863 10251
rect 14473 10217 14507 10251
rect 17049 10217 17083 10251
rect 20913 10217 20947 10251
rect 21452 10217 21486 10251
rect 22937 10217 22971 10251
rect 28917 10217 28951 10251
rect 30297 10217 30331 10251
rect 31861 10217 31895 10251
rect 11345 10149 11379 10183
rect 11713 10149 11747 10183
rect 18797 10149 18831 10183
rect 20085 10149 20119 10183
rect 29193 10149 29227 10183
rect 8953 10081 8987 10115
rect 11069 10081 11103 10115
rect 17233 10081 17267 10115
rect 18337 10081 18371 10115
rect 20361 10081 20395 10115
rect 21189 10081 21223 10115
rect 26249 10081 26283 10115
rect 26709 10081 26743 10115
rect 26893 10081 26927 10115
rect 30849 10081 30883 10115
rect 10977 10013 11011 10047
rect 11437 10013 11471 10047
rect 12725 10013 12759 10047
rect 12817 10013 12851 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 13737 10013 13771 10047
rect 13921 10013 13955 10047
rect 16221 10013 16255 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 17325 10013 17359 10047
rect 18429 10013 18463 10047
rect 20453 10013 20487 10047
rect 21004 10013 21038 10047
rect 21097 10013 21131 10047
rect 23765 10013 23799 10047
rect 24041 10013 24075 10047
rect 25329 10013 25363 10047
rect 25697 10013 25731 10047
rect 25789 10013 25823 10047
rect 25973 10013 26007 10047
rect 26341 10013 26375 10047
rect 27169 10013 27203 10047
rect 27353 10013 27387 10047
rect 28917 10013 28951 10047
rect 29009 10013 29043 10047
rect 29285 10013 29319 10047
rect 30205 10013 30239 10047
rect 30389 10015 30423 10049
rect 31125 10013 31159 10047
rect 9229 9945 9263 9979
rect 14105 9945 14139 9979
rect 14289 9945 14323 9979
rect 16497 9945 16531 9979
rect 25421 9945 25455 9979
rect 25513 9945 25547 9979
rect 25881 9945 25915 9979
rect 27031 9945 27065 9979
rect 27261 9945 27295 9979
rect 11897 9877 11931 9911
rect 16773 9877 16807 9911
rect 23029 9877 23063 9911
rect 25145 9877 25179 9911
rect 27537 9877 27571 9911
rect 9321 9673 9355 9707
rect 12541 9673 12575 9707
rect 22201 9673 22235 9707
rect 24041 9673 24075 9707
rect 25789 9673 25823 9707
rect 27997 9673 28031 9707
rect 30205 9673 30239 9707
rect 14657 9605 14691 9639
rect 19809 9605 19843 9639
rect 25421 9605 25455 9639
rect 25605 9605 25639 9639
rect 30297 9605 30331 9639
rect 9505 9537 9539 9571
rect 10149 9537 10183 9571
rect 12173 9537 12207 9571
rect 14565 9537 14599 9571
rect 14749 9537 14783 9571
rect 14933 9537 14967 9571
rect 19533 9537 19567 9571
rect 19717 9537 19751 9571
rect 19901 9537 19935 9571
rect 22109 9537 22143 9571
rect 23029 9537 23063 9571
rect 23305 9537 23339 9571
rect 27997 9537 28031 9571
rect 28181 9537 28215 9571
rect 29561 9537 29595 9571
rect 9873 9469 9907 9503
rect 12265 9469 12299 9503
rect 30389 9469 30423 9503
rect 29837 9401 29871 9435
rect 10885 9333 10919 9367
rect 14381 9333 14415 9367
rect 20085 9333 20119 9367
rect 29745 9333 29779 9367
rect 11529 9129 11563 9163
rect 15301 9129 15335 9163
rect 15945 9129 15979 9163
rect 16957 9129 16991 9163
rect 18429 9129 18463 9163
rect 19073 9129 19107 9163
rect 28457 9129 28491 9163
rect 31309 9129 31343 9163
rect 14749 9061 14783 9095
rect 17877 9061 17911 9095
rect 20269 9061 20303 9095
rect 24409 9061 24443 9095
rect 25237 9061 25271 9095
rect 26157 9061 26191 9095
rect 29193 9061 29227 9095
rect 17233 8993 17267 9027
rect 18613 8993 18647 9027
rect 19625 8993 19659 9027
rect 22109 8993 22143 9027
rect 25053 8993 25087 9027
rect 25697 8993 25731 9027
rect 27353 8993 27387 9027
rect 29837 8993 29871 9027
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 15577 8925 15611 8959
rect 15761 8925 15795 8959
rect 16405 8925 16439 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17049 8925 17083 8959
rect 17141 8925 17175 8959
rect 17325 8925 17359 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 18061 8925 18095 8959
rect 18245 8925 18279 8959
rect 18705 8925 18739 8959
rect 19901 8925 19935 8959
rect 21833 8925 21867 8959
rect 23397 8925 23431 8959
rect 24777 8925 24811 8959
rect 25605 8925 25639 8959
rect 27077 8925 27111 8959
rect 28273 8925 28307 8959
rect 28365 8925 28399 8959
rect 28549 8925 28583 8959
rect 29561 8925 29595 8959
rect 14749 8857 14783 8891
rect 15117 8857 15151 8891
rect 16589 8857 16623 8891
rect 18153 8857 18187 8891
rect 19809 8857 19843 8891
rect 25881 8857 25915 8891
rect 27905 8857 27939 8891
rect 28089 8857 28123 8891
rect 28917 8857 28951 8891
rect 15317 8789 15351 8823
rect 15485 8789 15519 8823
rect 17693 8789 17727 8823
rect 21097 8789 21131 8823
rect 23213 8789 23247 8823
rect 24869 8789 24903 8823
rect 26341 8789 26375 8823
rect 26709 8789 26743 8823
rect 27169 8789 27203 8823
rect 29377 8789 29411 8823
rect 17049 8585 17083 8619
rect 18337 8585 18371 8619
rect 26525 8585 26559 8619
rect 27905 8585 27939 8619
rect 28641 8585 28675 8619
rect 30113 8585 30147 8619
rect 13829 8517 13863 8551
rect 18797 8517 18831 8551
rect 21373 8517 21407 8551
rect 22845 8517 22879 8551
rect 11621 8449 11655 8483
rect 14657 8449 14691 8483
rect 14933 8449 14967 8483
rect 18245 8449 18279 8483
rect 19441 8449 19475 8483
rect 21465 8449 21499 8483
rect 22569 8449 22603 8483
rect 24685 8449 24719 8483
rect 25789 8449 25823 8483
rect 26801 8449 26835 8483
rect 27537 8449 27571 8483
rect 29377 8449 29411 8483
rect 29653 8449 29687 8483
rect 30021 8449 30055 8483
rect 38209 8449 38243 8483
rect 11897 8381 11931 8415
rect 13921 8381 13955 8415
rect 14105 8381 14139 8415
rect 14749 8381 14783 8415
rect 15393 8381 15427 8415
rect 17141 8381 17175 8415
rect 17233 8381 17267 8415
rect 17785 8381 17819 8415
rect 19717 8381 19751 8415
rect 21189 8381 21223 8415
rect 24317 8381 24351 8415
rect 24409 8381 24443 8415
rect 25513 8381 25547 8415
rect 27445 8381 27479 8415
rect 13461 8313 13495 8347
rect 14289 8313 14323 8347
rect 15301 8313 15335 8347
rect 17877 8313 17911 8347
rect 18429 8313 18463 8347
rect 25421 8313 25455 8347
rect 38393 8313 38427 8347
rect 13369 8245 13403 8279
rect 16681 8245 16715 8279
rect 26617 8245 26651 8279
rect 12265 8041 12299 8075
rect 12633 8041 12667 8075
rect 15209 8041 15243 8075
rect 17325 8041 17359 8075
rect 17969 8041 18003 8075
rect 19993 8041 20027 8075
rect 23581 8041 23615 8075
rect 15577 7905 15611 7939
rect 20637 7905 20671 7939
rect 26249 7905 26283 7939
rect 26525 7905 26559 7939
rect 28089 7905 28123 7939
rect 12425 7833 12459 7867
rect 12549 7837 12583 7871
rect 12909 7837 12943 7871
rect 13185 7837 13219 7871
rect 14197 7837 14231 7871
rect 14473 7837 14507 7871
rect 17601 7837 17635 7871
rect 18705 7837 18739 7871
rect 18981 7837 19015 7871
rect 20177 7837 20211 7871
rect 20913 7837 20947 7871
rect 23489 7837 23523 7871
rect 28365 7837 28399 7871
rect 15853 7769 15887 7803
rect 17509 7769 17543 7803
rect 13921 7701 13955 7735
rect 21649 7701 21683 7735
rect 27997 7701 28031 7735
rect 29101 7701 29135 7735
rect 16037 7497 16071 7531
rect 27353 7497 27387 7531
rect 16221 7361 16255 7395
rect 17601 7361 17635 7395
rect 27261 7361 27295 7395
rect 17325 7293 17359 7327
rect 18337 7157 18371 7191
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 15470 37408 15476 37460
rect 15528 37448 15534 37460
rect 15749 37451 15807 37457
rect 15749 37448 15761 37451
rect 15528 37420 15761 37448
rect 15528 37408 15534 37420
rect 15749 37417 15761 37420
rect 15795 37417 15807 37451
rect 15749 37411 15807 37417
rect 17402 37408 17408 37460
rect 17460 37448 17466 37460
rect 17681 37451 17739 37457
rect 17681 37448 17693 37451
rect 17460 37420 17693 37448
rect 17460 37408 17466 37420
rect 17681 37417 17693 37420
rect 17727 37417 17739 37451
rect 17681 37411 17739 37417
rect 19334 37408 19340 37460
rect 19392 37448 19398 37460
rect 19613 37451 19671 37457
rect 19613 37448 19625 37451
rect 19392 37420 19625 37448
rect 19392 37408 19398 37420
rect 19613 37417 19625 37420
rect 19659 37417 19671 37451
rect 19613 37411 19671 37417
rect 21910 37408 21916 37460
rect 21968 37448 21974 37460
rect 22097 37451 22155 37457
rect 22097 37448 22109 37451
rect 21968 37420 22109 37448
rect 21968 37408 21974 37420
rect 22097 37417 22109 37420
rect 22143 37417 22155 37451
rect 22097 37411 22155 37417
rect 15654 37136 15660 37188
rect 15712 37136 15718 37188
rect 17310 37136 17316 37188
rect 17368 37176 17374 37188
rect 17589 37179 17647 37185
rect 17589 37176 17601 37179
rect 17368 37148 17601 37176
rect 17368 37136 17374 37148
rect 17589 37145 17601 37148
rect 17635 37145 17647 37179
rect 17589 37139 17647 37145
rect 19518 37136 19524 37188
rect 19576 37136 19582 37188
rect 22370 37136 22376 37188
rect 22428 37136 22434 37188
rect 1104 37018 38824 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 38824 33754
rect 1104 33680 38824 33702
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 38824 31578
rect 1104 31504 38824 31526
rect 7558 31220 7564 31272
rect 7616 31220 7622 31272
rect 8202 31084 8208 31136
rect 8260 31084 8266 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 7285 30923 7343 30929
rect 7285 30889 7297 30923
rect 7331 30920 7343 30923
rect 7558 30920 7564 30932
rect 7331 30892 7564 30920
rect 7331 30889 7343 30892
rect 7285 30883 7343 30889
rect 7558 30880 7564 30892
rect 7616 30880 7622 30932
rect 8202 30880 8208 30932
rect 8260 30880 8266 30932
rect 6825 30787 6883 30793
rect 6825 30753 6837 30787
rect 6871 30784 6883 30787
rect 7377 30787 7435 30793
rect 6871 30756 7236 30784
rect 6871 30753 6883 30756
rect 6825 30747 6883 30753
rect 7208 30728 7236 30756
rect 7377 30753 7389 30787
rect 7423 30784 7435 30787
rect 7834 30784 7840 30796
rect 7423 30756 7840 30784
rect 7423 30753 7435 30756
rect 7377 30747 7435 30753
rect 7834 30744 7840 30756
rect 7892 30784 7898 30796
rect 8113 30787 8171 30793
rect 8113 30784 8125 30787
rect 7892 30756 8125 30784
rect 7892 30744 7898 30756
rect 8113 30753 8125 30756
rect 8159 30753 8171 30787
rect 8113 30747 8171 30753
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30716 6791 30719
rect 7101 30719 7159 30725
rect 7101 30716 7113 30719
rect 6779 30688 7113 30716
rect 6779 30685 6791 30688
rect 6733 30679 6791 30685
rect 7101 30685 7113 30688
rect 7147 30685 7159 30719
rect 7101 30679 7159 30685
rect 7116 30592 7144 30679
rect 7190 30676 7196 30728
rect 7248 30676 7254 30728
rect 7466 30676 7472 30728
rect 7524 30676 7530 30728
rect 8220 30725 8248 30880
rect 8205 30719 8263 30725
rect 8205 30685 8217 30719
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30716 8447 30719
rect 8435 30688 8524 30716
rect 8435 30685 8447 30688
rect 8389 30679 8447 30685
rect 8496 30592 8524 30688
rect 10594 30676 10600 30728
rect 10652 30676 10658 30728
rect 11790 30676 11796 30728
rect 11848 30676 11854 30728
rect 12250 30676 12256 30728
rect 12308 30676 12314 30728
rect 15562 30676 15568 30728
rect 15620 30716 15626 30728
rect 16945 30719 17003 30725
rect 16945 30716 16957 30719
rect 15620 30688 16957 30716
rect 15620 30676 15626 30688
rect 16945 30685 16957 30688
rect 16991 30685 17003 30719
rect 16945 30679 17003 30685
rect 6362 30540 6368 30592
rect 6420 30540 6426 30592
rect 7098 30540 7104 30592
rect 7156 30540 7162 30592
rect 8386 30540 8392 30592
rect 8444 30540 8450 30592
rect 8478 30540 8484 30592
rect 8536 30540 8542 30592
rect 10778 30540 10784 30592
rect 10836 30540 10842 30592
rect 11238 30540 11244 30592
rect 11296 30540 11302 30592
rect 12894 30540 12900 30592
rect 12952 30540 12958 30592
rect 17586 30540 17592 30592
rect 17644 30540 17650 30592
rect 1104 30490 38824 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 38824 30490
rect 1104 30416 38824 30438
rect 7466 30336 7472 30388
rect 7524 30336 7530 30388
rect 10594 30336 10600 30388
rect 10652 30376 10658 30388
rect 10781 30379 10839 30385
rect 10781 30376 10793 30379
rect 10652 30348 10793 30376
rect 10652 30336 10658 30348
rect 10781 30345 10793 30348
rect 10827 30345 10839 30379
rect 10781 30339 10839 30345
rect 11333 30379 11391 30385
rect 11333 30345 11345 30379
rect 11379 30376 11391 30379
rect 12250 30376 12256 30388
rect 11379 30348 12256 30376
rect 11379 30345 11391 30348
rect 11333 30339 11391 30345
rect 12250 30336 12256 30348
rect 12308 30336 12314 30388
rect 8386 30268 8392 30320
rect 8444 30308 8450 30320
rect 8582 30311 8640 30317
rect 8582 30308 8594 30311
rect 8444 30280 8594 30308
rect 8444 30268 8450 30280
rect 8582 30277 8594 30280
rect 8628 30277 8640 30311
rect 8582 30271 8640 30277
rect 10321 30311 10379 30317
rect 10321 30277 10333 30311
rect 10367 30308 10379 30311
rect 11238 30308 11244 30320
rect 10367 30280 11244 30308
rect 10367 30277 10379 30280
rect 10321 30271 10379 30277
rect 11238 30268 11244 30280
rect 11296 30268 11302 30320
rect 11790 30268 11796 30320
rect 11848 30268 11854 30320
rect 6362 30200 6368 30252
rect 6420 30240 6426 30252
rect 6549 30243 6607 30249
rect 6549 30240 6561 30243
rect 6420 30212 6561 30240
rect 6420 30200 6426 30212
rect 6549 30209 6561 30212
rect 6595 30209 6607 30243
rect 6549 30203 6607 30209
rect 8849 30243 8907 30249
rect 8849 30209 8861 30243
rect 8895 30209 8907 30243
rect 8849 30203 8907 30209
rect 10873 30243 10931 30249
rect 10873 30209 10885 30243
rect 10919 30240 10931 30243
rect 11146 30240 11152 30252
rect 10919 30212 11152 30240
rect 10919 30209 10931 30212
rect 10873 30203 10931 30209
rect 8864 30172 8892 30203
rect 11146 30200 11152 30212
rect 11204 30240 11210 30252
rect 11808 30240 11836 30268
rect 11204 30212 11836 30240
rect 11204 30200 11210 30212
rect 12710 30200 12716 30252
rect 12768 30240 12774 30252
rect 13153 30243 13211 30249
rect 13153 30240 13165 30243
rect 12768 30212 13165 30240
rect 12768 30200 12774 30212
rect 13153 30209 13165 30212
rect 13199 30209 13211 30243
rect 13153 30203 13211 30209
rect 13722 30200 13728 30252
rect 13780 30240 13786 30252
rect 15749 30243 15807 30249
rect 15749 30240 15761 30243
rect 13780 30212 15761 30240
rect 13780 30200 13786 30212
rect 15749 30209 15761 30212
rect 15795 30209 15807 30243
rect 15749 30203 15807 30209
rect 11054 30172 11060 30184
rect 8864 30144 11060 30172
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 12434 30132 12440 30184
rect 12492 30132 12498 30184
rect 12897 30175 12955 30181
rect 12897 30141 12909 30175
rect 12943 30141 12955 30175
rect 15562 30172 15568 30184
rect 12897 30135 12955 30141
rect 14292 30144 15568 30172
rect 10689 30107 10747 30113
rect 10689 30073 10701 30107
rect 10735 30104 10747 30107
rect 10735 30076 11192 30104
rect 10735 30073 10747 30076
rect 10689 30067 10747 30073
rect 7193 30039 7251 30045
rect 7193 30005 7205 30039
rect 7239 30036 7251 30039
rect 7374 30036 7380 30048
rect 7239 30008 7380 30036
rect 7239 30005 7251 30008
rect 7193 29999 7251 30005
rect 7374 29996 7380 30008
rect 7432 29996 7438 30048
rect 11164 30045 11192 30076
rect 11149 30039 11207 30045
rect 11149 30005 11161 30039
rect 11195 30036 11207 30039
rect 11885 30039 11943 30045
rect 11885 30036 11897 30039
rect 11195 30008 11897 30036
rect 11195 30005 11207 30008
rect 11149 29999 11207 30005
rect 11885 30005 11897 30008
rect 11931 30005 11943 30039
rect 11885 29999 11943 30005
rect 12342 29996 12348 30048
rect 12400 30036 12406 30048
rect 12912 30036 12940 30135
rect 14292 30113 14320 30144
rect 15562 30132 15568 30144
rect 15620 30132 15626 30184
rect 15764 30172 15792 30203
rect 17586 30200 17592 30252
rect 17644 30240 17650 30252
rect 19593 30243 19651 30249
rect 19593 30240 19605 30243
rect 17644 30212 19605 30240
rect 17644 30200 17650 30212
rect 19593 30209 19605 30212
rect 19639 30209 19651 30243
rect 19593 30203 19651 30209
rect 19337 30175 19395 30181
rect 15764 30144 18184 30172
rect 14277 30107 14335 30113
rect 14277 30073 14289 30107
rect 14323 30073 14335 30107
rect 14277 30067 14335 30073
rect 18156 30048 18184 30144
rect 19337 30141 19349 30175
rect 19383 30141 19395 30175
rect 20901 30175 20959 30181
rect 20901 30172 20913 30175
rect 19337 30135 19395 30141
rect 20732 30144 20913 30172
rect 14090 30036 14096 30048
rect 12400 30008 14096 30036
rect 12400 29996 12406 30008
rect 14090 29996 14096 30008
rect 14148 29996 14154 30048
rect 15657 30039 15715 30045
rect 15657 30005 15669 30039
rect 15703 30036 15715 30039
rect 15746 30036 15752 30048
rect 15703 30008 15752 30036
rect 15703 30005 15715 30008
rect 15657 29999 15715 30005
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 18138 29996 18144 30048
rect 18196 29996 18202 30048
rect 19352 30036 19380 30135
rect 20732 30113 20760 30144
rect 20901 30141 20913 30144
rect 20947 30141 20959 30175
rect 20901 30135 20959 30141
rect 20717 30107 20775 30113
rect 20717 30073 20729 30107
rect 20763 30073 20775 30107
rect 20717 30067 20775 30073
rect 19978 30036 19984 30048
rect 19352 30008 19984 30036
rect 19978 29996 19984 30008
rect 20036 29996 20042 30048
rect 21542 29996 21548 30048
rect 21600 29996 21606 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 11977 29835 12035 29841
rect 11977 29801 11989 29835
rect 12023 29832 12035 29835
rect 12434 29832 12440 29844
rect 12023 29804 12440 29832
rect 12023 29801 12035 29804
rect 11977 29795 12035 29801
rect 12434 29792 12440 29804
rect 12492 29792 12498 29844
rect 12621 29835 12679 29841
rect 12621 29801 12633 29835
rect 12667 29832 12679 29835
rect 12710 29832 12716 29844
rect 12667 29804 12716 29832
rect 12667 29801 12679 29804
rect 12621 29795 12679 29801
rect 12710 29792 12716 29804
rect 12768 29792 12774 29844
rect 17586 29832 17592 29844
rect 13188 29804 17592 29832
rect 7834 29724 7840 29776
rect 7892 29724 7898 29776
rect 7653 29699 7711 29705
rect 7653 29665 7665 29699
rect 7699 29696 7711 29699
rect 12253 29699 12311 29705
rect 7699 29668 8340 29696
rect 7699 29665 7711 29668
rect 7653 29659 7711 29665
rect 8312 29640 8340 29668
rect 12253 29665 12265 29699
rect 12299 29696 12311 29699
rect 12894 29696 12900 29708
rect 12299 29668 12900 29696
rect 12299 29665 12311 29668
rect 12253 29659 12311 29665
rect 12894 29656 12900 29668
rect 12952 29656 12958 29708
rect 5810 29588 5816 29640
rect 5868 29588 5874 29640
rect 5997 29631 6055 29637
rect 5997 29597 6009 29631
rect 6043 29597 6055 29631
rect 5997 29591 6055 29597
rect 6181 29631 6239 29637
rect 6181 29597 6193 29631
rect 6227 29628 6239 29631
rect 6270 29628 6276 29640
rect 6227 29600 6276 29628
rect 6227 29597 6239 29600
rect 6181 29591 6239 29597
rect 6012 29560 6040 29591
rect 6270 29588 6276 29600
rect 6328 29588 6334 29640
rect 7374 29588 7380 29640
rect 7432 29637 7438 29640
rect 7432 29628 7444 29637
rect 7745 29631 7803 29637
rect 7432 29600 7477 29628
rect 7432 29591 7444 29600
rect 7745 29597 7757 29631
rect 7791 29597 7803 29631
rect 7745 29591 7803 29597
rect 8021 29631 8079 29637
rect 8021 29597 8033 29631
rect 8067 29597 8079 29631
rect 8021 29591 8079 29597
rect 7432 29588 7438 29591
rect 6086 29560 6092 29572
rect 6012 29532 6092 29560
rect 6086 29520 6092 29532
rect 6144 29560 6150 29572
rect 7190 29560 7196 29572
rect 6144 29532 7196 29560
rect 6144 29520 6150 29532
rect 7190 29520 7196 29532
rect 7248 29560 7254 29572
rect 7760 29560 7788 29591
rect 7248 29532 7788 29560
rect 7248 29520 7254 29532
rect 5261 29495 5319 29501
rect 5261 29461 5273 29495
rect 5307 29492 5319 29495
rect 5350 29492 5356 29504
rect 5307 29464 5356 29492
rect 5307 29461 5319 29464
rect 5261 29455 5319 29461
rect 5350 29452 5356 29464
rect 5408 29452 5414 29504
rect 5994 29452 6000 29504
rect 6052 29452 6058 29504
rect 6273 29495 6331 29501
rect 6273 29461 6285 29495
rect 6319 29492 6331 29495
rect 7098 29492 7104 29504
rect 6319 29464 7104 29492
rect 6319 29461 6331 29464
rect 6273 29455 6331 29461
rect 7098 29452 7104 29464
rect 7156 29492 7162 29504
rect 8036 29492 8064 29591
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 8941 29631 8999 29637
rect 8941 29597 8953 29631
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29628 9183 29631
rect 9674 29628 9680 29640
rect 9171 29600 9680 29628
rect 9171 29597 9183 29600
rect 9125 29591 9183 29597
rect 8478 29520 8484 29572
rect 8536 29560 8542 29572
rect 8956 29560 8984 29591
rect 9674 29588 9680 29600
rect 9732 29588 9738 29640
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 10864 29631 10922 29637
rect 10864 29597 10876 29631
rect 10910 29597 10922 29631
rect 10864 29591 10922 29597
rect 12345 29631 12403 29637
rect 12345 29597 12357 29631
rect 12391 29628 12403 29631
rect 13188 29628 13216 29804
rect 17586 29792 17592 29804
rect 17644 29832 17650 29844
rect 17644 29804 20300 29832
rect 17644 29792 17650 29804
rect 20272 29773 20300 29804
rect 20257 29767 20315 29773
rect 20257 29733 20269 29767
rect 20303 29733 20315 29767
rect 20257 29727 20315 29733
rect 13722 29656 13728 29708
rect 13780 29656 13786 29708
rect 14090 29656 14096 29708
rect 14148 29696 14154 29708
rect 14461 29699 14519 29705
rect 14461 29696 14473 29699
rect 14148 29668 14473 29696
rect 14148 29656 14154 29668
rect 14461 29665 14473 29668
rect 14507 29696 14519 29699
rect 16577 29699 16635 29705
rect 16577 29696 16589 29699
rect 14507 29668 16589 29696
rect 14507 29665 14519 29668
rect 14461 29659 14519 29665
rect 16577 29665 16589 29668
rect 16623 29665 16635 29699
rect 20165 29699 20223 29705
rect 20165 29696 20177 29699
rect 16577 29659 16635 29665
rect 19904 29668 20177 29696
rect 12391 29600 13216 29628
rect 12391 29597 12403 29600
rect 12345 29591 12403 29597
rect 9582 29560 9588 29572
rect 8536 29532 9588 29560
rect 8536 29520 8542 29532
rect 9582 29520 9588 29532
rect 9640 29520 9646 29572
rect 7156 29464 8064 29492
rect 7156 29452 7162 29464
rect 8662 29452 8668 29504
rect 8720 29492 8726 29504
rect 9033 29495 9091 29501
rect 9033 29492 9045 29495
rect 8720 29464 9045 29492
rect 8720 29452 8726 29464
rect 9033 29461 9045 29464
rect 9079 29461 9091 29495
rect 10612 29492 10640 29591
rect 10778 29520 10784 29572
rect 10836 29560 10842 29572
rect 10888 29560 10916 29591
rect 13262 29588 13268 29640
rect 13320 29628 13326 29640
rect 13740 29628 13768 29656
rect 13320 29600 13768 29628
rect 13320 29588 13326 29600
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 19904 29637 19932 29668
rect 20165 29665 20177 29668
rect 20211 29665 20223 29699
rect 20165 29659 20223 29665
rect 20625 29699 20683 29705
rect 20625 29665 20637 29699
rect 20671 29696 20683 29699
rect 20671 29668 20944 29696
rect 20671 29665 20683 29668
rect 20625 29659 20683 29665
rect 19889 29631 19947 29637
rect 15804 29600 15870 29628
rect 15804 29588 15810 29600
rect 19889 29597 19901 29631
rect 19935 29597 19947 29631
rect 19889 29591 19947 29597
rect 19978 29588 19984 29640
rect 20036 29628 20042 29640
rect 20809 29631 20867 29637
rect 20809 29628 20821 29631
rect 20036 29600 20821 29628
rect 20036 29588 20042 29600
rect 20809 29597 20821 29600
rect 20855 29597 20867 29631
rect 20916 29628 20944 29668
rect 21076 29631 21134 29637
rect 21076 29628 21088 29631
rect 20916 29600 21088 29628
rect 20809 29591 20867 29597
rect 21076 29597 21088 29600
rect 21122 29628 21134 29631
rect 21542 29628 21548 29640
rect 21122 29600 21548 29628
rect 21122 29597 21134 29600
rect 21076 29591 21134 29597
rect 21542 29588 21548 29600
rect 21600 29588 21606 29640
rect 10836 29532 10916 29560
rect 10836 29520 10842 29532
rect 14734 29520 14740 29572
rect 14792 29520 14798 29572
rect 16482 29520 16488 29572
rect 16540 29520 16546 29572
rect 16850 29520 16856 29572
rect 16908 29520 16914 29572
rect 17586 29520 17592 29572
rect 17644 29520 17650 29572
rect 18601 29563 18659 29569
rect 18601 29529 18613 29563
rect 18647 29529 18659 29563
rect 18601 29523 18659 29529
rect 11054 29492 11060 29504
rect 10612 29464 11060 29492
rect 9033 29455 9091 29461
rect 11054 29452 11060 29464
rect 11112 29452 11118 29504
rect 13354 29452 13360 29504
rect 13412 29452 13418 29504
rect 17034 29452 17040 29504
rect 17092 29492 17098 29504
rect 18616 29492 18644 29523
rect 17092 29464 18644 29492
rect 20073 29495 20131 29501
rect 17092 29452 17098 29464
rect 20073 29461 20085 29495
rect 20119 29492 20131 29495
rect 20438 29492 20444 29504
rect 20119 29464 20444 29492
rect 20119 29461 20131 29464
rect 20073 29455 20131 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 22186 29452 22192 29504
rect 22244 29452 22250 29504
rect 1104 29402 38824 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 38824 29402
rect 1104 29328 38824 29350
rect 4801 29291 4859 29297
rect 4801 29257 4813 29291
rect 4847 29288 4859 29291
rect 5810 29288 5816 29300
rect 4847 29260 5816 29288
rect 4847 29257 4859 29260
rect 4801 29251 4859 29257
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 5994 29248 6000 29300
rect 6052 29248 6058 29300
rect 9674 29248 9680 29300
rect 9732 29248 9738 29300
rect 11146 29248 11152 29300
rect 11204 29248 11210 29300
rect 14734 29248 14740 29300
rect 14792 29288 14798 29300
rect 15013 29291 15071 29297
rect 15013 29288 15025 29291
rect 14792 29260 15025 29288
rect 14792 29248 14798 29260
rect 15013 29257 15025 29260
rect 15059 29257 15071 29291
rect 15013 29251 15071 29257
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 16761 29291 16819 29297
rect 15252 29260 16712 29288
rect 15252 29248 15258 29260
rect 5925 29155 5983 29161
rect 5925 29121 5937 29155
rect 5971 29152 5983 29155
rect 6012 29152 6040 29248
rect 6362 29220 6368 29232
rect 6196 29192 6368 29220
rect 6196 29161 6224 29192
rect 6362 29180 6368 29192
rect 6420 29220 6426 29232
rect 6420 29192 8340 29220
rect 6420 29180 6426 29192
rect 8312 29164 8340 29192
rect 9784 29192 11100 29220
rect 5971 29124 6040 29152
rect 6181 29155 6239 29161
rect 5971 29121 5983 29124
rect 5925 29115 5983 29121
rect 6181 29121 6193 29155
rect 6227 29121 6239 29155
rect 6181 29115 6239 29121
rect 6270 29112 6276 29164
rect 6328 29112 6334 29164
rect 6638 29112 6644 29164
rect 6696 29152 6702 29164
rect 7101 29155 7159 29161
rect 7101 29152 7113 29155
rect 6696 29124 7113 29152
rect 6696 29112 6702 29124
rect 7101 29121 7113 29124
rect 7147 29121 7159 29155
rect 7101 29115 7159 29121
rect 8294 29112 8300 29164
rect 8352 29112 8358 29164
rect 8564 29155 8622 29161
rect 8564 29121 8576 29155
rect 8610 29152 8622 29155
rect 8938 29152 8944 29164
rect 8610 29124 8944 29152
rect 8610 29121 8622 29124
rect 8564 29115 8622 29121
rect 8938 29112 8944 29124
rect 8996 29112 9002 29164
rect 9784 29161 9812 29192
rect 10042 29161 10048 29164
rect 9769 29155 9827 29161
rect 9769 29121 9781 29155
rect 9815 29121 9827 29155
rect 10036 29152 10048 29161
rect 10003 29124 10048 29152
rect 9769 29115 9827 29121
rect 10036 29115 10048 29124
rect 10042 29112 10048 29115
rect 10100 29112 10106 29164
rect 6288 29084 6316 29112
rect 11072 29096 11100 29192
rect 13354 29180 13360 29232
rect 13412 29180 13418 29232
rect 15102 29180 15108 29232
rect 15160 29220 15166 29232
rect 15381 29223 15439 29229
rect 15381 29220 15393 29223
rect 15160 29192 15393 29220
rect 15160 29180 15166 29192
rect 15381 29189 15393 29192
rect 15427 29189 15439 29223
rect 16482 29220 16488 29232
rect 15381 29183 15439 29189
rect 15488 29192 16488 29220
rect 15194 29112 15200 29164
rect 15252 29112 15258 29164
rect 15289 29155 15347 29161
rect 15289 29121 15301 29155
rect 15335 29152 15347 29155
rect 15488 29152 15516 29192
rect 16482 29180 16488 29192
rect 16540 29180 16546 29232
rect 16684 29220 16712 29260
rect 16761 29257 16773 29291
rect 16807 29288 16819 29291
rect 16850 29288 16856 29300
rect 16807 29260 16856 29288
rect 16807 29257 16819 29260
rect 16761 29251 16819 29257
rect 16850 29248 16856 29260
rect 16908 29248 16914 29300
rect 17494 29288 17500 29300
rect 16960 29260 17500 29288
rect 16960 29220 16988 29260
rect 17494 29248 17500 29260
rect 17552 29248 17558 29300
rect 17586 29248 17592 29300
rect 17644 29288 17650 29300
rect 17681 29291 17739 29297
rect 17681 29288 17693 29291
rect 17644 29260 17693 29288
rect 17644 29248 17650 29260
rect 17681 29257 17693 29260
rect 17727 29257 17739 29291
rect 19978 29288 19984 29300
rect 17681 29251 17739 29257
rect 18248 29260 19984 29288
rect 18046 29220 18052 29232
rect 16684 29192 16988 29220
rect 16960 29161 16988 29192
rect 17328 29192 18052 29220
rect 15335 29124 15516 29152
rect 15565 29155 15623 29161
rect 15335 29121 15347 29124
rect 15289 29115 15347 29121
rect 15565 29121 15577 29155
rect 15611 29152 15623 29155
rect 16945 29155 17003 29161
rect 15611 29124 15792 29152
rect 15611 29121 15623 29124
rect 15565 29115 15623 29121
rect 6365 29087 6423 29093
rect 6365 29084 6377 29087
rect 6288 29056 6377 29084
rect 6365 29053 6377 29056
rect 6411 29053 6423 29087
rect 6365 29047 6423 29053
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 6917 29087 6975 29093
rect 6917 29084 6929 29087
rect 6604 29056 6929 29084
rect 6604 29044 6610 29056
rect 6917 29053 6929 29056
rect 6963 29053 6975 29087
rect 6917 29047 6975 29053
rect 7377 29087 7435 29093
rect 7377 29053 7389 29087
rect 7423 29084 7435 29087
rect 7423 29056 7512 29084
rect 7423 29053 7435 29056
rect 7377 29047 7435 29053
rect 6454 28976 6460 29028
rect 6512 29016 6518 29028
rect 7193 29019 7251 29025
rect 7193 29016 7205 29019
rect 6512 28988 7205 29016
rect 6512 28976 6518 28988
rect 7193 28985 7205 28988
rect 7239 28985 7251 29019
rect 7193 28979 7251 28985
rect 7484 28960 7512 29056
rect 8018 29044 8024 29096
rect 8076 29044 8082 29096
rect 11054 29044 11060 29096
rect 11112 29084 11118 29096
rect 12342 29084 12348 29096
rect 11112 29056 12348 29084
rect 11112 29044 11118 29056
rect 12342 29044 12348 29056
rect 12400 29044 12406 29096
rect 12618 29044 12624 29096
rect 12676 29044 12682 29096
rect 14093 29087 14151 29093
rect 14093 29053 14105 29087
rect 14139 29084 14151 29087
rect 14550 29084 14556 29096
rect 14139 29056 14556 29084
rect 14139 29053 14151 29056
rect 14093 29047 14151 29053
rect 14550 29044 14556 29056
rect 14608 29084 14614 29096
rect 14829 29087 14887 29093
rect 14829 29084 14841 29087
rect 14608 29056 14841 29084
rect 14608 29044 14614 29056
rect 14829 29053 14841 29056
rect 14875 29053 14887 29087
rect 14829 29047 14887 29053
rect 15764 29084 15792 29124
rect 16945 29121 16957 29155
rect 16991 29121 17003 29155
rect 16945 29115 17003 29121
rect 17034 29112 17040 29164
rect 17092 29112 17098 29164
rect 17126 29112 17132 29164
rect 17184 29112 17190 29164
rect 17328 29161 17356 29192
rect 18046 29180 18052 29192
rect 18104 29180 18110 29232
rect 18248 29161 18276 29260
rect 19978 29248 19984 29260
rect 20036 29248 20042 29300
rect 19518 29180 19524 29232
rect 19576 29180 19582 29232
rect 17313 29155 17371 29161
rect 17313 29152 17325 29155
rect 17236 29124 17325 29152
rect 17236 29084 17264 29124
rect 17313 29121 17325 29124
rect 17359 29121 17371 29155
rect 17313 29115 17371 29121
rect 17589 29155 17647 29161
rect 17589 29121 17601 29155
rect 17635 29121 17647 29155
rect 17589 29115 17647 29121
rect 18233 29155 18291 29161
rect 18233 29121 18245 29155
rect 18279 29121 18291 29155
rect 18233 29115 18291 29121
rect 15764 29056 17264 29084
rect 14182 28976 14188 29028
rect 14240 29016 14246 29028
rect 15764 29016 15792 29056
rect 17494 29044 17500 29096
rect 17552 29044 17558 29096
rect 14240 28988 15792 29016
rect 14240 28976 14246 28988
rect 5534 28908 5540 28960
rect 5592 28948 5598 28960
rect 6638 28948 6644 28960
rect 5592 28920 6644 28948
rect 5592 28908 5598 28920
rect 6638 28908 6644 28920
rect 6696 28908 6702 28960
rect 7282 28908 7288 28960
rect 7340 28908 7346 28960
rect 7466 28908 7472 28960
rect 7524 28908 7530 28960
rect 14274 28908 14280 28960
rect 14332 28908 14338 28960
rect 17512 28948 17540 29044
rect 17604 29016 17632 29115
rect 18138 29044 18144 29096
rect 18196 29044 18202 29096
rect 18506 29044 18512 29096
rect 18564 29084 18570 29096
rect 20257 29087 20315 29093
rect 20257 29084 20269 29087
rect 18564 29056 20269 29084
rect 18564 29044 18570 29056
rect 20257 29053 20269 29056
rect 20303 29053 20315 29087
rect 20257 29047 20315 29053
rect 18156 29016 18184 29044
rect 17604 28988 18184 29016
rect 17954 28948 17960 28960
rect 17512 28920 17960 28948
rect 17954 28908 17960 28920
rect 18012 28908 18018 28960
rect 18230 28908 18236 28960
rect 18288 28948 18294 28960
rect 18490 28951 18548 28957
rect 18490 28948 18502 28951
rect 18288 28920 18502 28948
rect 18288 28908 18294 28920
rect 18490 28917 18502 28920
rect 18536 28917 18548 28951
rect 18490 28911 18548 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 5353 28747 5411 28753
rect 5353 28713 5365 28747
rect 5399 28744 5411 28747
rect 6546 28744 6552 28756
rect 5399 28716 6552 28744
rect 5399 28713 5411 28716
rect 5353 28707 5411 28713
rect 6546 28704 6552 28716
rect 6604 28704 6610 28756
rect 7745 28747 7803 28753
rect 7745 28713 7757 28747
rect 7791 28744 7803 28747
rect 8018 28744 8024 28756
rect 7791 28716 8024 28744
rect 7791 28713 7803 28716
rect 7745 28707 7803 28713
rect 5813 28679 5871 28685
rect 5813 28645 5825 28679
rect 5859 28645 5871 28679
rect 5813 28639 5871 28645
rect 5123 28611 5181 28617
rect 5123 28577 5135 28611
rect 5169 28608 5181 28611
rect 5534 28608 5540 28620
rect 5169 28580 5540 28608
rect 5169 28577 5181 28580
rect 5123 28571 5181 28577
rect 5534 28568 5540 28580
rect 5592 28608 5598 28620
rect 5684 28611 5742 28617
rect 5684 28608 5696 28611
rect 5592 28580 5696 28608
rect 5592 28568 5598 28580
rect 5684 28577 5696 28580
rect 5730 28577 5742 28611
rect 5684 28571 5742 28577
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28540 5043 28543
rect 5261 28543 5319 28549
rect 5031 28512 5212 28540
rect 5031 28509 5043 28512
rect 4985 28503 5043 28509
rect 5184 28404 5212 28512
rect 5261 28509 5273 28543
rect 5307 28509 5319 28543
rect 5261 28503 5319 28509
rect 5276 28472 5304 28503
rect 5350 28500 5356 28552
rect 5408 28540 5414 28552
rect 5445 28543 5503 28549
rect 5445 28540 5457 28543
rect 5408 28512 5457 28540
rect 5408 28500 5414 28512
rect 5445 28509 5457 28512
rect 5491 28540 5503 28543
rect 5828 28540 5856 28639
rect 5905 28611 5963 28617
rect 5905 28577 5917 28611
rect 5951 28577 5963 28611
rect 5905 28571 5963 28577
rect 5491 28512 5856 28540
rect 5920 28540 5948 28571
rect 6086 28568 6092 28620
rect 6144 28568 6150 28620
rect 6362 28568 6368 28620
rect 6420 28568 6426 28620
rect 7760 28540 7788 28707
rect 8018 28704 8024 28716
rect 8076 28704 8082 28756
rect 8938 28704 8944 28756
rect 8996 28704 9002 28756
rect 12618 28704 12624 28756
rect 12676 28744 12682 28756
rect 12805 28747 12863 28753
rect 12805 28744 12817 28747
rect 12676 28716 12817 28744
rect 12676 28704 12682 28716
rect 12805 28713 12817 28716
rect 12851 28713 12863 28747
rect 12805 28707 12863 28713
rect 18230 28704 18236 28756
rect 18288 28704 18294 28756
rect 18322 28704 18328 28756
rect 18380 28744 18386 28756
rect 19337 28747 19395 28753
rect 18380 28716 19288 28744
rect 18380 28704 18386 28716
rect 8665 28679 8723 28685
rect 8665 28645 8677 28679
rect 8711 28645 8723 28679
rect 13262 28676 13268 28688
rect 8665 28639 8723 28645
rect 12636 28648 13268 28676
rect 8680 28608 8708 28639
rect 9493 28611 9551 28617
rect 9493 28608 9505 28611
rect 8680 28580 9505 28608
rect 9493 28577 9505 28580
rect 9539 28577 9551 28611
rect 9493 28571 9551 28577
rect 9582 28568 9588 28620
rect 9640 28608 9646 28620
rect 9640 28580 9904 28608
rect 9640 28568 9646 28580
rect 5920 28512 7788 28540
rect 8573 28543 8631 28549
rect 5491 28509 5503 28512
rect 5445 28503 5503 28509
rect 5537 28475 5595 28481
rect 5537 28472 5549 28475
rect 5276 28444 5549 28472
rect 5537 28441 5549 28444
rect 5583 28472 5595 28475
rect 5810 28472 5816 28484
rect 5583 28444 5816 28472
rect 5583 28441 5595 28444
rect 5537 28435 5595 28441
rect 5810 28432 5816 28444
rect 5868 28432 5874 28484
rect 6012 28404 6040 28512
rect 8573 28509 8585 28543
rect 8619 28540 8631 28543
rect 8662 28540 8668 28552
rect 8619 28512 8668 28540
rect 8619 28509 8631 28512
rect 8573 28503 8631 28509
rect 8662 28500 8668 28512
rect 8720 28500 8726 28552
rect 8757 28543 8815 28549
rect 8757 28509 8769 28543
rect 8803 28540 8815 28543
rect 8803 28512 9628 28540
rect 8803 28509 8815 28512
rect 8757 28503 8815 28509
rect 6638 28481 6644 28484
rect 6632 28435 6644 28481
rect 6638 28432 6644 28435
rect 6696 28432 6702 28484
rect 9600 28416 9628 28512
rect 9674 28500 9680 28552
rect 9732 28500 9738 28552
rect 9876 28549 9904 28580
rect 12342 28568 12348 28620
rect 12400 28568 12406 28620
rect 12636 28549 12664 28648
rect 13262 28636 13268 28648
rect 13320 28636 13326 28688
rect 18506 28676 18512 28688
rect 16408 28648 18512 28676
rect 16408 28620 16436 28648
rect 18506 28636 18512 28648
rect 18564 28636 18570 28688
rect 13096 28580 14320 28608
rect 13096 28549 13124 28580
rect 14292 28552 14320 28580
rect 16390 28568 16396 28620
rect 16448 28568 16454 28620
rect 16669 28611 16727 28617
rect 16669 28577 16681 28611
rect 16715 28608 16727 28611
rect 16758 28608 16764 28620
rect 16715 28580 16764 28608
rect 16715 28577 16727 28580
rect 16669 28571 16727 28577
rect 16758 28568 16764 28580
rect 16816 28568 16822 28620
rect 18046 28568 18052 28620
rect 18104 28608 18110 28620
rect 18104 28580 18828 28608
rect 18104 28568 18110 28580
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 12621 28543 12679 28549
rect 12621 28509 12633 28543
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 13081 28543 13139 28549
rect 13081 28509 13093 28543
rect 13127 28509 13139 28543
rect 13081 28503 13139 28509
rect 13357 28543 13415 28549
rect 13357 28509 13369 28543
rect 13403 28540 13415 28543
rect 13814 28540 13820 28552
rect 13403 28512 13820 28540
rect 13403 28509 13415 28512
rect 13357 28503 13415 28509
rect 10321 28475 10379 28481
rect 10321 28441 10333 28475
rect 10367 28472 10379 28475
rect 10686 28472 10692 28484
rect 10367 28444 10692 28472
rect 10367 28441 10379 28444
rect 10321 28435 10379 28441
rect 10686 28432 10692 28444
rect 10744 28432 10750 28484
rect 11638 28444 11744 28472
rect 5184 28376 6040 28404
rect 9582 28364 9588 28416
rect 9640 28404 9646 28416
rect 9953 28407 10011 28413
rect 9953 28404 9965 28407
rect 9640 28376 9965 28404
rect 9640 28364 9646 28376
rect 9953 28373 9965 28376
rect 9999 28373 10011 28407
rect 11716 28404 11744 28444
rect 12066 28432 12072 28484
rect 12124 28432 12130 28484
rect 12529 28407 12587 28413
rect 12529 28404 12541 28407
rect 11716 28376 12541 28404
rect 9953 28367 10011 28373
rect 12529 28373 12541 28376
rect 12575 28373 12587 28407
rect 13004 28404 13032 28503
rect 13814 28500 13820 28512
rect 13872 28540 13878 28552
rect 14182 28540 14188 28552
rect 13872 28512 14188 28540
rect 13872 28500 13878 28512
rect 14182 28500 14188 28512
rect 14240 28500 14246 28552
rect 14274 28500 14280 28552
rect 14332 28500 14338 28552
rect 16298 28500 16304 28552
rect 16356 28540 16362 28552
rect 17034 28540 17040 28552
rect 16356 28512 17040 28540
rect 16356 28500 16362 28512
rect 17034 28500 17040 28512
rect 17092 28540 17098 28552
rect 17402 28540 17408 28552
rect 17092 28512 17408 28540
rect 17092 28500 17098 28512
rect 17402 28500 17408 28512
rect 17460 28500 17466 28552
rect 17954 28500 17960 28552
rect 18012 28540 18018 28552
rect 18800 28549 18828 28580
rect 19260 28549 19288 28716
rect 19337 28713 19349 28747
rect 19383 28744 19395 28747
rect 19518 28744 19524 28756
rect 19383 28716 19524 28744
rect 19383 28713 19395 28716
rect 19337 28707 19395 28713
rect 19518 28704 19524 28716
rect 19576 28704 19582 28756
rect 18417 28543 18475 28549
rect 18417 28540 18429 28543
rect 18012 28512 18429 28540
rect 18012 28500 18018 28512
rect 18417 28509 18429 28512
rect 18463 28509 18475 28543
rect 18417 28503 18475 28509
rect 18785 28543 18843 28549
rect 18785 28509 18797 28543
rect 18831 28509 18843 28543
rect 18785 28503 18843 28509
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28540 19303 28543
rect 19291 28512 19380 28540
rect 19291 28509 19303 28512
rect 19245 28503 19303 28509
rect 13170 28432 13176 28484
rect 13228 28432 13234 28484
rect 13998 28404 14004 28416
rect 13004 28376 14004 28404
rect 12529 28367 12587 28373
rect 13998 28364 14004 28376
rect 14056 28364 14062 28416
rect 18432 28404 18460 28503
rect 18506 28432 18512 28484
rect 18564 28432 18570 28484
rect 18598 28432 18604 28484
rect 18656 28432 18662 28484
rect 18800 28472 18828 28503
rect 19352 28472 19380 28512
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20349 28543 20407 28549
rect 20349 28540 20361 28543
rect 20036 28512 20361 28540
rect 20036 28500 20042 28512
rect 20349 28509 20361 28512
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20605 28543 20663 28549
rect 20605 28540 20617 28543
rect 20496 28512 20617 28540
rect 20496 28500 20502 28512
rect 20605 28509 20617 28512
rect 20651 28509 20663 28543
rect 20605 28503 20663 28509
rect 21082 28472 21088 28484
rect 18800 28444 19288 28472
rect 19352 28444 21088 28472
rect 19260 28416 19288 28444
rect 21082 28432 21088 28444
rect 21140 28432 21146 28484
rect 19150 28404 19156 28416
rect 18432 28376 19156 28404
rect 19150 28364 19156 28376
rect 19208 28364 19214 28416
rect 19242 28364 19248 28416
rect 19300 28364 19306 28416
rect 20990 28364 20996 28416
rect 21048 28404 21054 28416
rect 21729 28407 21787 28413
rect 21729 28404 21741 28407
rect 21048 28376 21741 28404
rect 21048 28364 21054 28376
rect 21729 28373 21741 28376
rect 21775 28373 21787 28407
rect 21729 28367 21787 28373
rect 1104 28314 38824 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 38824 28314
rect 1104 28240 38824 28262
rect 5810 28160 5816 28212
rect 5868 28200 5874 28212
rect 6454 28200 6460 28212
rect 5868 28172 6460 28200
rect 5868 28160 5874 28172
rect 6454 28160 6460 28172
rect 6512 28160 6518 28212
rect 6638 28160 6644 28212
rect 6696 28160 6702 28212
rect 6733 28203 6791 28209
rect 6733 28169 6745 28203
rect 6779 28200 6791 28203
rect 7009 28203 7067 28209
rect 7009 28200 7021 28203
rect 6779 28172 7021 28200
rect 6779 28169 6791 28172
rect 6733 28163 6791 28169
rect 7009 28169 7021 28172
rect 7055 28169 7067 28203
rect 7009 28163 7067 28169
rect 7282 28160 7288 28212
rect 7340 28160 7346 28212
rect 9401 28203 9459 28209
rect 9401 28200 9413 28203
rect 8588 28172 9413 28200
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28064 6423 28067
rect 6472 28064 6500 28160
rect 6411 28036 6500 28064
rect 6411 28033 6423 28036
rect 6365 28027 6423 28033
rect 6457 27999 6515 28005
rect 6457 27965 6469 27999
rect 6503 27965 6515 27999
rect 6457 27959 6515 27965
rect 5534 27820 5540 27872
rect 5592 27860 5598 27872
rect 6365 27863 6423 27869
rect 6365 27860 6377 27863
rect 5592 27832 6377 27860
rect 5592 27820 5598 27832
rect 6365 27829 6377 27832
rect 6411 27829 6423 27863
rect 6472 27860 6500 27959
rect 6656 27928 6684 28160
rect 6825 28135 6883 28141
rect 6825 28101 6837 28135
rect 6871 28132 6883 28135
rect 6914 28132 6920 28144
rect 6871 28104 6920 28132
rect 6871 28101 6883 28104
rect 6825 28095 6883 28101
rect 6914 28092 6920 28104
rect 6972 28092 6978 28144
rect 7101 28067 7159 28073
rect 7101 28033 7113 28067
rect 7147 28064 7159 28067
rect 7300 28064 7328 28160
rect 8588 28073 8616 28172
rect 9401 28169 9413 28172
rect 9447 28200 9459 28203
rect 10778 28200 10784 28212
rect 9447 28172 10784 28200
rect 9447 28169 9459 28172
rect 9401 28163 9459 28169
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 12066 28160 12072 28212
rect 12124 28200 12130 28212
rect 12897 28203 12955 28209
rect 12897 28200 12909 28203
rect 12124 28172 12909 28200
rect 12124 28160 12130 28172
rect 12897 28169 12909 28172
rect 12943 28169 12955 28203
rect 13722 28200 13728 28212
rect 12897 28163 12955 28169
rect 13188 28172 13728 28200
rect 9582 28132 9588 28144
rect 9232 28104 9588 28132
rect 9232 28076 9260 28104
rect 9582 28092 9588 28104
rect 9640 28132 9646 28144
rect 13188 28141 13216 28172
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 13817 28203 13875 28209
rect 13817 28169 13829 28203
rect 13863 28169 13875 28203
rect 13817 28163 13875 28169
rect 13173 28135 13231 28141
rect 9640 28104 9996 28132
rect 9640 28092 9646 28104
rect 7147 28036 7328 28064
rect 8389 28067 8447 28073
rect 7147 28033 7159 28036
rect 7101 28027 7159 28033
rect 8389 28033 8401 28067
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28033 8631 28067
rect 8573 28027 8631 28033
rect 8404 27996 8432 28027
rect 9214 28024 9220 28076
rect 9272 28024 9278 28076
rect 9398 28024 9404 28076
rect 9456 28024 9462 28076
rect 9968 28073 9996 28104
rect 13173 28101 13185 28135
rect 13219 28101 13231 28135
rect 13173 28095 13231 28101
rect 13265 28135 13323 28141
rect 13265 28101 13277 28135
rect 13311 28132 13323 28135
rect 13832 28132 13860 28163
rect 13998 28160 14004 28212
rect 14056 28200 14062 28212
rect 15194 28200 15200 28212
rect 14056 28172 15200 28200
rect 14056 28160 14062 28172
rect 15194 28160 15200 28172
rect 15252 28160 15258 28212
rect 15764 28172 16528 28200
rect 13311 28104 13860 28132
rect 13311 28101 13323 28104
rect 13265 28095 13323 28101
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 10226 28024 10232 28076
rect 10284 28024 10290 28076
rect 13078 28024 13084 28076
rect 13136 28024 13142 28076
rect 13354 28024 13360 28076
rect 13412 28064 13418 28076
rect 14016 28073 14044 28160
rect 14108 28104 15056 28132
rect 13449 28067 13507 28073
rect 13449 28064 13461 28067
rect 13412 28036 13461 28064
rect 13412 28024 13418 28036
rect 13449 28033 13461 28036
rect 13495 28033 13507 28067
rect 13449 28027 13507 28033
rect 14001 28067 14059 28073
rect 14001 28033 14013 28067
rect 14047 28033 14059 28067
rect 14001 28027 14059 28033
rect 9674 27996 9680 28008
rect 8404 27968 9680 27996
rect 9674 27956 9680 27968
rect 9732 27956 9738 28008
rect 9766 27956 9772 28008
rect 9824 27956 9830 28008
rect 13262 27956 13268 28008
rect 13320 27996 13326 28008
rect 14108 27996 14136 28104
rect 14185 28067 14243 28073
rect 14185 28033 14197 28067
rect 14231 28064 14243 28067
rect 14231 28036 14596 28064
rect 14231 28033 14243 28036
rect 14185 28027 14243 28033
rect 13320 27968 14136 27996
rect 13320 27956 13326 27968
rect 6825 27931 6883 27937
rect 6825 27928 6837 27931
rect 6656 27900 6837 27928
rect 6825 27897 6837 27900
rect 6871 27897 6883 27931
rect 6825 27891 6883 27897
rect 7466 27860 7472 27872
rect 6472 27832 7472 27860
rect 6365 27823 6423 27829
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 8478 27820 8484 27872
rect 8536 27820 8542 27872
rect 10134 27820 10140 27872
rect 10192 27820 10198 27872
rect 10410 27820 10416 27872
rect 10468 27820 10474 27872
rect 14185 27863 14243 27869
rect 14185 27829 14197 27863
rect 14231 27860 14243 27863
rect 14366 27860 14372 27872
rect 14231 27832 14372 27860
rect 14231 27829 14243 27832
rect 14185 27823 14243 27829
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 14568 27869 14596 28036
rect 15028 28005 15056 28104
rect 15764 28076 15792 28172
rect 16500 28144 16528 28172
rect 18598 28160 18604 28212
rect 18656 28200 18662 28212
rect 18877 28203 18935 28209
rect 18877 28200 18889 28203
rect 18656 28172 18889 28200
rect 18656 28160 18662 28172
rect 18877 28169 18889 28172
rect 18923 28169 18935 28203
rect 18877 28163 18935 28169
rect 19150 28160 19156 28212
rect 19208 28160 19214 28212
rect 19242 28160 19248 28212
rect 19300 28200 19306 28212
rect 19797 28203 19855 28209
rect 19797 28200 19809 28203
rect 19300 28172 19809 28200
rect 19300 28160 19306 28172
rect 19797 28169 19809 28172
rect 19843 28200 19855 28203
rect 20533 28203 20591 28209
rect 20533 28200 20545 28203
rect 19843 28172 20545 28200
rect 19843 28169 19855 28172
rect 19797 28163 19855 28169
rect 20533 28169 20545 28172
rect 20579 28169 20591 28203
rect 20533 28163 20591 28169
rect 16285 28135 16343 28141
rect 16285 28132 16297 28135
rect 16040 28104 16297 28132
rect 15746 28024 15752 28076
rect 15804 28024 15810 28076
rect 16040 28073 16068 28104
rect 16285 28101 16297 28104
rect 16331 28132 16343 28135
rect 16390 28132 16396 28144
rect 16331 28104 16396 28132
rect 16331 28101 16343 28104
rect 16285 28095 16343 28101
rect 16390 28092 16396 28104
rect 16448 28092 16454 28144
rect 16482 28092 16488 28144
rect 16540 28092 16546 28144
rect 18506 28092 18512 28144
rect 18564 28132 18570 28144
rect 20990 28132 20996 28144
rect 18564 28104 19196 28132
rect 18564 28092 18570 28104
rect 19168 28076 19196 28104
rect 20732 28104 20996 28132
rect 15933 28067 15991 28073
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16025 28067 16083 28073
rect 16025 28033 16037 28067
rect 16071 28033 16083 28067
rect 16025 28027 16083 28033
rect 15013 27999 15071 28005
rect 15013 27965 15025 27999
rect 15059 27965 15071 27999
rect 15948 27996 15976 28027
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 18690 28024 18696 28076
rect 18748 28024 18754 28076
rect 19150 28024 19156 28076
rect 19208 28024 19214 28076
rect 20732 28073 20760 28104
rect 20990 28092 20996 28104
rect 21048 28092 21054 28144
rect 22002 28092 22008 28144
rect 22060 28132 22066 28144
rect 22370 28132 22376 28144
rect 22060 28104 22376 28132
rect 22060 28092 22066 28104
rect 22370 28092 22376 28104
rect 22428 28092 22434 28144
rect 22646 28132 22652 28144
rect 22480 28104 22652 28132
rect 20717 28067 20775 28073
rect 20717 28033 20729 28067
rect 20763 28033 20775 28067
rect 20717 28027 20775 28033
rect 20898 28024 20904 28076
rect 20956 28064 20962 28076
rect 22480 28064 22508 28104
rect 22646 28092 22652 28104
rect 22704 28132 22710 28144
rect 23017 28135 23075 28141
rect 23017 28132 23029 28135
rect 22704 28104 23029 28132
rect 22704 28092 22710 28104
rect 23017 28101 23029 28104
rect 23063 28101 23075 28135
rect 23017 28095 23075 28101
rect 20956 28036 22508 28064
rect 22557 28067 22615 28073
rect 20956 28024 20962 28036
rect 22557 28033 22569 28067
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 15948 27968 16344 27996
rect 15013 27959 15071 27965
rect 14734 27888 14740 27940
rect 14792 27888 14798 27940
rect 15028 27928 15056 27959
rect 16117 27931 16175 27937
rect 16117 27928 16129 27931
rect 15028 27900 16129 27928
rect 16117 27897 16129 27900
rect 16163 27897 16175 27931
rect 16117 27891 16175 27897
rect 16316 27872 16344 27968
rect 19334 27956 19340 28008
rect 19392 27956 19398 28008
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27996 19487 27999
rect 20993 27999 21051 28005
rect 19475 27968 19748 27996
rect 19475 27965 19487 27968
rect 19429 27959 19487 27965
rect 19720 27928 19748 27968
rect 20993 27965 21005 27999
rect 21039 27965 21051 27999
rect 20993 27959 21051 27965
rect 21008 27928 21036 27959
rect 22002 27956 22008 28008
rect 22060 27956 22066 28008
rect 22572 27996 22600 28027
rect 22830 28024 22836 28076
rect 22888 28024 22894 28076
rect 23201 27999 23259 28005
rect 23201 27996 23213 27999
rect 22572 27968 23213 27996
rect 23201 27965 23213 27968
rect 23247 27965 23259 27999
rect 23201 27959 23259 27965
rect 19720 27900 21036 27928
rect 19720 27872 19748 27900
rect 22186 27888 22192 27940
rect 22244 27928 22250 27940
rect 22281 27931 22339 27937
rect 22281 27928 22293 27931
rect 22244 27900 22293 27928
rect 22244 27888 22250 27900
rect 22281 27897 22293 27900
rect 22327 27897 22339 27931
rect 22281 27891 22339 27897
rect 22741 27931 22799 27937
rect 22741 27897 22753 27931
rect 22787 27928 22799 27931
rect 23474 27928 23480 27940
rect 22787 27900 23480 27928
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 23474 27888 23480 27900
rect 23532 27888 23538 27940
rect 14553 27863 14611 27869
rect 14553 27829 14565 27863
rect 14599 27860 14611 27863
rect 14642 27860 14648 27872
rect 14599 27832 14648 27860
rect 14599 27829 14611 27832
rect 14553 27823 14611 27829
rect 14642 27820 14648 27832
rect 14700 27820 14706 27872
rect 15378 27820 15384 27872
rect 15436 27860 15442 27872
rect 15565 27863 15623 27869
rect 15565 27860 15577 27863
rect 15436 27832 15577 27860
rect 15436 27820 15442 27832
rect 15565 27829 15577 27832
rect 15611 27829 15623 27863
rect 15565 27823 15623 27829
rect 16298 27820 16304 27872
rect 16356 27820 16362 27872
rect 19702 27820 19708 27872
rect 19760 27820 19766 27872
rect 22462 27820 22468 27872
rect 22520 27820 22526 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 4062 27616 4068 27668
rect 4120 27656 4126 27668
rect 5534 27656 5540 27668
rect 4120 27628 5540 27656
rect 4120 27616 4126 27628
rect 5534 27616 5540 27628
rect 5592 27616 5598 27668
rect 6365 27659 6423 27665
rect 6365 27625 6377 27659
rect 6411 27656 6423 27659
rect 6454 27656 6460 27668
rect 6411 27628 6460 27656
rect 6411 27625 6423 27628
rect 6365 27619 6423 27625
rect 6454 27616 6460 27628
rect 6512 27616 6518 27668
rect 8941 27659 8999 27665
rect 8941 27625 8953 27659
rect 8987 27656 8999 27659
rect 9398 27656 9404 27668
rect 8987 27628 9404 27656
rect 8987 27625 8999 27628
rect 8941 27619 8999 27625
rect 9398 27616 9404 27628
rect 9456 27616 9462 27668
rect 12713 27659 12771 27665
rect 12713 27625 12725 27659
rect 12759 27656 12771 27659
rect 12897 27659 12955 27665
rect 12759 27628 12848 27656
rect 12759 27625 12771 27628
rect 12713 27619 12771 27625
rect 5169 27591 5227 27597
rect 5169 27557 5181 27591
rect 5215 27557 5227 27591
rect 5169 27551 5227 27557
rect 12253 27591 12311 27597
rect 12253 27557 12265 27591
rect 12299 27557 12311 27591
rect 12820 27588 12848 27628
rect 12897 27625 12909 27659
rect 12943 27656 12955 27659
rect 13170 27656 13176 27668
rect 12943 27628 13176 27656
rect 12943 27625 12955 27628
rect 12897 27619 12955 27625
rect 13170 27616 13176 27628
rect 13228 27616 13234 27668
rect 13280 27628 14136 27656
rect 13280 27588 13308 27628
rect 14108 27597 14136 27628
rect 14734 27616 14740 27668
rect 14792 27656 14798 27668
rect 14792 27628 15240 27656
rect 14792 27616 14798 27628
rect 12820 27560 13308 27588
rect 14093 27591 14151 27597
rect 12253 27551 12311 27557
rect 14093 27557 14105 27591
rect 14139 27557 14151 27591
rect 14093 27551 14151 27557
rect 15013 27591 15071 27597
rect 15013 27557 15025 27591
rect 15059 27588 15071 27591
rect 15102 27588 15108 27600
rect 15059 27560 15108 27588
rect 15059 27557 15071 27560
rect 15013 27551 15071 27557
rect 5184 27520 5212 27551
rect 5813 27523 5871 27529
rect 5813 27520 5825 27523
rect 5184 27492 5825 27520
rect 5813 27489 5825 27492
rect 5859 27489 5871 27523
rect 8478 27520 8484 27532
rect 5813 27483 5871 27489
rect 7576 27492 8484 27520
rect 3786 27412 3792 27464
rect 3844 27412 3850 27464
rect 5828 27452 5856 27483
rect 7576 27461 7604 27492
rect 8478 27480 8484 27492
rect 8536 27480 8542 27532
rect 5997 27455 6055 27461
rect 5997 27452 6009 27455
rect 5828 27424 6009 27452
rect 5997 27421 6009 27424
rect 6043 27421 6055 27455
rect 5997 27415 6055 27421
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27421 7435 27455
rect 7377 27415 7435 27421
rect 7561 27455 7619 27461
rect 7561 27421 7573 27455
rect 7607 27421 7619 27455
rect 7561 27415 7619 27421
rect 4056 27387 4114 27393
rect 4056 27353 4068 27387
rect 4102 27384 4114 27387
rect 4154 27384 4160 27396
rect 4102 27356 4160 27384
rect 4102 27353 4114 27356
rect 4056 27347 4114 27353
rect 4154 27344 4160 27356
rect 4212 27344 4218 27396
rect 6181 27387 6239 27393
rect 6181 27384 6193 27387
rect 6104 27356 6193 27384
rect 6104 27328 6132 27356
rect 6181 27353 6193 27356
rect 6227 27353 6239 27387
rect 7392 27384 7420 27415
rect 8386 27412 8392 27464
rect 8444 27412 8450 27464
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27452 9643 27455
rect 9766 27452 9772 27464
rect 9631 27424 9772 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 7745 27387 7803 27393
rect 7745 27384 7757 27387
rect 7392 27356 7757 27384
rect 6181 27347 6239 27353
rect 7745 27353 7757 27356
rect 7791 27353 7803 27387
rect 7745 27347 7803 27353
rect 5258 27276 5264 27328
rect 5316 27276 5322 27328
rect 6086 27276 6092 27328
rect 6144 27276 6150 27328
rect 7374 27276 7380 27328
rect 7432 27276 7438 27328
rect 9692 27325 9720 27424
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 10410 27412 10416 27464
rect 10468 27452 10474 27464
rect 10790 27455 10848 27461
rect 10790 27452 10802 27455
rect 10468 27424 10802 27452
rect 10468 27412 10474 27424
rect 10790 27421 10802 27424
rect 10836 27421 10848 27455
rect 10790 27415 10848 27421
rect 11054 27412 11060 27464
rect 11112 27412 11118 27464
rect 11974 27412 11980 27464
rect 12032 27412 12038 27464
rect 12268 27452 12296 27551
rect 15102 27548 15108 27560
rect 15160 27548 15166 27600
rect 15212 27588 15240 27628
rect 17052 27628 17356 27656
rect 17052 27588 17080 27628
rect 15212 27560 17080 27588
rect 13262 27480 13268 27532
rect 13320 27480 13326 27532
rect 13630 27480 13636 27532
rect 13688 27520 13694 27532
rect 14461 27523 14519 27529
rect 13688 27492 14044 27520
rect 13688 27480 13694 27492
rect 12345 27455 12403 27461
rect 12345 27452 12357 27455
rect 12268 27424 12357 27452
rect 12345 27421 12357 27424
rect 12391 27421 12403 27455
rect 12345 27415 12403 27421
rect 12618 27412 12624 27464
rect 12676 27412 12682 27464
rect 13909 27455 13967 27461
rect 13909 27452 13921 27455
rect 13740 27424 13921 27452
rect 12253 27387 12311 27393
rect 12253 27353 12265 27387
rect 12299 27384 12311 27387
rect 13148 27387 13206 27393
rect 12299 27356 13032 27384
rect 12299 27353 12311 27356
rect 12253 27347 12311 27353
rect 9677 27319 9735 27325
rect 9677 27285 9689 27319
rect 9723 27316 9735 27319
rect 10318 27316 10324 27328
rect 9723 27288 10324 27316
rect 9723 27285 9735 27288
rect 9677 27279 9735 27285
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 12069 27319 12127 27325
rect 12069 27285 12081 27319
rect 12115 27316 12127 27319
rect 12434 27316 12440 27328
rect 12115 27288 12440 27316
rect 12115 27285 12127 27288
rect 12069 27279 12127 27285
rect 12434 27276 12440 27288
rect 12492 27276 12498 27328
rect 13004 27325 13032 27356
rect 13148 27353 13160 27387
rect 13194 27384 13206 27387
rect 13538 27384 13544 27396
rect 13194 27356 13544 27384
rect 13194 27353 13206 27356
rect 13148 27347 13206 27353
rect 13538 27344 13544 27356
rect 13596 27344 13602 27396
rect 12989 27319 13047 27325
rect 12989 27285 13001 27319
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 13740 27316 13768 27424
rect 13909 27421 13921 27424
rect 13955 27421 13967 27455
rect 13909 27415 13967 27421
rect 14016 27384 14044 27492
rect 14461 27489 14473 27523
rect 14507 27520 14519 27523
rect 14642 27520 14648 27532
rect 14507 27492 14648 27520
rect 14507 27489 14519 27492
rect 14461 27483 14519 27489
rect 14642 27480 14648 27492
rect 14700 27520 14706 27532
rect 14700 27492 15516 27520
rect 14700 27480 14706 27492
rect 14274 27412 14280 27464
rect 14332 27412 14338 27464
rect 14366 27412 14372 27464
rect 14424 27412 14430 27464
rect 14550 27412 14556 27464
rect 14608 27412 14614 27464
rect 15010 27412 15016 27464
rect 15068 27452 15074 27464
rect 15151 27455 15209 27461
rect 15151 27452 15163 27455
rect 15068 27424 15163 27452
rect 15068 27412 15074 27424
rect 15151 27421 15163 27424
rect 15197 27452 15209 27455
rect 15197 27421 15235 27452
rect 15151 27415 15235 27421
rect 14568 27384 14596 27412
rect 14016 27356 14596 27384
rect 13412 27288 13768 27316
rect 13412 27276 13418 27288
rect 13814 27276 13820 27328
rect 13872 27276 13878 27328
rect 15207 27316 15235 27415
rect 15286 27412 15292 27464
rect 15344 27412 15350 27464
rect 15378 27412 15384 27464
rect 15436 27412 15442 27464
rect 15488 27461 15516 27492
rect 15488 27455 15567 27461
rect 15488 27424 15521 27455
rect 15509 27421 15521 27424
rect 15555 27421 15567 27455
rect 15509 27415 15567 27421
rect 15654 27412 15660 27464
rect 15712 27412 15718 27464
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 16684 27461 16712 27560
rect 17126 27548 17132 27600
rect 17184 27588 17190 27600
rect 17221 27591 17279 27597
rect 17221 27588 17233 27591
rect 17184 27560 17233 27588
rect 17184 27548 17190 27560
rect 17221 27557 17233 27560
rect 17267 27557 17279 27591
rect 17328 27588 17356 27628
rect 18690 27616 18696 27668
rect 18748 27616 18754 27668
rect 20898 27656 20904 27668
rect 20364 27628 20904 27656
rect 20364 27588 20392 27628
rect 20898 27616 20904 27628
rect 20956 27616 20962 27668
rect 22557 27659 22615 27665
rect 22557 27625 22569 27659
rect 22603 27656 22615 27659
rect 22830 27656 22836 27668
rect 22603 27628 22836 27656
rect 22603 27625 22615 27628
rect 22557 27619 22615 27625
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 17328 27560 20392 27588
rect 17221 27551 17279 27557
rect 16942 27480 16948 27532
rect 17000 27520 17006 27532
rect 19245 27523 19303 27529
rect 19245 27520 19257 27523
rect 17000 27492 19257 27520
rect 17000 27480 17006 27492
rect 16670 27455 16728 27461
rect 16670 27421 16682 27455
rect 16716 27421 16728 27455
rect 16670 27415 16728 27421
rect 16758 27412 16764 27464
rect 16816 27412 16822 27464
rect 17042 27455 17100 27461
rect 17042 27421 17054 27455
rect 17088 27452 17100 27455
rect 18141 27455 18199 27461
rect 17088 27424 17264 27452
rect 17088 27421 17100 27424
rect 17042 27415 17100 27421
rect 16776 27384 16804 27412
rect 16853 27387 16911 27393
rect 16853 27384 16865 27387
rect 16776 27356 16865 27384
rect 16853 27353 16865 27356
rect 16899 27353 16911 27387
rect 16853 27347 16911 27353
rect 16965 27387 17023 27393
rect 16965 27353 16977 27387
rect 17011 27384 17023 27387
rect 17126 27384 17132 27396
rect 17011 27356 17132 27384
rect 17011 27353 17023 27356
rect 16965 27347 17023 27353
rect 17126 27344 17132 27356
rect 17184 27344 17190 27396
rect 17236 27384 17264 27424
rect 18141 27421 18153 27455
rect 18187 27452 18199 27455
rect 18230 27452 18236 27464
rect 18187 27424 18236 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 18524 27461 18552 27492
rect 19245 27489 19257 27492
rect 19291 27489 19303 27523
rect 19536 27520 19564 27560
rect 22554 27520 22560 27532
rect 19245 27483 19303 27489
rect 19444 27492 19564 27520
rect 19628 27492 22560 27520
rect 19444 27461 19472 27492
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 18969 27455 19027 27461
rect 18969 27421 18981 27455
rect 19015 27421 19027 27455
rect 18969 27415 19027 27421
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 18046 27384 18052 27396
rect 17236 27356 18052 27384
rect 17236 27316 17264 27356
rect 18046 27344 18052 27356
rect 18104 27344 18110 27396
rect 18322 27344 18328 27396
rect 18380 27344 18386 27396
rect 18417 27387 18475 27393
rect 18417 27353 18429 27387
rect 18463 27384 18475 27387
rect 18877 27387 18935 27393
rect 18877 27384 18889 27387
rect 18463 27356 18889 27384
rect 18463 27353 18475 27356
rect 18417 27347 18475 27353
rect 18877 27353 18889 27356
rect 18923 27353 18935 27387
rect 18877 27347 18935 27353
rect 15207 27288 17264 27316
rect 18984 27316 19012 27415
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 19628 27461 19656 27492
rect 22554 27480 22560 27492
rect 22612 27480 22618 27532
rect 19613 27455 19671 27461
rect 19613 27452 19625 27455
rect 19576 27424 19625 27452
rect 19576 27412 19582 27424
rect 19613 27421 19625 27424
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27452 19763 27455
rect 19751 27424 19840 27452
rect 19751 27421 19763 27424
rect 19705 27415 19763 27421
rect 19058 27344 19064 27396
rect 19116 27384 19122 27396
rect 19536 27384 19564 27412
rect 19116 27356 19564 27384
rect 19116 27344 19122 27356
rect 19812 27328 19840 27424
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20257 27455 20315 27461
rect 20257 27452 20269 27455
rect 20036 27424 20269 27452
rect 20036 27412 20042 27424
rect 20257 27421 20269 27424
rect 20303 27421 20315 27455
rect 20257 27415 20315 27421
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 22373 27455 22431 27461
rect 22373 27421 22385 27455
rect 22419 27452 22431 27455
rect 22419 27424 22876 27452
rect 22419 27421 22431 27424
rect 22373 27415 22431 27421
rect 20530 27344 20536 27396
rect 20588 27344 20594 27396
rect 21266 27344 21272 27396
rect 21324 27344 21330 27396
rect 22296 27384 22324 27415
rect 22296 27356 22692 27384
rect 19150 27316 19156 27328
rect 18984 27288 19156 27316
rect 19150 27276 19156 27288
rect 19208 27276 19214 27328
rect 19794 27276 19800 27328
rect 19852 27276 19858 27328
rect 22002 27276 22008 27328
rect 22060 27276 22066 27328
rect 22664 27325 22692 27356
rect 22848 27328 22876 27424
rect 23474 27412 23480 27464
rect 23532 27452 23538 27464
rect 23762 27455 23820 27461
rect 23762 27452 23774 27455
rect 23532 27424 23774 27452
rect 23532 27412 23538 27424
rect 23762 27421 23774 27424
rect 23808 27421 23820 27455
rect 23762 27415 23820 27421
rect 23934 27412 23940 27464
rect 23992 27452 23998 27464
rect 24029 27455 24087 27461
rect 24029 27452 24041 27455
rect 23992 27424 24041 27452
rect 23992 27412 23998 27424
rect 24029 27421 24041 27424
rect 24075 27421 24087 27455
rect 24029 27415 24087 27421
rect 22649 27319 22707 27325
rect 22649 27285 22661 27319
rect 22695 27316 22707 27319
rect 22738 27316 22744 27328
rect 22695 27288 22744 27316
rect 22695 27285 22707 27288
rect 22649 27279 22707 27285
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 22830 27276 22836 27328
rect 22888 27276 22894 27328
rect 1104 27226 38824 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 38824 27226
rect 1104 27152 38824 27174
rect 4154 27072 4160 27124
rect 4212 27072 4218 27124
rect 5258 27072 5264 27124
rect 5316 27072 5322 27124
rect 5534 27072 5540 27124
rect 5592 27072 5598 27124
rect 7374 27072 7380 27124
rect 7432 27072 7438 27124
rect 10226 27072 10232 27124
rect 10284 27112 10290 27124
rect 10965 27115 11023 27121
rect 10965 27112 10977 27115
rect 10284 27084 10977 27112
rect 10284 27072 10290 27084
rect 10965 27081 10977 27084
rect 11011 27081 11023 27115
rect 10965 27075 11023 27081
rect 12529 27115 12587 27121
rect 12529 27081 12541 27115
rect 12575 27112 12587 27115
rect 12618 27112 12624 27124
rect 12575 27084 12624 27112
rect 12575 27081 12587 27084
rect 12529 27075 12587 27081
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 13078 27072 13084 27124
rect 13136 27112 13142 27124
rect 13449 27115 13507 27121
rect 13449 27112 13461 27115
rect 13136 27084 13461 27112
rect 13136 27072 13142 27084
rect 13449 27081 13461 27084
rect 13495 27081 13507 27115
rect 13449 27075 13507 27081
rect 13538 27072 13544 27124
rect 13596 27112 13602 27124
rect 13722 27112 13728 27124
rect 13596 27084 13728 27112
rect 13596 27072 13602 27084
rect 13722 27072 13728 27084
rect 13780 27072 13786 27124
rect 13814 27072 13820 27124
rect 13872 27072 13878 27124
rect 14093 27115 14151 27121
rect 14093 27081 14105 27115
rect 14139 27112 14151 27115
rect 14274 27112 14280 27124
rect 14139 27084 14280 27112
rect 14139 27081 14151 27084
rect 14093 27075 14151 27081
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 15565 27115 15623 27121
rect 15565 27081 15577 27115
rect 15611 27112 15623 27115
rect 15654 27112 15660 27124
rect 15611 27084 15660 27112
rect 15611 27081 15623 27084
rect 15565 27075 15623 27081
rect 15654 27072 15660 27084
rect 15712 27072 15718 27124
rect 17034 27112 17040 27124
rect 15764 27084 17040 27112
rect 5276 26985 5304 27072
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26945 5319 26979
rect 5552 26976 5580 27072
rect 5721 26979 5779 26985
rect 5721 26976 5733 26979
rect 5552 26948 5733 26976
rect 5261 26939 5319 26945
rect 5721 26945 5733 26948
rect 5767 26976 5779 26979
rect 5997 26979 6055 26985
rect 5997 26976 6009 26979
rect 5767 26948 6009 26976
rect 5767 26945 5779 26948
rect 5721 26939 5779 26945
rect 5997 26945 6009 26948
rect 6043 26945 6055 26979
rect 5997 26939 6055 26945
rect 6086 26936 6092 26988
rect 6144 26976 6150 26988
rect 6181 26979 6239 26985
rect 6181 26976 6193 26979
rect 6144 26948 6193 26976
rect 6144 26936 6150 26948
rect 6181 26945 6193 26948
rect 6227 26976 6239 26979
rect 6917 26979 6975 26985
rect 6917 26976 6929 26979
rect 6227 26948 6929 26976
rect 6227 26945 6239 26948
rect 6181 26939 6239 26945
rect 6917 26945 6929 26948
rect 6963 26945 6975 26979
rect 6917 26939 6975 26945
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26976 7343 26979
rect 7392 26976 7420 27072
rect 11054 27044 11060 27056
rect 8404 27016 11060 27044
rect 7331 26948 7420 26976
rect 7331 26945 7343 26948
rect 7285 26939 7343 26945
rect 3326 26868 3332 26920
rect 3384 26868 3390 26920
rect 4801 26911 4859 26917
rect 4801 26877 4813 26911
rect 4847 26908 4859 26911
rect 4893 26911 4951 26917
rect 4893 26908 4905 26911
rect 4847 26880 4905 26908
rect 4847 26877 4859 26880
rect 4801 26871 4859 26877
rect 4893 26877 4905 26880
rect 4939 26877 4951 26911
rect 4893 26871 4951 26877
rect 5353 26911 5411 26917
rect 5353 26877 5365 26911
rect 5399 26877 5411 26911
rect 5353 26871 5411 26877
rect 5905 26911 5963 26917
rect 5905 26877 5917 26911
rect 5951 26908 5963 26911
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 5951 26880 6377 26908
rect 5951 26877 5963 26880
rect 5905 26871 5963 26877
rect 6365 26877 6377 26880
rect 6411 26877 6423 26911
rect 7116 26908 7144 26939
rect 8202 26936 8208 26988
rect 8260 26936 8266 26988
rect 8404 26985 8432 27016
rect 11054 27004 11060 27016
rect 11112 27004 11118 27056
rect 11992 27016 12848 27044
rect 8389 26979 8447 26985
rect 8389 26945 8401 26979
rect 8435 26945 8447 26979
rect 8389 26939 8447 26945
rect 8656 26979 8714 26985
rect 8656 26945 8668 26979
rect 8702 26976 8714 26979
rect 8702 26948 9904 26976
rect 8702 26945 8714 26948
rect 8656 26939 8714 26945
rect 7834 26908 7840 26920
rect 7116 26880 7840 26908
rect 6365 26871 6423 26877
rect 5368 26840 5396 26871
rect 7834 26868 7840 26880
rect 7892 26868 7898 26920
rect 9876 26908 9904 26948
rect 10134 26936 10140 26988
rect 10192 26976 10198 26988
rect 10597 26979 10655 26985
rect 10597 26976 10609 26979
rect 10192 26948 10609 26976
rect 10192 26936 10198 26948
rect 10597 26945 10609 26948
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 10778 26936 10784 26988
rect 10836 26976 10842 26988
rect 11241 26979 11299 26985
rect 11241 26976 11253 26979
rect 10836 26948 11253 26976
rect 10836 26936 10842 26948
rect 11241 26945 11253 26948
rect 11287 26945 11299 26979
rect 11241 26939 11299 26945
rect 11333 26979 11391 26985
rect 11333 26945 11345 26979
rect 11379 26945 11391 26979
rect 11333 26939 11391 26945
rect 11793 26979 11851 26985
rect 11793 26945 11805 26979
rect 11839 26945 11851 26979
rect 11793 26939 11851 26945
rect 9876 26880 9996 26908
rect 5626 26840 5632 26852
rect 5368 26812 5632 26840
rect 5626 26800 5632 26812
rect 5684 26840 5690 26852
rect 5997 26843 6055 26849
rect 5997 26840 6009 26843
rect 5684 26812 6009 26840
rect 5684 26800 5690 26812
rect 5997 26809 6009 26812
rect 6043 26809 6055 26843
rect 5997 26803 6055 26809
rect 9766 26800 9772 26852
rect 9824 26800 9830 26852
rect 3973 26775 4031 26781
rect 3973 26741 3985 26775
rect 4019 26772 4031 26775
rect 4614 26772 4620 26784
rect 4019 26744 4620 26772
rect 4019 26741 4031 26744
rect 3973 26735 4031 26741
rect 4614 26732 4620 26744
rect 4672 26732 4678 26784
rect 5534 26732 5540 26784
rect 5592 26732 5598 26784
rect 7190 26732 7196 26784
rect 7248 26732 7254 26784
rect 9490 26732 9496 26784
rect 9548 26772 9554 26784
rect 9861 26775 9919 26781
rect 9861 26772 9873 26775
rect 9548 26744 9873 26772
rect 9548 26732 9554 26744
rect 9861 26741 9873 26744
rect 9907 26741 9919 26775
rect 9968 26772 9996 26880
rect 10318 26868 10324 26920
rect 10376 26919 10382 26920
rect 10376 26917 10456 26919
rect 10376 26911 10471 26917
rect 10376 26891 10425 26911
rect 10376 26868 10382 26891
rect 10413 26877 10425 26891
rect 10459 26877 10471 26911
rect 10413 26871 10471 26877
rect 10962 26868 10968 26920
rect 11020 26908 11026 26920
rect 11057 26911 11115 26917
rect 11057 26908 11069 26911
rect 11020 26880 11069 26908
rect 11020 26868 11026 26880
rect 11057 26877 11069 26880
rect 11103 26877 11115 26911
rect 11057 26871 11115 26877
rect 10502 26800 10508 26852
rect 10560 26840 10566 26852
rect 11348 26840 11376 26939
rect 10560 26812 11376 26840
rect 11808 26840 11836 26939
rect 11882 26936 11888 26988
rect 11940 26976 11946 26988
rect 11992 26985 12020 27016
rect 11977 26979 12035 26985
rect 11977 26976 11989 26979
rect 11940 26948 11989 26976
rect 11940 26936 11946 26948
rect 11977 26945 11989 26948
rect 12023 26945 12035 26979
rect 11977 26939 12035 26945
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12526 26976 12532 26988
rect 12391 26948 12532 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 12820 26985 12848 27016
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26945 12863 26979
rect 12805 26939 12863 26945
rect 13262 26936 13268 26988
rect 13320 26936 13326 26988
rect 13633 26979 13691 26985
rect 13633 26945 13645 26979
rect 13679 26976 13691 26979
rect 13740 26976 13768 27072
rect 13832 26985 13860 27072
rect 15289 27047 15347 27053
rect 15289 27044 15301 27047
rect 14384 27016 15301 27044
rect 13679 26948 13768 26976
rect 13817 26979 13875 26985
rect 13679 26945 13691 26948
rect 13633 26939 13691 26945
rect 13817 26945 13829 26979
rect 13863 26976 13875 26979
rect 14277 26979 14335 26985
rect 14277 26976 14289 26979
rect 13863 26948 14289 26976
rect 13863 26945 13875 26948
rect 13817 26939 13875 26945
rect 14277 26945 14289 26948
rect 14323 26945 14335 26979
rect 14277 26939 14335 26945
rect 12069 26911 12127 26917
rect 12069 26877 12081 26911
rect 12115 26908 12127 26911
rect 12621 26911 12679 26917
rect 12621 26908 12633 26911
rect 12115 26880 12633 26908
rect 12115 26877 12127 26880
rect 12069 26871 12127 26877
rect 12621 26877 12633 26880
rect 12667 26877 12679 26911
rect 12621 26871 12679 26877
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26908 13047 26911
rect 13170 26908 13176 26920
rect 13035 26880 13176 26908
rect 13035 26877 13047 26880
rect 12989 26871 13047 26877
rect 12434 26840 12440 26852
rect 11808 26812 12440 26840
rect 10560 26800 10566 26812
rect 12434 26800 12440 26812
rect 12492 26840 12498 26852
rect 13004 26840 13032 26871
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 13280 26908 13308 26936
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13280 26880 13737 26908
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 13906 26868 13912 26920
rect 13964 26868 13970 26920
rect 12492 26812 13032 26840
rect 12492 26800 12498 26812
rect 11149 26775 11207 26781
rect 11149 26772 11161 26775
rect 9968 26744 11161 26772
rect 9861 26735 9919 26741
rect 11149 26741 11161 26744
rect 11195 26741 11207 26775
rect 11149 26735 11207 26741
rect 11977 26775 12035 26781
rect 11977 26741 11989 26775
rect 12023 26772 12035 26775
rect 12161 26775 12219 26781
rect 12161 26772 12173 26775
rect 12023 26744 12173 26772
rect 12023 26741 12035 26744
rect 11977 26735 12035 26741
rect 12161 26741 12173 26744
rect 12207 26741 12219 26775
rect 12161 26735 12219 26741
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 14384 26772 14412 27016
rect 15289 27013 15301 27016
rect 15335 27044 15347 27047
rect 15764 27044 15792 27084
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 17221 27115 17279 27121
rect 17221 27081 17233 27115
rect 17267 27112 17279 27115
rect 17957 27115 18015 27121
rect 17957 27112 17969 27115
rect 17267 27084 17356 27112
rect 17267 27081 17279 27084
rect 17221 27075 17279 27081
rect 17328 27056 17356 27084
rect 17788 27084 17969 27112
rect 15335 27016 15608 27044
rect 15335 27013 15347 27016
rect 15289 27007 15347 27013
rect 15580 26988 15608 27016
rect 15672 27016 15792 27044
rect 15672 26988 15700 27016
rect 16298 27004 16304 27056
rect 16356 27044 16362 27056
rect 16695 27047 16753 27053
rect 16695 27044 16707 27047
rect 16356 27016 16707 27044
rect 16356 27004 16362 27016
rect 16695 27013 16707 27016
rect 16741 27013 16753 27047
rect 16695 27007 16753 27013
rect 16899 27013 16957 27019
rect 14458 26936 14464 26988
rect 14516 26976 14522 26988
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14516 26948 15025 26976
rect 14516 26936 14522 26948
rect 15013 26945 15025 26948
rect 15059 26945 15071 26979
rect 15013 26939 15071 26945
rect 14553 26911 14611 26917
rect 14553 26877 14565 26911
rect 14599 26908 14611 26911
rect 14734 26908 14740 26920
rect 14599 26880 14740 26908
rect 14599 26877 14611 26880
rect 14553 26871 14611 26877
rect 14734 26868 14740 26880
rect 14792 26868 14798 26920
rect 15028 26908 15056 26939
rect 15194 26936 15200 26988
rect 15252 26936 15258 26988
rect 15378 26936 15384 26988
rect 15436 26936 15442 26988
rect 15562 26936 15568 26988
rect 15620 26936 15626 26988
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 15746 26936 15752 26988
rect 15804 26936 15810 26988
rect 16117 26979 16175 26985
rect 16117 26976 16129 26979
rect 16040 26948 16129 26976
rect 15933 26911 15991 26917
rect 15933 26908 15945 26911
rect 15028 26880 15945 26908
rect 15933 26877 15945 26880
rect 15979 26877 15991 26911
rect 15933 26871 15991 26877
rect 14461 26843 14519 26849
rect 14461 26809 14473 26843
rect 14507 26840 14519 26843
rect 16040 26840 16068 26948
rect 16117 26945 16129 26948
rect 16163 26945 16175 26979
rect 16899 26979 16911 27013
rect 16945 26988 16957 27013
rect 17310 27004 17316 27056
rect 17368 27004 17374 27056
rect 17788 27044 17816 27084
rect 17957 27081 17969 27084
rect 18003 27081 18015 27115
rect 17957 27075 18015 27081
rect 18322 27072 18328 27124
rect 18380 27072 18386 27124
rect 18414 27072 18420 27124
rect 18472 27072 18478 27124
rect 19518 27072 19524 27124
rect 19576 27072 19582 27124
rect 20441 27115 20499 27121
rect 20441 27081 20453 27115
rect 20487 27112 20499 27115
rect 20530 27112 20536 27124
rect 20487 27084 20536 27112
rect 20487 27081 20499 27084
rect 20441 27075 20499 27081
rect 20530 27072 20536 27084
rect 20588 27072 20594 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 21361 27115 21419 27121
rect 21361 27112 21373 27115
rect 21324 27084 21373 27112
rect 21324 27072 21330 27084
rect 21361 27081 21373 27084
rect 21407 27081 21419 27115
rect 21361 27075 21419 27081
rect 22462 27072 22468 27124
rect 22520 27072 22526 27124
rect 22646 27072 22652 27124
rect 22704 27072 22710 27124
rect 23201 27115 23259 27121
rect 23201 27081 23213 27115
rect 23247 27112 23259 27115
rect 23934 27112 23940 27124
rect 23247 27084 23940 27112
rect 23247 27081 23259 27084
rect 23201 27075 23259 27081
rect 23934 27072 23940 27084
rect 23992 27072 23998 27124
rect 18690 27044 18696 27056
rect 17788 27016 18696 27044
rect 17788 26988 17816 27016
rect 18690 27004 18696 27016
rect 18748 27004 18754 27056
rect 18782 27004 18788 27056
rect 18840 27004 18846 27056
rect 16945 26979 16948 26988
rect 16899 26973 16948 26979
rect 16900 26948 16948 26973
rect 16117 26939 16175 26945
rect 16942 26936 16948 26948
rect 17000 26976 17006 26988
rect 17129 26980 17187 26985
rect 17052 26979 17187 26980
rect 17052 26976 17141 26979
rect 17000 26952 17141 26976
rect 17000 26948 17080 26952
rect 17000 26936 17006 26948
rect 17129 26945 17141 26952
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 17402 26936 17408 26988
rect 17460 26936 17466 26988
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26945 17555 26979
rect 17497 26939 17555 26945
rect 17512 26908 17540 26939
rect 17678 26936 17684 26988
rect 17736 26936 17742 26988
rect 17770 26936 17776 26988
rect 17828 26936 17834 26988
rect 17868 26979 17926 26985
rect 17868 26945 17880 26979
rect 17914 26976 17926 26979
rect 17914 26948 18000 26976
rect 17914 26945 17926 26948
rect 17868 26939 17926 26945
rect 17423 26880 17540 26908
rect 17972 26908 18000 26948
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18141 26979 18199 26985
rect 18141 26976 18153 26979
rect 18104 26948 18153 26976
rect 18104 26936 18110 26948
rect 18141 26945 18153 26948
rect 18187 26945 18199 26979
rect 18141 26939 18199 26945
rect 18601 26979 18659 26985
rect 18601 26945 18613 26979
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18414 26908 18420 26920
rect 17972 26880 18420 26908
rect 16942 26840 16948 26852
rect 14507 26812 16948 26840
rect 14507 26809 14519 26812
rect 14461 26803 14519 26809
rect 16942 26800 16948 26812
rect 17000 26800 17006 26852
rect 17423 26849 17451 26880
rect 18414 26868 18420 26880
rect 18472 26908 18478 26920
rect 18616 26908 18644 26939
rect 18472 26880 18644 26908
rect 18472 26868 18478 26880
rect 17405 26843 17463 26849
rect 17405 26809 17417 26843
rect 17451 26809 17463 26843
rect 17405 26803 17463 26809
rect 17494 26800 17500 26852
rect 17552 26800 17558 26852
rect 18800 26840 18828 27004
rect 18969 26979 19027 26985
rect 18969 26945 18981 26979
rect 19015 26976 19027 26979
rect 19153 26979 19211 26985
rect 19153 26976 19165 26979
rect 19015 26948 19165 26976
rect 19015 26945 19027 26948
rect 18969 26939 19027 26945
rect 19153 26945 19165 26948
rect 19199 26945 19211 26979
rect 19153 26939 19211 26945
rect 19245 26979 19303 26985
rect 19245 26945 19257 26979
rect 19291 26976 19303 26979
rect 19536 26976 19564 27072
rect 19613 27047 19671 27053
rect 19613 27013 19625 27047
rect 19659 27044 19671 27047
rect 20714 27044 20720 27056
rect 19659 27016 20720 27044
rect 19659 27013 19671 27016
rect 19613 27007 19671 27013
rect 20714 27004 20720 27016
rect 20772 27044 20778 27056
rect 20993 27047 21051 27053
rect 20993 27044 21005 27047
rect 20772 27016 21005 27044
rect 20772 27004 20778 27016
rect 20993 27013 21005 27016
rect 21039 27013 21051 27047
rect 20993 27007 21051 27013
rect 21082 27004 21088 27056
rect 21140 27044 21146 27056
rect 22480 27044 22508 27072
rect 21140 27016 21312 27044
rect 22480 27016 23060 27044
rect 21140 27004 21146 27016
rect 21284 26985 21312 27016
rect 20855 26979 20913 26985
rect 20855 26976 20867 26979
rect 19291 26948 19564 26976
rect 20364 26948 20867 26976
rect 19291 26945 19303 26948
rect 19245 26939 19303 26945
rect 20364 26852 20392 26948
rect 20855 26945 20867 26948
rect 20901 26945 20913 26979
rect 20855 26939 20913 26945
rect 21269 26979 21327 26985
rect 21269 26945 21281 26979
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 20625 26911 20683 26917
rect 20625 26877 20637 26911
rect 20671 26877 20683 26911
rect 20625 26871 20683 26877
rect 20717 26911 20775 26917
rect 20717 26877 20729 26911
rect 20763 26908 20775 26911
rect 20990 26908 20996 26920
rect 20763 26880 20996 26908
rect 20763 26877 20775 26880
rect 20717 26871 20775 26877
rect 19429 26843 19487 26849
rect 19429 26840 19441 26843
rect 18800 26812 19441 26840
rect 19429 26809 19441 26812
rect 19475 26840 19487 26843
rect 19794 26840 19800 26852
rect 19475 26812 19800 26840
rect 19475 26809 19487 26812
rect 19429 26803 19487 26809
rect 19794 26800 19800 26812
rect 19852 26800 19858 26852
rect 19981 26843 20039 26849
rect 19981 26809 19993 26843
rect 20027 26840 20039 26843
rect 20346 26840 20352 26852
rect 20027 26812 20352 26840
rect 20027 26809 20039 26812
rect 19981 26803 20039 26809
rect 20346 26800 20352 26812
rect 20404 26800 20410 26852
rect 20640 26840 20668 26871
rect 20990 26868 20996 26880
rect 21048 26868 21054 26920
rect 21085 26911 21143 26917
rect 21085 26877 21097 26911
rect 21131 26908 21143 26911
rect 21174 26908 21180 26920
rect 21131 26880 21180 26908
rect 21131 26877 21143 26880
rect 21085 26871 21143 26877
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 21284 26908 21312 26939
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 22373 26979 22431 26985
rect 22373 26976 22385 26979
rect 22060 26948 22385 26976
rect 22060 26936 22066 26948
rect 22373 26945 22385 26948
rect 22419 26945 22431 26979
rect 22373 26939 22431 26945
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26945 22707 26979
rect 22649 26939 22707 26945
rect 21726 26908 21732 26920
rect 21284 26880 21732 26908
rect 21726 26868 21732 26880
rect 21784 26868 21790 26920
rect 22664 26908 22692 26939
rect 22830 26936 22836 26988
rect 22888 26936 22894 26988
rect 23032 26985 23060 27016
rect 23017 26979 23075 26985
rect 23017 26945 23029 26979
rect 23063 26945 23075 26979
rect 23017 26939 23075 26945
rect 22664 26880 22784 26908
rect 21821 26843 21879 26849
rect 21821 26840 21833 26843
rect 20640 26812 21833 26840
rect 21821 26809 21833 26812
rect 21867 26809 21879 26843
rect 21821 26803 21879 26809
rect 22756 26784 22784 26880
rect 12584 26744 14412 26772
rect 16853 26775 16911 26781
rect 12584 26732 12590 26744
rect 16853 26741 16865 26775
rect 16899 26772 16911 26775
rect 17310 26772 17316 26784
rect 16899 26744 17316 26772
rect 16899 26741 16911 26744
rect 16853 26735 16911 26741
rect 17310 26732 17316 26744
rect 17368 26772 17374 26784
rect 19150 26772 19156 26784
rect 17368 26744 19156 26772
rect 17368 26732 17374 26744
rect 19150 26732 19156 26744
rect 19208 26732 19214 26784
rect 19613 26775 19671 26781
rect 19613 26741 19625 26775
rect 19659 26772 19671 26775
rect 19702 26772 19708 26784
rect 19659 26744 19708 26772
rect 19659 26741 19671 26744
rect 19613 26735 19671 26741
rect 19702 26732 19708 26744
rect 19760 26732 19766 26784
rect 22738 26732 22744 26784
rect 22796 26732 22802 26784
rect 22848 26772 22876 26936
rect 23382 26772 23388 26784
rect 22848 26744 23388 26772
rect 23382 26732 23388 26744
rect 23440 26732 23446 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 2225 26571 2283 26577
rect 2225 26537 2237 26571
rect 2271 26568 2283 26571
rect 3326 26568 3332 26580
rect 2271 26540 3332 26568
rect 2271 26537 2283 26540
rect 2225 26531 2283 26537
rect 3326 26528 3332 26540
rect 3384 26528 3390 26580
rect 5997 26571 6055 26577
rect 5997 26537 6009 26571
rect 6043 26568 6055 26571
rect 6086 26568 6092 26580
rect 6043 26540 6092 26568
rect 6043 26537 6055 26540
rect 5997 26531 6055 26537
rect 6086 26528 6092 26540
rect 6144 26528 6150 26580
rect 8202 26528 8208 26580
rect 8260 26568 8266 26580
rect 8389 26571 8447 26577
rect 8389 26568 8401 26571
rect 8260 26540 8401 26568
rect 8260 26528 8266 26540
rect 8389 26537 8401 26540
rect 8435 26537 8447 26571
rect 8389 26531 8447 26537
rect 9214 26528 9220 26580
rect 9272 26568 9278 26580
rect 9401 26571 9459 26577
rect 9401 26568 9413 26571
rect 9272 26540 9413 26568
rect 9272 26528 9278 26540
rect 9401 26537 9413 26540
rect 9447 26537 9459 26571
rect 9401 26531 9459 26537
rect 9490 26528 9496 26580
rect 9548 26528 9554 26580
rect 9766 26528 9772 26580
rect 9824 26528 9830 26580
rect 11054 26528 11060 26580
rect 11112 26568 11118 26580
rect 11149 26571 11207 26577
rect 11149 26568 11161 26571
rect 11112 26540 11161 26568
rect 11112 26528 11118 26540
rect 11149 26537 11161 26540
rect 11195 26537 11207 26571
rect 11149 26531 11207 26537
rect 15194 26528 15200 26580
rect 15252 26528 15258 26580
rect 16301 26571 16359 26577
rect 16301 26537 16313 26571
rect 16347 26568 16359 26571
rect 16574 26568 16580 26580
rect 16347 26540 16580 26568
rect 16347 26537 16359 26540
rect 16301 26531 16359 26537
rect 16574 26528 16580 26540
rect 16632 26528 16638 26580
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 19245 26571 19303 26577
rect 19245 26568 19257 26571
rect 18104 26540 19257 26568
rect 18104 26528 18110 26540
rect 19245 26537 19257 26540
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 19429 26571 19487 26577
rect 19429 26537 19441 26571
rect 19475 26568 19487 26571
rect 19702 26568 19708 26580
rect 19475 26540 19708 26568
rect 19475 26537 19487 26540
rect 19429 26531 19487 26537
rect 19702 26528 19708 26540
rect 19760 26568 19766 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 19760 26540 20177 26568
rect 19760 26528 19766 26540
rect 20165 26537 20177 26540
rect 20211 26568 20223 26571
rect 21637 26571 21695 26577
rect 21637 26568 21649 26571
rect 20211 26540 21649 26568
rect 20211 26537 20223 26540
rect 20165 26531 20223 26537
rect 21637 26537 21649 26540
rect 21683 26537 21695 26571
rect 21637 26531 21695 26537
rect 21821 26571 21879 26577
rect 21821 26537 21833 26571
rect 21867 26568 21879 26571
rect 21867 26540 22094 26568
rect 21867 26537 21879 26540
rect 21821 26531 21879 26537
rect 9309 26503 9367 26509
rect 9309 26469 9321 26503
rect 9355 26469 9367 26503
rect 9309 26463 9367 26469
rect 3605 26435 3663 26441
rect 3605 26401 3617 26435
rect 3651 26432 3663 26435
rect 3786 26432 3792 26444
rect 3651 26404 3792 26432
rect 3651 26401 3663 26404
rect 3605 26395 3663 26401
rect 3786 26392 3792 26404
rect 3844 26432 3850 26444
rect 3844 26404 4660 26432
rect 3844 26392 3850 26404
rect 4430 26324 4436 26376
rect 4488 26324 4494 26376
rect 4632 26373 4660 26404
rect 6362 26392 6368 26444
rect 6420 26432 6426 26444
rect 6549 26435 6607 26441
rect 6549 26432 6561 26435
rect 6420 26404 6561 26432
rect 6420 26392 6426 26404
rect 6549 26401 6561 26404
rect 6595 26401 6607 26435
rect 6549 26395 6607 26401
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26364 4675 26367
rect 6380 26364 6408 26392
rect 4663 26336 6408 26364
rect 6816 26367 6874 26373
rect 4663 26333 4675 26336
rect 4617 26327 4675 26333
rect 6816 26333 6828 26367
rect 6862 26364 6874 26367
rect 7190 26364 7196 26376
rect 6862 26336 7196 26364
rect 6862 26333 6874 26336
rect 6816 26327 6874 26333
rect 7190 26324 7196 26336
rect 7248 26324 7254 26376
rect 8021 26367 8079 26373
rect 8021 26333 8033 26367
rect 8067 26364 8079 26367
rect 8478 26364 8484 26376
rect 8067 26336 8484 26364
rect 8067 26333 8079 26336
rect 8021 26327 8079 26333
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 8941 26367 8999 26373
rect 8941 26333 8953 26367
rect 8987 26333 8999 26367
rect 9324 26364 9352 26463
rect 9508 26441 9536 26528
rect 9784 26500 9812 26528
rect 9784 26472 10548 26500
rect 9493 26435 9551 26441
rect 9493 26401 9505 26435
rect 9539 26401 9551 26435
rect 9493 26395 9551 26401
rect 9674 26392 9680 26444
rect 9732 26432 9738 26444
rect 10410 26432 10416 26444
rect 9732 26404 10416 26432
rect 9732 26392 9738 26404
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 10520 26441 10548 26472
rect 18690 26460 18696 26512
rect 18748 26500 18754 26512
rect 19981 26503 20039 26509
rect 19981 26500 19993 26503
rect 18748 26472 19993 26500
rect 18748 26460 18754 26472
rect 19981 26469 19993 26472
rect 20027 26469 20039 26503
rect 19981 26463 20039 26469
rect 10505 26435 10563 26441
rect 10505 26401 10517 26435
rect 10551 26401 10563 26435
rect 16850 26432 16856 26444
rect 10505 26395 10563 26401
rect 16500 26404 16856 26432
rect 9858 26364 9864 26376
rect 9324 26336 9864 26364
rect 8941 26327 8999 26333
rect 3360 26299 3418 26305
rect 3360 26265 3372 26299
rect 3406 26296 3418 26299
rect 3602 26296 3608 26308
rect 3406 26268 3608 26296
rect 3406 26265 3418 26268
rect 3360 26259 3418 26265
rect 3602 26256 3608 26268
rect 3660 26256 3666 26308
rect 4884 26299 4942 26305
rect 4884 26265 4896 26299
rect 4930 26265 4942 26299
rect 8205 26299 8263 26305
rect 8205 26296 8217 26299
rect 4884 26259 4942 26265
rect 7944 26268 8217 26296
rect 3878 26188 3884 26240
rect 3936 26188 3942 26240
rect 4798 26188 4804 26240
rect 4856 26228 4862 26240
rect 4908 26228 4936 26259
rect 7944 26237 7972 26268
rect 8205 26265 8217 26268
rect 8251 26296 8263 26299
rect 8386 26296 8392 26308
rect 8251 26268 8392 26296
rect 8251 26265 8263 26268
rect 8205 26259 8263 26265
rect 8386 26256 8392 26268
rect 8444 26296 8450 26308
rect 8956 26296 8984 26327
rect 9858 26324 9864 26336
rect 9916 26364 9922 26376
rect 9953 26367 10011 26373
rect 9953 26364 9965 26367
rect 9916 26336 9965 26364
rect 9916 26324 9922 26336
rect 9953 26333 9965 26336
rect 9999 26333 10011 26367
rect 9953 26327 10011 26333
rect 10962 26324 10968 26376
rect 11020 26324 11026 26376
rect 11974 26324 11980 26376
rect 12032 26364 12038 26376
rect 13722 26364 13728 26376
rect 12032 26336 13728 26364
rect 12032 26324 12038 26336
rect 13722 26324 13728 26336
rect 13780 26364 13786 26376
rect 15010 26364 15016 26376
rect 13780 26336 15016 26364
rect 13780 26324 13786 26336
rect 15010 26324 15016 26336
rect 15068 26324 15074 26376
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26364 15623 26367
rect 15654 26364 15660 26376
rect 15611 26336 15660 26364
rect 15611 26333 15623 26336
rect 15565 26327 15623 26333
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 15746 26324 15752 26376
rect 15804 26324 15810 26376
rect 16500 26373 16528 26404
rect 16850 26392 16856 26404
rect 16908 26392 16914 26444
rect 22066 26432 22094 26540
rect 22189 26503 22247 26509
rect 22189 26469 22201 26503
rect 22235 26500 22247 26503
rect 22278 26500 22284 26512
rect 22235 26472 22284 26500
rect 22235 26469 22247 26472
rect 22189 26463 22247 26469
rect 22278 26460 22284 26472
rect 22336 26500 22342 26512
rect 22336 26472 23336 26500
rect 22336 26460 22342 26472
rect 22738 26432 22744 26444
rect 22066 26404 22744 26432
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26333 16543 26367
rect 16485 26327 16543 26333
rect 16942 26324 16948 26376
rect 17000 26324 17006 26376
rect 17494 26324 17500 26376
rect 17552 26324 17558 26376
rect 22480 26373 22508 26404
rect 22738 26392 22744 26404
rect 22796 26392 22802 26444
rect 23308 26376 23336 26472
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 22465 26367 22523 26373
rect 19843 26336 20392 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 10980 26296 11008 26324
rect 8444 26268 8984 26296
rect 9784 26268 11008 26296
rect 8444 26256 8450 26268
rect 9784 26237 9812 26268
rect 11146 26256 11152 26308
rect 11204 26296 11210 26308
rect 12621 26299 12679 26305
rect 12621 26296 12633 26299
rect 11204 26268 12633 26296
rect 11204 26256 11210 26268
rect 12621 26265 12633 26268
rect 12667 26265 12679 26299
rect 12621 26259 12679 26265
rect 15381 26299 15439 26305
rect 15381 26265 15393 26299
rect 15427 26296 15439 26299
rect 15764 26296 15792 26324
rect 15427 26268 15792 26296
rect 15427 26265 15439 26268
rect 15381 26259 15439 26265
rect 16574 26256 16580 26308
rect 16632 26256 16638 26308
rect 16669 26299 16727 26305
rect 16669 26265 16681 26299
rect 16715 26265 16727 26299
rect 16669 26259 16727 26265
rect 16807 26299 16865 26305
rect 16807 26265 16819 26299
rect 16853 26296 16865 26299
rect 17512 26296 17540 26324
rect 20364 26308 20392 26336
rect 22465 26333 22477 26367
rect 22511 26333 22523 26367
rect 23109 26367 23167 26373
rect 23109 26364 23121 26367
rect 22465 26327 22523 26333
rect 22664 26336 23121 26364
rect 16853 26268 17540 26296
rect 19429 26299 19487 26305
rect 16853 26265 16865 26268
rect 16807 26259 16865 26265
rect 19429 26265 19441 26299
rect 19475 26296 19487 26299
rect 20162 26296 20168 26308
rect 19475 26268 20168 26296
rect 19475 26265 19487 26268
rect 19429 26259 19487 26265
rect 4856 26200 4936 26228
rect 7929 26231 7987 26237
rect 4856 26188 4862 26200
rect 7929 26197 7941 26231
rect 7975 26197 7987 26231
rect 7929 26191 7987 26197
rect 9769 26231 9827 26237
rect 9769 26197 9781 26231
rect 9815 26197 9827 26231
rect 9769 26191 9827 26197
rect 15562 26188 15568 26240
rect 15620 26228 15626 26240
rect 16684 26228 16712 26259
rect 20162 26256 20168 26268
rect 20220 26256 20226 26308
rect 20346 26256 20352 26308
rect 20404 26256 20410 26308
rect 21821 26299 21879 26305
rect 21821 26265 21833 26299
rect 21867 26296 21879 26299
rect 22094 26296 22100 26308
rect 21867 26268 22100 26296
rect 21867 26265 21879 26268
rect 21821 26259 21879 26265
rect 22094 26256 22100 26268
rect 22152 26296 22158 26308
rect 22664 26296 22692 26336
rect 23109 26333 23121 26336
rect 23155 26333 23167 26367
rect 23109 26327 23167 26333
rect 23290 26324 23296 26376
rect 23348 26324 23354 26376
rect 23385 26367 23443 26373
rect 23385 26333 23397 26367
rect 23431 26333 23443 26367
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 23385 26327 23443 26333
rect 23492 26336 23581 26364
rect 23400 26296 23428 26327
rect 22152 26268 22692 26296
rect 23124 26268 23428 26296
rect 22152 26256 22158 26268
rect 17770 26228 17776 26240
rect 15620 26200 17776 26228
rect 15620 26188 15626 26200
rect 17770 26188 17776 26200
rect 17828 26188 17834 26240
rect 20990 26188 20996 26240
rect 21048 26228 21054 26240
rect 22002 26228 22008 26240
rect 21048 26200 22008 26228
rect 21048 26188 21054 26200
rect 22002 26188 22008 26200
rect 22060 26188 22066 26240
rect 22370 26188 22376 26240
rect 22428 26188 22434 26240
rect 22922 26188 22928 26240
rect 22980 26228 22986 26240
rect 23124 26237 23152 26268
rect 23109 26231 23167 26237
rect 23109 26228 23121 26231
rect 22980 26200 23121 26228
rect 22980 26188 22986 26200
rect 23109 26197 23121 26200
rect 23155 26197 23167 26231
rect 23109 26191 23167 26197
rect 23382 26188 23388 26240
rect 23440 26228 23446 26240
rect 23492 26228 23520 26336
rect 23569 26333 23581 26336
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26364 28227 26367
rect 28445 26367 28503 26373
rect 28215 26336 28304 26364
rect 28215 26333 28227 26336
rect 28169 26327 28227 26333
rect 28276 26240 28304 26336
rect 28445 26333 28457 26367
rect 28491 26333 28503 26367
rect 28445 26327 28503 26333
rect 28460 26296 28488 26327
rect 28902 26296 28908 26308
rect 28460 26268 28908 26296
rect 28902 26256 28908 26268
rect 28960 26256 28966 26308
rect 23440 26200 23520 26228
rect 23440 26188 23446 26200
rect 23566 26188 23572 26240
rect 23624 26188 23630 26240
rect 26970 26188 26976 26240
rect 27028 26228 27034 26240
rect 28258 26228 28264 26240
rect 27028 26200 28264 26228
rect 27028 26188 27034 26200
rect 28258 26188 28264 26200
rect 28316 26188 28322 26240
rect 29178 26188 29184 26240
rect 29236 26228 29242 26240
rect 30558 26228 30564 26240
rect 29236 26200 30564 26228
rect 29236 26188 29242 26200
rect 30558 26188 30564 26200
rect 30616 26188 30622 26240
rect 1104 26138 38824 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 38824 26138
rect 1104 26064 38824 26086
rect 4341 26027 4399 26033
rect 4341 25993 4353 26027
rect 4387 26024 4399 26027
rect 4430 26024 4436 26036
rect 4387 25996 4436 26024
rect 4387 25993 4399 25996
rect 4341 25987 4399 25993
rect 4430 25984 4436 25996
rect 4488 25984 4494 26036
rect 4614 25984 4620 26036
rect 4672 25984 4678 26036
rect 4798 25984 4804 26036
rect 4856 26024 4862 26036
rect 5077 26027 5135 26033
rect 5077 26024 5089 26027
rect 4856 25996 5089 26024
rect 4856 25984 4862 25996
rect 5077 25993 5089 25996
rect 5123 25993 5135 26027
rect 5077 25987 5135 25993
rect 5534 25984 5540 26036
rect 5592 25984 5598 26036
rect 9674 25984 9680 26036
rect 9732 26024 9738 26036
rect 9769 26027 9827 26033
rect 9769 26024 9781 26027
rect 9732 25996 9781 26024
rect 9732 25984 9738 25996
rect 9769 25993 9781 25996
rect 9815 25993 9827 26027
rect 9769 25987 9827 25993
rect 9858 25984 9864 26036
rect 9916 25984 9922 26036
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 11238 26024 11244 26036
rect 10744 25996 11244 26024
rect 10744 25984 10750 25996
rect 11238 25984 11244 25996
rect 11296 25984 11302 26036
rect 13630 25984 13636 26036
rect 13688 25984 13694 26036
rect 13722 25984 13728 26036
rect 13780 25984 13786 26036
rect 13817 26027 13875 26033
rect 13817 25993 13829 26027
rect 13863 26024 13875 26027
rect 13906 26024 13912 26036
rect 13863 25996 13912 26024
rect 13863 25993 13875 25996
rect 13817 25987 13875 25993
rect 13906 25984 13912 25996
rect 13964 25984 13970 26036
rect 16850 25984 16856 26036
rect 16908 25984 16914 26036
rect 17497 26027 17555 26033
rect 17497 25993 17509 26027
rect 17543 26024 17555 26027
rect 17543 25996 18184 26024
rect 17543 25993 17555 25996
rect 17497 25987 17555 25993
rect 4632 25956 4660 25984
rect 4356 25928 4660 25956
rect 2774 25848 2780 25900
rect 2832 25897 2838 25900
rect 2832 25851 2844 25897
rect 2832 25848 2838 25851
rect 3510 25848 3516 25900
rect 3568 25848 3574 25900
rect 3786 25848 3792 25900
rect 3844 25848 3850 25900
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25820 3111 25823
rect 3804 25820 3832 25848
rect 3099 25792 3832 25820
rect 3099 25789 3111 25792
rect 3053 25783 3111 25789
rect 4062 25780 4068 25832
rect 4120 25780 4126 25832
rect 4356 25829 4384 25928
rect 4617 25891 4675 25897
rect 4617 25857 4629 25891
rect 4663 25857 4675 25891
rect 4617 25851 4675 25857
rect 5261 25891 5319 25897
rect 5261 25857 5273 25891
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 5445 25891 5503 25897
rect 5445 25857 5457 25891
rect 5491 25888 5503 25891
rect 5552 25888 5580 25984
rect 5491 25860 5580 25888
rect 5491 25857 5503 25860
rect 5445 25851 5503 25857
rect 4341 25823 4399 25829
rect 4341 25789 4353 25823
rect 4387 25789 4399 25823
rect 4341 25783 4399 25789
rect 4632 25752 4660 25851
rect 3068 25724 4660 25752
rect 1670 25644 1676 25696
rect 1728 25684 1734 25696
rect 3068 25684 3096 25724
rect 5276 25696 5304 25851
rect 5626 25848 5632 25900
rect 5684 25848 5690 25900
rect 7285 25891 7343 25897
rect 7285 25857 7297 25891
rect 7331 25888 7343 25891
rect 7834 25888 7840 25900
rect 7331 25860 7840 25888
rect 7331 25857 7343 25860
rect 7285 25851 7343 25857
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 9876 25897 9904 25984
rect 12161 25959 12219 25965
rect 12161 25956 12173 25959
rect 11072 25928 12173 25956
rect 11072 25897 11100 25928
rect 12161 25925 12173 25928
rect 12207 25925 12219 25959
rect 13648 25956 13676 25984
rect 12161 25919 12219 25925
rect 12268 25928 13676 25956
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25888 9367 25891
rect 9401 25891 9459 25897
rect 9401 25888 9413 25891
rect 9355 25860 9413 25888
rect 9355 25857 9367 25860
rect 9309 25851 9367 25857
rect 9401 25857 9413 25860
rect 9447 25857 9459 25891
rect 9401 25851 9459 25857
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9861 25891 9919 25897
rect 9861 25857 9873 25891
rect 9907 25857 9919 25891
rect 9861 25851 9919 25857
rect 11057 25891 11115 25897
rect 11057 25857 11069 25891
rect 11103 25857 11115 25891
rect 11057 25851 11115 25857
rect 11333 25891 11391 25897
rect 11333 25857 11345 25891
rect 11379 25888 11391 25891
rect 11606 25888 11612 25900
rect 11379 25860 11612 25888
rect 11379 25857 11391 25860
rect 11333 25851 11391 25857
rect 5537 25823 5595 25829
rect 5537 25789 5549 25823
rect 5583 25820 5595 25823
rect 5644 25820 5672 25848
rect 5583 25792 5672 25820
rect 5583 25789 5595 25792
rect 5537 25783 5595 25789
rect 8662 25780 8668 25832
rect 8720 25780 8726 25832
rect 6914 25712 6920 25764
rect 6972 25752 6978 25764
rect 7285 25755 7343 25761
rect 7285 25752 7297 25755
rect 6972 25724 7297 25752
rect 6972 25712 6978 25724
rect 7285 25721 7297 25724
rect 7331 25752 7343 25755
rect 8202 25752 8208 25764
rect 7331 25724 8208 25752
rect 7331 25721 7343 25724
rect 7285 25715 7343 25721
rect 8202 25712 8208 25724
rect 8260 25752 8266 25764
rect 9600 25752 9628 25851
rect 11606 25848 11612 25860
rect 11664 25848 11670 25900
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25888 11759 25891
rect 12268 25888 12296 25928
rect 11747 25860 12296 25888
rect 12345 25894 12403 25897
rect 12434 25894 12440 25900
rect 12345 25891 12440 25894
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 12345 25857 12357 25891
rect 12391 25866 12440 25891
rect 12391 25857 12403 25866
rect 12345 25851 12403 25857
rect 12434 25848 12440 25866
rect 12492 25848 12498 25900
rect 12526 25848 12532 25900
rect 12584 25888 12590 25900
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 12584 25860 13277 25888
rect 12584 25848 12590 25860
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 13446 25848 13452 25900
rect 13504 25848 13510 25900
rect 13541 25891 13599 25897
rect 13541 25857 13553 25891
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 13633 25891 13691 25897
rect 13633 25857 13645 25891
rect 13679 25888 13691 25891
rect 13740 25888 13768 25984
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25925 17831 25959
rect 17773 25919 17831 25925
rect 18156 25956 18184 25996
rect 18414 25984 18420 26036
rect 18472 25984 18478 26036
rect 19334 25984 19340 26036
rect 19392 26024 19398 26036
rect 20070 26024 20076 26036
rect 19392 25996 20076 26024
rect 19392 25984 19398 25996
rect 20070 25984 20076 25996
rect 20128 26024 20134 26036
rect 20625 26027 20683 26033
rect 20625 26024 20637 26027
rect 20128 25996 20637 26024
rect 20128 25984 20134 25996
rect 20625 25993 20637 25996
rect 20671 25993 20683 26027
rect 20625 25987 20683 25993
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 22370 26024 22376 26036
rect 22235 25996 22376 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 18432 25956 18460 25984
rect 18156 25928 18460 25956
rect 13679 25860 13768 25888
rect 16301 25891 16359 25897
rect 13679 25857 13691 25860
rect 13633 25851 13691 25857
rect 16301 25857 16313 25891
rect 16347 25857 16359 25891
rect 16301 25851 16359 25857
rect 16485 25891 16543 25897
rect 16485 25857 16497 25891
rect 16531 25888 16543 25891
rect 16758 25888 16764 25900
rect 16531 25860 16764 25888
rect 16531 25857 16543 25860
rect 16485 25851 16543 25857
rect 10873 25823 10931 25829
rect 10873 25789 10885 25823
rect 10919 25820 10931 25823
rect 11793 25823 11851 25829
rect 11793 25820 11805 25823
rect 10919 25792 11805 25820
rect 10919 25789 10931 25792
rect 10873 25783 10931 25789
rect 11793 25789 11805 25792
rect 11839 25789 11851 25823
rect 11793 25783 11851 25789
rect 12250 25780 12256 25832
rect 12308 25820 12314 25832
rect 12621 25823 12679 25829
rect 12621 25820 12633 25823
rect 12308 25792 12633 25820
rect 12308 25780 12314 25792
rect 12621 25789 12633 25792
rect 12667 25820 12679 25823
rect 13354 25820 13360 25832
rect 12667 25792 13360 25820
rect 12667 25789 12679 25792
rect 12621 25783 12679 25789
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 13556 25752 13584 25851
rect 8260 25724 9628 25752
rect 8260 25712 8266 25724
rect 3142 25684 3148 25696
rect 1728 25656 3148 25684
rect 1728 25644 1734 25656
rect 3142 25644 3148 25656
rect 3200 25644 3206 25696
rect 3694 25644 3700 25696
rect 3752 25684 3758 25696
rect 4525 25687 4583 25693
rect 4525 25684 4537 25687
rect 3752 25656 4537 25684
rect 3752 25644 3758 25656
rect 4525 25653 4537 25656
rect 4571 25653 4583 25687
rect 4525 25647 4583 25653
rect 5258 25644 5264 25696
rect 5316 25644 5322 25696
rect 9398 25644 9404 25696
rect 9456 25644 9462 25696
rect 9600 25684 9628 25724
rect 12636 25724 13584 25752
rect 12636 25696 12664 25724
rect 10042 25684 10048 25696
rect 9600 25656 10048 25684
rect 10042 25644 10048 25656
rect 10100 25684 10106 25696
rect 11514 25684 11520 25696
rect 10100 25656 11520 25684
rect 10100 25644 10106 25656
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 11882 25644 11888 25696
rect 11940 25684 11946 25696
rect 11977 25687 12035 25693
rect 11977 25684 11989 25687
rect 11940 25656 11989 25684
rect 11940 25644 11946 25656
rect 11977 25653 11989 25656
rect 12023 25653 12035 25687
rect 11977 25647 12035 25653
rect 12529 25687 12587 25693
rect 12529 25653 12541 25687
rect 12575 25684 12587 25687
rect 12618 25684 12624 25696
rect 12575 25656 12624 25684
rect 12575 25653 12587 25656
rect 12529 25647 12587 25653
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 15010 25644 15016 25696
rect 15068 25684 15074 25696
rect 16117 25687 16175 25693
rect 16117 25684 16129 25687
rect 15068 25656 16129 25684
rect 15068 25644 15074 25656
rect 16117 25653 16129 25656
rect 16163 25653 16175 25687
rect 16316 25684 16344 25851
rect 16758 25848 16764 25860
rect 16816 25888 16822 25900
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 16816 25860 17141 25888
rect 16816 25848 16822 25860
rect 17129 25857 17141 25860
rect 17175 25888 17187 25891
rect 17788 25888 17816 25919
rect 18156 25897 18184 25928
rect 20806 25916 20812 25968
rect 20864 25956 20870 25968
rect 21174 25956 21180 25968
rect 20864 25928 21180 25956
rect 20864 25916 20870 25928
rect 21174 25916 21180 25928
rect 21232 25956 21238 25968
rect 21361 25959 21419 25965
rect 21361 25956 21373 25959
rect 21232 25928 21373 25956
rect 21232 25916 21238 25928
rect 21361 25925 21373 25928
rect 21407 25925 21419 25959
rect 22296 25956 22324 25996
rect 22370 25984 22376 25996
rect 22428 25984 22434 26036
rect 23290 25984 23296 26036
rect 23348 26024 23354 26036
rect 25501 26027 25559 26033
rect 25501 26024 25513 26027
rect 23348 25996 25513 26024
rect 23348 25984 23354 25996
rect 25501 25993 25513 25996
rect 25547 25993 25559 26027
rect 30374 26024 30380 26036
rect 25501 25987 25559 25993
rect 29472 25996 30380 26024
rect 23382 25956 23388 25968
rect 21361 25919 21419 25925
rect 21468 25928 22324 25956
rect 22480 25928 23388 25956
rect 21468 25900 21496 25928
rect 17175 25860 17816 25888
rect 18141 25891 18199 25897
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 18141 25857 18153 25891
rect 18187 25857 18199 25891
rect 18141 25851 18199 25857
rect 18230 25848 18236 25900
rect 18288 25888 18294 25900
rect 18325 25891 18383 25897
rect 18325 25888 18337 25891
rect 18288 25860 18337 25888
rect 18288 25848 18294 25860
rect 18325 25857 18337 25860
rect 18371 25888 18383 25891
rect 18414 25888 18420 25900
rect 18371 25860 18420 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25857 18567 25891
rect 18509 25851 18567 25857
rect 18693 25891 18751 25897
rect 18693 25857 18705 25891
rect 18739 25888 18751 25891
rect 19242 25888 19248 25900
rect 18739 25860 19248 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 17037 25823 17095 25829
rect 17037 25789 17049 25823
rect 17083 25789 17095 25823
rect 18524 25820 18552 25851
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20533 25891 20591 25897
rect 20533 25888 20545 25891
rect 20220 25860 20545 25888
rect 20220 25848 20226 25860
rect 20533 25857 20545 25860
rect 20579 25857 20591 25891
rect 20533 25851 20591 25857
rect 20714 25848 20720 25900
rect 20772 25848 20778 25900
rect 20898 25848 20904 25900
rect 20956 25848 20962 25900
rect 21266 25848 21272 25900
rect 21324 25848 21330 25900
rect 21450 25848 21456 25900
rect 21508 25848 21514 25900
rect 22278 25898 22284 25900
rect 21821 25891 21879 25897
rect 21821 25857 21833 25891
rect 21867 25888 21879 25891
rect 22112 25888 22284 25898
rect 21867 25870 22284 25888
rect 21867 25860 22140 25870
rect 21867 25857 21879 25860
rect 21821 25851 21879 25857
rect 22278 25848 22284 25870
rect 22336 25848 22342 25900
rect 19150 25820 19156 25832
rect 18524 25792 19156 25820
rect 17037 25783 17095 25789
rect 17052 25752 17080 25783
rect 19150 25780 19156 25792
rect 19208 25780 19214 25832
rect 21284 25820 21312 25848
rect 22480 25820 22508 25928
rect 23382 25916 23388 25928
rect 23440 25916 23446 25968
rect 23566 25916 23572 25968
rect 23624 25956 23630 25968
rect 24366 25959 24424 25965
rect 24366 25956 24378 25959
rect 23624 25928 24378 25956
rect 23624 25916 23630 25928
rect 24366 25925 24378 25928
rect 24412 25925 24424 25959
rect 29472 25956 29500 25996
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 30558 25984 30564 26036
rect 30616 26024 30622 26036
rect 35434 26024 35440 26036
rect 30616 25996 35440 26024
rect 30616 25984 30622 25996
rect 35434 25984 35440 25996
rect 35492 25984 35498 26036
rect 24366 25919 24424 25925
rect 25148 25928 29500 25956
rect 22554 25848 22560 25900
rect 22612 25888 22618 25900
rect 23762 25891 23820 25897
rect 23762 25888 23774 25891
rect 22612 25860 23774 25888
rect 22612 25848 22618 25860
rect 23762 25857 23774 25860
rect 23808 25857 23820 25891
rect 23762 25851 23820 25857
rect 23934 25848 23940 25900
rect 23992 25888 23998 25900
rect 24029 25891 24087 25897
rect 24029 25888 24041 25891
rect 23992 25860 24041 25888
rect 23992 25848 23998 25860
rect 24029 25857 24041 25860
rect 24075 25888 24087 25891
rect 24121 25891 24179 25897
rect 24121 25888 24133 25891
rect 24075 25860 24133 25888
rect 24075 25857 24087 25860
rect 24029 25851 24087 25857
rect 24121 25857 24133 25860
rect 24167 25857 24179 25891
rect 24121 25851 24179 25857
rect 25148 25832 25176 25928
rect 28261 25891 28319 25897
rect 28261 25857 28273 25891
rect 28307 25888 28319 25891
rect 28350 25888 28356 25900
rect 28307 25860 28356 25888
rect 28307 25857 28319 25860
rect 28261 25851 28319 25857
rect 28350 25848 28356 25860
rect 28408 25848 28414 25900
rect 29089 25891 29147 25897
rect 29089 25857 29101 25891
rect 29135 25888 29147 25891
rect 29178 25888 29184 25900
rect 29135 25860 29184 25888
rect 29135 25857 29147 25860
rect 29089 25851 29147 25857
rect 29178 25848 29184 25860
rect 29236 25848 29242 25900
rect 29472 25897 29500 25928
rect 30466 25916 30472 25968
rect 30524 25916 30530 25968
rect 29457 25891 29515 25897
rect 29457 25857 29469 25891
rect 29503 25857 29515 25891
rect 29457 25851 29515 25857
rect 21284 25792 22508 25820
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 29365 25823 29423 25829
rect 29365 25789 29377 25823
rect 29411 25820 29423 25823
rect 29411 25792 29592 25820
rect 29411 25789 29423 25792
rect 29365 25783 29423 25789
rect 17310 25752 17316 25764
rect 17052 25724 17316 25752
rect 17310 25712 17316 25724
rect 17368 25752 17374 25764
rect 22649 25755 22707 25761
rect 22649 25752 22661 25755
rect 17368 25724 17816 25752
rect 17368 25712 17374 25724
rect 16574 25684 16580 25696
rect 16316 25656 16580 25684
rect 16117 25647 16175 25653
rect 16574 25644 16580 25656
rect 16632 25684 16638 25696
rect 17494 25684 17500 25696
rect 16632 25656 17500 25684
rect 16632 25644 16638 25656
rect 17494 25644 17500 25656
rect 17552 25644 17558 25696
rect 17586 25644 17592 25696
rect 17644 25644 17650 25696
rect 17788 25693 17816 25724
rect 22204 25724 22661 25752
rect 17773 25687 17831 25693
rect 17773 25653 17785 25687
rect 17819 25653 17831 25687
rect 17773 25647 17831 25653
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 19978 25684 19984 25696
rect 19484 25656 19984 25684
rect 19484 25644 19490 25656
rect 19978 25644 19984 25656
rect 20036 25644 20042 25696
rect 21085 25687 21143 25693
rect 21085 25653 21097 25687
rect 21131 25684 21143 25687
rect 21910 25684 21916 25696
rect 21131 25656 21916 25684
rect 21131 25653 21143 25656
rect 21085 25647 21143 25653
rect 21910 25644 21916 25656
rect 21968 25644 21974 25696
rect 22094 25644 22100 25696
rect 22152 25684 22158 25696
rect 22204 25693 22232 25724
rect 22649 25721 22661 25724
rect 22695 25721 22707 25755
rect 22649 25715 22707 25721
rect 22189 25687 22247 25693
rect 22189 25684 22201 25687
rect 22152 25656 22201 25684
rect 22152 25644 22158 25656
rect 22189 25653 22201 25656
rect 22235 25653 22247 25687
rect 22189 25647 22247 25653
rect 22370 25644 22376 25696
rect 22428 25644 22434 25696
rect 28258 25644 28264 25696
rect 28316 25684 28322 25696
rect 29564 25684 29592 25792
rect 29730 25780 29736 25832
rect 29788 25780 29794 25832
rect 33318 25780 33324 25832
rect 33376 25780 33382 25832
rect 33336 25752 33364 25780
rect 30760 25724 33364 25752
rect 30760 25684 30788 25724
rect 28316 25656 30788 25684
rect 28316 25644 28322 25656
rect 31202 25644 31208 25696
rect 31260 25644 31266 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 2593 25483 2651 25489
rect 2593 25449 2605 25483
rect 2639 25480 2651 25483
rect 2774 25480 2780 25492
rect 2639 25452 2780 25480
rect 2639 25449 2651 25452
rect 2593 25443 2651 25449
rect 2774 25440 2780 25452
rect 2832 25440 2838 25492
rect 3034 25483 3092 25489
rect 3034 25449 3046 25483
rect 3080 25480 3092 25483
rect 3326 25480 3332 25492
rect 3080 25452 3332 25480
rect 3080 25449 3092 25452
rect 3034 25443 3092 25449
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 3510 25440 3516 25492
rect 3568 25440 3574 25492
rect 3602 25440 3608 25492
rect 3660 25480 3666 25492
rect 3881 25483 3939 25489
rect 3881 25480 3893 25483
rect 3660 25452 3893 25480
rect 3660 25440 3666 25452
rect 3881 25449 3893 25452
rect 3927 25449 3939 25483
rect 3881 25443 3939 25449
rect 8021 25483 8079 25489
rect 8021 25449 8033 25483
rect 8067 25480 8079 25483
rect 8662 25480 8668 25492
rect 8067 25452 8668 25480
rect 8067 25449 8079 25452
rect 8021 25443 8079 25449
rect 8662 25440 8668 25452
rect 8720 25440 8726 25492
rect 9858 25480 9864 25492
rect 9140 25452 9864 25480
rect 3142 25372 3148 25424
rect 3200 25372 3206 25424
rect 9140 25412 9168 25452
rect 9858 25440 9864 25452
rect 9916 25480 9922 25492
rect 10505 25483 10563 25489
rect 10505 25480 10517 25483
rect 9916 25452 10517 25480
rect 9916 25440 9922 25452
rect 10505 25449 10517 25452
rect 10551 25480 10563 25483
rect 10962 25480 10968 25492
rect 10551 25452 10968 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12618 25440 12624 25492
rect 12676 25440 12682 25492
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 13446 25480 13452 25492
rect 12851 25452 13452 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 13446 25440 13452 25452
rect 13504 25440 13510 25492
rect 15010 25440 15016 25492
rect 15068 25440 15074 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15378 25480 15384 25492
rect 15151 25452 15384 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15378 25440 15384 25452
rect 15436 25440 15442 25492
rect 15565 25483 15623 25489
rect 15565 25449 15577 25483
rect 15611 25480 15623 25483
rect 15611 25452 16252 25480
rect 15611 25449 15623 25452
rect 15565 25443 15623 25449
rect 7760 25384 9168 25412
rect 3234 25304 3240 25356
rect 3292 25304 3298 25356
rect 4062 25344 4068 25356
rect 3804 25316 4068 25344
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25245 1915 25279
rect 1857 25239 1915 25245
rect 934 25100 940 25152
rect 992 25140 998 25152
rect 1673 25143 1731 25149
rect 1673 25140 1685 25143
rect 992 25112 1685 25140
rect 992 25100 998 25112
rect 1673 25109 1685 25112
rect 1719 25109 1731 25143
rect 1872 25140 1900 25239
rect 1946 25236 1952 25288
rect 2004 25236 2010 25288
rect 3804 25285 3832 25316
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 3789 25279 3847 25285
rect 3789 25245 3801 25279
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 3878 25236 3884 25288
rect 3936 25276 3942 25288
rect 3973 25279 4031 25285
rect 3973 25276 3985 25279
rect 3936 25248 3985 25276
rect 3936 25236 3942 25248
rect 3973 25245 3985 25248
rect 4019 25245 4031 25279
rect 3973 25239 4031 25245
rect 5258 25236 5264 25288
rect 5316 25236 5322 25288
rect 5442 25236 5448 25288
rect 5500 25236 5506 25288
rect 5534 25236 5540 25288
rect 5592 25236 5598 25288
rect 7760 25285 7788 25384
rect 11606 25372 11612 25424
rect 11664 25412 11670 25424
rect 12636 25412 12664 25440
rect 11664 25384 12664 25412
rect 14369 25415 14427 25421
rect 11664 25372 11670 25384
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25344 7895 25347
rect 8018 25344 8024 25356
rect 7883 25316 8024 25344
rect 7883 25313 7895 25316
rect 7837 25307 7895 25313
rect 8018 25304 8024 25316
rect 8076 25304 8082 25356
rect 11900 25353 11928 25384
rect 14369 25381 14381 25415
rect 14415 25412 14427 25415
rect 15028 25412 15056 25440
rect 14415 25384 15056 25412
rect 14415 25381 14427 25384
rect 14369 25375 14427 25381
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25313 11943 25347
rect 11885 25307 11943 25313
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12710 25344 12716 25356
rect 12667 25316 12716 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 14185 25347 14243 25353
rect 14185 25313 14197 25347
rect 14231 25344 14243 25347
rect 14231 25316 14688 25344
rect 14231 25313 14243 25316
rect 14185 25307 14243 25313
rect 7745 25279 7803 25285
rect 7745 25245 7757 25279
rect 7791 25245 7803 25279
rect 7745 25239 7803 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25276 9183 25279
rect 9950 25276 9956 25288
rect 9171 25248 9956 25276
rect 9171 25245 9183 25248
rect 9125 25239 9183 25245
rect 9950 25236 9956 25248
rect 10008 25236 10014 25288
rect 10778 25236 10784 25288
rect 10836 25236 10842 25288
rect 11238 25236 11244 25288
rect 11296 25276 11302 25288
rect 11793 25279 11851 25285
rect 11793 25276 11805 25279
rect 11296 25248 11805 25276
rect 11296 25236 11302 25248
rect 11793 25245 11805 25248
rect 11839 25276 11851 25279
rect 12250 25276 12256 25288
rect 11839 25248 12256 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12529 25239 12587 25245
rect 2866 25168 2872 25220
rect 2924 25168 2930 25220
rect 5276 25208 5304 25236
rect 7834 25208 7840 25220
rect 4724 25180 5212 25208
rect 5276 25180 7840 25208
rect 4724 25140 4752 25180
rect 1872 25112 4752 25140
rect 1673 25103 1731 25109
rect 4798 25100 4804 25152
rect 4856 25140 4862 25152
rect 5077 25143 5135 25149
rect 5077 25140 5089 25143
rect 4856 25112 5089 25140
rect 4856 25100 4862 25112
rect 5077 25109 5089 25112
rect 5123 25109 5135 25143
rect 5184 25140 5212 25180
rect 7834 25168 7840 25180
rect 7892 25168 7898 25220
rect 9398 25217 9404 25220
rect 9392 25208 9404 25217
rect 9359 25180 9404 25208
rect 9392 25171 9404 25180
rect 9398 25168 9404 25171
rect 9456 25168 9462 25220
rect 9508 25180 11468 25208
rect 9508 25140 9536 25180
rect 11440 25152 11468 25180
rect 12434 25168 12440 25220
rect 12492 25208 12498 25220
rect 12544 25208 12572 25239
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14185 25211 14243 25217
rect 14185 25208 14197 25211
rect 12492 25180 14197 25208
rect 12492 25168 12498 25180
rect 14185 25177 14197 25180
rect 14231 25177 14243 25211
rect 14185 25171 14243 25177
rect 5184 25112 9536 25140
rect 5077 25103 5135 25109
rect 11330 25100 11336 25152
rect 11388 25100 11394 25152
rect 11422 25100 11428 25152
rect 11480 25100 11486 25152
rect 12161 25143 12219 25149
rect 12161 25109 12173 25143
rect 12207 25140 12219 25143
rect 12710 25140 12716 25152
rect 12207 25112 12716 25140
rect 12207 25109 12219 25112
rect 12161 25103 12219 25109
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 14660 25140 14688 25316
rect 14752 25285 14780 25384
rect 14829 25347 14887 25353
rect 14829 25313 14841 25347
rect 14875 25344 14887 25347
rect 16025 25347 16083 25353
rect 16025 25344 16037 25347
rect 14875 25316 16037 25344
rect 14875 25313 14887 25316
rect 14829 25307 14887 25313
rect 16025 25313 16037 25316
rect 16071 25313 16083 25347
rect 16025 25307 16083 25313
rect 14737 25279 14795 25285
rect 14737 25245 14749 25279
rect 14783 25245 14795 25279
rect 15286 25276 15292 25288
rect 14737 25239 14795 25245
rect 15212 25248 15292 25276
rect 14826 25168 14832 25220
rect 14884 25208 14890 25220
rect 15212 25217 15240 25248
rect 15286 25236 15292 25248
rect 15344 25276 15350 25288
rect 15657 25279 15715 25285
rect 15657 25276 15669 25279
rect 15344 25248 15669 25276
rect 15344 25236 15350 25248
rect 15657 25245 15669 25248
rect 15703 25245 15715 25279
rect 15657 25239 15715 25245
rect 15746 25236 15752 25288
rect 15804 25276 15810 25288
rect 15841 25279 15899 25285
rect 15841 25276 15853 25279
rect 15804 25248 15853 25276
rect 15804 25236 15810 25248
rect 15841 25245 15853 25248
rect 15887 25245 15899 25279
rect 15841 25239 15899 25245
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25245 15991 25279
rect 15933 25239 15991 25245
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16224 25276 16252 25452
rect 16758 25440 16764 25492
rect 16816 25440 16822 25492
rect 17310 25440 17316 25492
rect 17368 25440 17374 25492
rect 17494 25440 17500 25492
rect 17552 25440 17558 25492
rect 17586 25440 17592 25492
rect 17644 25440 17650 25492
rect 20714 25440 20720 25492
rect 20772 25440 20778 25492
rect 20898 25440 20904 25492
rect 20956 25440 20962 25492
rect 22094 25440 22100 25492
rect 22152 25480 22158 25492
rect 22152 25452 22324 25480
rect 22152 25440 22158 25452
rect 17034 25344 17040 25356
rect 16684 25316 17040 25344
rect 16163 25248 16252 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 15197 25211 15255 25217
rect 15197 25208 15209 25211
rect 14884 25180 15209 25208
rect 14884 25168 14890 25180
rect 15197 25177 15209 25180
rect 15243 25177 15255 25211
rect 15197 25171 15255 25177
rect 15378 25168 15384 25220
rect 15436 25168 15442 25220
rect 15948 25208 15976 25239
rect 16298 25236 16304 25288
rect 16356 25276 16362 25288
rect 16684 25285 16712 25316
rect 17034 25304 17040 25316
rect 17092 25344 17098 25356
rect 17092 25316 17172 25344
rect 17092 25304 17098 25316
rect 17144 25285 17172 25316
rect 17604 25285 17632 25440
rect 20622 25412 20628 25424
rect 19812 25384 20628 25412
rect 19812 25285 19840 25384
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 20732 25412 20760 25440
rect 20993 25415 21051 25421
rect 20993 25412 21005 25415
rect 20732 25384 21005 25412
rect 20993 25381 21005 25384
rect 21039 25381 21051 25415
rect 20993 25375 21051 25381
rect 21361 25347 21419 25353
rect 21361 25344 21373 25347
rect 20272 25316 21373 25344
rect 20272 25288 20300 25316
rect 21361 25313 21373 25316
rect 21407 25313 21419 25347
rect 21361 25307 21419 25313
rect 16669 25279 16727 25285
rect 16669 25276 16681 25279
rect 16356 25248 16681 25276
rect 16356 25236 16362 25248
rect 16669 25245 16681 25248
rect 16715 25245 16727 25279
rect 16669 25239 16727 25245
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25245 16911 25279
rect 16853 25239 16911 25245
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17589 25279 17647 25285
rect 17589 25245 17601 25279
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 15764 25180 15976 25208
rect 16868 25208 16896 25239
rect 20070 25236 20076 25288
rect 20128 25276 20134 25288
rect 20165 25279 20223 25285
rect 20165 25276 20177 25279
rect 20128 25248 20177 25276
rect 20128 25236 20134 25248
rect 20165 25245 20177 25248
rect 20211 25245 20223 25279
rect 20165 25239 20223 25245
rect 20254 25236 20260 25288
rect 20312 25236 20318 25288
rect 20533 25279 20591 25285
rect 20533 25245 20545 25279
rect 20579 25276 20591 25279
rect 21174 25276 21180 25288
rect 20579 25248 21180 25276
rect 20579 25245 20591 25248
rect 20533 25239 20591 25245
rect 21174 25236 21180 25248
rect 21232 25236 21238 25288
rect 22094 25236 22100 25288
rect 22152 25236 22158 25288
rect 22296 25276 22324 25452
rect 22370 25440 22376 25492
rect 22428 25440 22434 25492
rect 22554 25440 22560 25492
rect 22612 25440 22618 25492
rect 23382 25440 23388 25492
rect 23440 25440 23446 25492
rect 29730 25440 29736 25492
rect 29788 25440 29794 25492
rect 30466 25440 30472 25492
rect 30524 25480 30530 25492
rect 30561 25483 30619 25489
rect 30561 25480 30573 25483
rect 30524 25452 30573 25480
rect 30524 25440 30530 25452
rect 30561 25449 30573 25452
rect 30607 25449 30619 25483
rect 30561 25443 30619 25449
rect 22388 25353 22416 25440
rect 28074 25372 28080 25424
rect 28132 25412 28138 25424
rect 28261 25415 28319 25421
rect 28261 25412 28273 25415
rect 28132 25384 28273 25412
rect 28132 25372 28138 25384
rect 28261 25381 28273 25384
rect 28307 25412 28319 25415
rect 35434 25412 35440 25424
rect 28307 25384 35440 25412
rect 28307 25381 28319 25384
rect 28261 25375 28319 25381
rect 35434 25372 35440 25384
rect 35492 25372 35498 25424
rect 22373 25347 22431 25353
rect 22373 25313 22385 25347
rect 22419 25313 22431 25347
rect 22373 25307 22431 25313
rect 22480 25316 23244 25344
rect 22480 25285 22508 25316
rect 22465 25279 22523 25285
rect 22465 25276 22477 25279
rect 22296 25248 22477 25276
rect 22465 25245 22477 25248
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 22738 25236 22744 25288
rect 22796 25236 22802 25288
rect 22922 25236 22928 25288
rect 22980 25236 22986 25288
rect 23216 25285 23244 25316
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25245 23259 25279
rect 23201 25239 23259 25245
rect 23290 25236 23296 25288
rect 23348 25236 23354 25288
rect 25130 25236 25136 25288
rect 25188 25276 25194 25288
rect 25409 25279 25467 25285
rect 25409 25276 25421 25279
rect 25188 25248 25421 25276
rect 25188 25236 25194 25248
rect 25409 25245 25421 25248
rect 25455 25245 25467 25279
rect 25409 25239 25467 25245
rect 26970 25236 26976 25288
rect 27028 25276 27034 25288
rect 27249 25279 27307 25285
rect 27249 25276 27261 25279
rect 27028 25248 27261 25276
rect 27028 25236 27034 25248
rect 27249 25245 27261 25248
rect 27295 25245 27307 25279
rect 27249 25239 27307 25245
rect 27525 25279 27583 25285
rect 27525 25245 27537 25279
rect 27571 25245 27583 25279
rect 27525 25239 27583 25245
rect 16945 25211 17003 25217
rect 16945 25208 16957 25211
rect 16868 25180 16957 25208
rect 15764 25149 15792 25180
rect 16945 25177 16957 25180
rect 16991 25208 17003 25211
rect 19889 25211 19947 25217
rect 16991 25180 17172 25208
rect 16991 25177 17003 25180
rect 16945 25171 17003 25177
rect 17144 25152 17172 25180
rect 19889 25177 19901 25211
rect 19935 25177 19947 25211
rect 19889 25171 19947 25177
rect 19981 25211 20039 25217
rect 19981 25177 19993 25211
rect 20027 25208 20039 25211
rect 20742 25211 20800 25217
rect 20742 25208 20754 25211
rect 20027 25180 20754 25208
rect 20027 25177 20039 25180
rect 19981 25171 20039 25177
rect 20742 25177 20754 25180
rect 20788 25208 20800 25211
rect 22833 25211 22891 25217
rect 22833 25208 22845 25211
rect 20788 25180 22845 25208
rect 20788 25177 20800 25180
rect 20742 25171 20800 25177
rect 22833 25177 22845 25180
rect 22879 25177 22891 25211
rect 22833 25171 22891 25177
rect 23017 25211 23075 25217
rect 23017 25177 23029 25211
rect 23063 25208 23075 25211
rect 23308 25208 23336 25236
rect 23063 25180 23336 25208
rect 23063 25177 23075 25180
rect 23017 25171 23075 25177
rect 15749 25143 15807 25149
rect 15749 25140 15761 25143
rect 14660 25112 15761 25140
rect 15749 25109 15761 25112
rect 15795 25109 15807 25143
rect 15749 25103 15807 25109
rect 17126 25100 17132 25152
rect 17184 25100 17190 25152
rect 19058 25100 19064 25152
rect 19116 25140 19122 25152
rect 19613 25143 19671 25149
rect 19613 25140 19625 25143
rect 19116 25112 19625 25140
rect 19116 25100 19122 25112
rect 19613 25109 19625 25112
rect 19659 25109 19671 25143
rect 19904 25140 19932 25171
rect 25682 25168 25688 25220
rect 25740 25168 25746 25220
rect 26418 25168 26424 25220
rect 26476 25168 26482 25220
rect 27540 25208 27568 25239
rect 29546 25236 29552 25288
rect 29604 25236 29610 25288
rect 30469 25279 30527 25285
rect 30469 25245 30481 25279
rect 30515 25276 30527 25279
rect 30515 25248 30696 25276
rect 30515 25245 30527 25248
rect 30469 25239 30527 25245
rect 27172 25180 27568 25208
rect 27172 25152 27200 25180
rect 30668 25152 30696 25248
rect 20162 25140 20168 25152
rect 19904 25112 20168 25140
rect 19613 25103 19671 25109
rect 20162 25100 20168 25112
rect 20220 25100 20226 25152
rect 20346 25100 20352 25152
rect 20404 25140 20410 25152
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 20404 25112 20637 25140
rect 20404 25100 20410 25112
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 27154 25100 27160 25152
rect 27212 25100 27218 25152
rect 30650 25100 30656 25152
rect 30708 25100 30714 25152
rect 1104 25050 38824 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 38824 25050
rect 1104 24976 38824 24998
rect 1946 24896 1952 24948
rect 2004 24896 2010 24948
rect 2409 24939 2467 24945
rect 2409 24905 2421 24939
rect 2455 24936 2467 24939
rect 3694 24936 3700 24948
rect 2455 24908 3700 24936
rect 2455 24905 2467 24908
rect 2409 24899 2467 24905
rect 2130 24868 2136 24880
rect 1504 24840 2136 24868
rect 1504 24741 1532 24840
rect 2130 24828 2136 24840
rect 2188 24868 2194 24880
rect 2424 24868 2452 24899
rect 3694 24896 3700 24908
rect 3752 24896 3758 24948
rect 5534 24896 5540 24948
rect 5592 24936 5598 24948
rect 5997 24939 6055 24945
rect 5997 24936 6009 24939
rect 5592 24908 6009 24936
rect 5592 24896 5598 24908
rect 5997 24905 6009 24908
rect 6043 24905 6055 24939
rect 5997 24899 6055 24905
rect 3234 24868 3240 24880
rect 2188 24840 2452 24868
rect 2700 24840 3240 24868
rect 2188 24828 2194 24840
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 1670 24800 1676 24812
rect 1627 24772 1676 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 1670 24760 1676 24772
rect 1728 24760 1734 24812
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24769 2375 24803
rect 2317 24763 2375 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 2700 24800 2728 24840
rect 3234 24828 3240 24840
rect 3292 24828 3298 24880
rect 4700 24871 4758 24877
rect 4700 24837 4712 24871
rect 4746 24868 4758 24871
rect 4798 24868 4804 24880
rect 4746 24840 4804 24868
rect 4746 24837 4758 24840
rect 4700 24831 4758 24837
rect 4798 24828 4804 24840
rect 4856 24828 4862 24880
rect 6012 24868 6040 24899
rect 10778 24896 10784 24948
rect 10836 24896 10842 24948
rect 11330 24896 11336 24948
rect 11388 24896 11394 24948
rect 11422 24896 11428 24948
rect 11480 24936 11486 24948
rect 13357 24939 13415 24945
rect 13357 24936 13369 24939
rect 11480 24908 13369 24936
rect 11480 24896 11486 24908
rect 13357 24905 13369 24908
rect 13403 24905 13415 24939
rect 13357 24899 13415 24905
rect 13814 24896 13820 24948
rect 13872 24936 13878 24948
rect 13872 24908 14412 24936
rect 13872 24896 13878 24908
rect 9953 24871 10011 24877
rect 6012 24840 6684 24868
rect 2639 24772 2728 24800
rect 2777 24803 2835 24809
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 2777 24769 2789 24803
rect 2823 24800 2835 24803
rect 2866 24800 2872 24812
rect 2823 24772 2872 24800
rect 2823 24769 2835 24772
rect 2777 24763 2835 24769
rect 1489 24735 1547 24741
rect 1489 24701 1501 24735
rect 1535 24701 1547 24735
rect 1489 24695 1547 24701
rect 2332 24664 2360 24763
rect 2866 24760 2872 24772
rect 2924 24800 2930 24812
rect 3326 24800 3332 24812
rect 2924 24772 3332 24800
rect 2924 24760 2930 24772
rect 3326 24760 3332 24772
rect 3384 24760 3390 24812
rect 3786 24760 3792 24812
rect 3844 24800 3850 24812
rect 4433 24803 4491 24809
rect 4433 24800 4445 24803
rect 3844 24772 4445 24800
rect 3844 24760 3850 24772
rect 4433 24769 4445 24772
rect 4479 24769 4491 24803
rect 5905 24803 5963 24809
rect 5905 24800 5917 24803
rect 4433 24763 4491 24769
rect 5552 24772 5917 24800
rect 5552 24744 5580 24772
rect 5905 24769 5917 24772
rect 5951 24769 5963 24803
rect 5905 24763 5963 24769
rect 6089 24803 6147 24809
rect 6089 24769 6101 24803
rect 6135 24769 6147 24803
rect 6089 24763 6147 24769
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 3936 24704 4261 24732
rect 3936 24692 3942 24704
rect 4249 24701 4261 24704
rect 4295 24701 4307 24735
rect 4249 24695 4307 24701
rect 5534 24692 5540 24744
rect 5592 24692 5598 24744
rect 6104 24664 6132 24763
rect 6178 24760 6184 24812
rect 6236 24800 6242 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 6236 24772 6561 24800
rect 6236 24760 6242 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6656 24741 6684 24840
rect 9953 24837 9965 24871
rect 9999 24868 10011 24871
rect 11146 24868 11152 24880
rect 9999 24840 11152 24868
rect 9999 24837 10011 24840
rect 9953 24831 10011 24837
rect 11146 24828 11152 24840
rect 11204 24828 11210 24880
rect 11348 24868 11376 24896
rect 11348 24840 11836 24868
rect 7653 24803 7711 24809
rect 7653 24769 7665 24803
rect 7699 24800 7711 24803
rect 7745 24803 7803 24809
rect 7745 24800 7757 24803
rect 7699 24772 7757 24800
rect 7699 24769 7711 24772
rect 7653 24763 7711 24769
rect 7745 24769 7757 24772
rect 7791 24769 7803 24803
rect 7745 24763 7803 24769
rect 7929 24803 7987 24809
rect 7929 24769 7941 24803
rect 7975 24800 7987 24803
rect 8202 24800 8208 24812
rect 7975 24772 8208 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 8202 24760 8208 24772
rect 8260 24760 8266 24812
rect 8294 24760 8300 24812
rect 8352 24760 8358 24812
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 10781 24803 10839 24809
rect 10781 24800 10793 24803
rect 10744 24772 10793 24800
rect 10744 24760 10750 24772
rect 10781 24769 10793 24772
rect 10827 24769 10839 24803
rect 10781 24763 10839 24769
rect 10870 24760 10876 24812
rect 10928 24800 10934 24812
rect 11241 24803 11299 24809
rect 11241 24800 11253 24803
rect 10928 24772 11253 24800
rect 10928 24760 10934 24772
rect 11241 24769 11253 24772
rect 11287 24769 11299 24803
rect 11241 24763 11299 24769
rect 11514 24760 11520 24812
rect 11572 24760 11578 24812
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 11808 24809 11836 24840
rect 13630 24828 13636 24880
rect 13688 24828 13694 24880
rect 14277 24871 14335 24877
rect 14277 24868 14289 24871
rect 14016 24840 14289 24868
rect 11793 24803 11851 24809
rect 11793 24769 11805 24803
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 13354 24760 13360 24812
rect 13412 24760 13418 24812
rect 13538 24760 13544 24812
rect 13596 24760 13602 24812
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24800 13783 24803
rect 13814 24800 13820 24812
rect 13771 24772 13820 24800
rect 13771 24769 13783 24772
rect 13725 24763 13783 24769
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 13906 24760 13912 24812
rect 13964 24760 13970 24812
rect 6641 24735 6699 24741
rect 6641 24701 6653 24735
rect 6687 24701 6699 24735
rect 6641 24695 6699 24701
rect 7009 24735 7067 24741
rect 7009 24701 7021 24735
rect 7055 24701 7067 24735
rect 7009 24695 7067 24701
rect 6822 24664 6828 24676
rect 2332 24636 4476 24664
rect 1118 24556 1124 24608
rect 1176 24596 1182 24608
rect 2133 24599 2191 24605
rect 2133 24596 2145 24599
rect 1176 24568 2145 24596
rect 1176 24556 1182 24568
rect 2133 24565 2145 24568
rect 2179 24565 2191 24599
rect 2133 24559 2191 24565
rect 3694 24556 3700 24608
rect 3752 24556 3758 24608
rect 4448 24596 4476 24636
rect 5460 24636 6040 24664
rect 6104 24636 6828 24664
rect 5460 24596 5488 24636
rect 4448 24568 5488 24596
rect 5534 24556 5540 24608
rect 5592 24596 5598 24608
rect 5813 24599 5871 24605
rect 5813 24596 5825 24599
rect 5592 24568 5825 24596
rect 5592 24556 5598 24568
rect 5813 24565 5825 24568
rect 5859 24565 5871 24599
rect 6012 24596 6040 24636
rect 6822 24624 6828 24636
rect 6880 24624 6886 24676
rect 6917 24667 6975 24673
rect 6917 24633 6929 24667
rect 6963 24664 6975 24667
rect 7024 24664 7052 24695
rect 10042 24692 10048 24744
rect 10100 24692 10106 24744
rect 13372 24732 13400 24760
rect 14016 24732 14044 24840
rect 14277 24837 14289 24840
rect 14323 24837 14335 24871
rect 14277 24831 14335 24837
rect 14384 24809 14412 24908
rect 14458 24896 14464 24948
rect 14516 24936 14522 24948
rect 14829 24939 14887 24945
rect 14829 24936 14841 24939
rect 14516 24908 14841 24936
rect 14516 24896 14522 24908
rect 14829 24905 14841 24908
rect 14875 24905 14887 24939
rect 15378 24936 15384 24948
rect 14829 24899 14887 24905
rect 15120 24908 15384 24936
rect 15120 24868 15148 24908
rect 15378 24896 15384 24908
rect 15436 24936 15442 24948
rect 15746 24936 15752 24948
rect 15436 24908 15752 24936
rect 15436 24896 15442 24908
rect 15746 24896 15752 24908
rect 15804 24896 15810 24948
rect 19058 24936 19064 24948
rect 16960 24908 19064 24936
rect 16960 24877 16988 24908
rect 19058 24896 19064 24908
rect 19116 24896 19122 24948
rect 20162 24896 20168 24948
rect 20220 24896 20226 24948
rect 22189 24939 22247 24945
rect 22189 24905 22201 24939
rect 22235 24936 22247 24939
rect 22554 24936 22560 24948
rect 22235 24908 22560 24936
rect 22235 24905 22247 24908
rect 22189 24899 22247 24905
rect 22554 24896 22560 24908
rect 22612 24896 22618 24948
rect 25682 24896 25688 24948
rect 25740 24936 25746 24948
rect 25961 24939 26019 24945
rect 25961 24936 25973 24939
rect 25740 24908 25973 24936
rect 25740 24896 25746 24908
rect 25961 24905 25973 24908
rect 26007 24905 26019 24939
rect 25961 24899 26019 24905
rect 26418 24896 26424 24948
rect 26476 24896 26482 24948
rect 27249 24939 27307 24945
rect 27249 24905 27261 24939
rect 27295 24936 27307 24939
rect 27522 24936 27528 24948
rect 27295 24908 27528 24936
rect 27295 24905 27307 24908
rect 27249 24899 27307 24905
rect 27522 24896 27528 24908
rect 27580 24936 27586 24948
rect 28442 24936 28448 24948
rect 27580 24908 28448 24936
rect 27580 24896 27586 24908
rect 28442 24896 28448 24908
rect 28500 24896 28506 24948
rect 29546 24896 29552 24948
rect 29604 24936 29610 24948
rect 29641 24939 29699 24945
rect 29641 24936 29653 24939
rect 29604 24908 29653 24936
rect 29604 24896 29610 24908
rect 29641 24905 29653 24908
rect 29687 24905 29699 24939
rect 29641 24899 29699 24905
rect 31202 24896 31208 24948
rect 31260 24896 31266 24948
rect 14936 24840 15148 24868
rect 15197 24871 15255 24877
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24769 14243 24803
rect 14185 24763 14243 24769
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24769 14427 24803
rect 14369 24763 14427 24769
rect 10428 24704 12756 24732
rect 13372 24704 14044 24732
rect 10428 24664 10456 24704
rect 6963 24636 7052 24664
rect 7300 24636 10456 24664
rect 12728 24664 12756 24704
rect 14001 24667 14059 24673
rect 14001 24664 14013 24667
rect 12728 24636 14013 24664
rect 6963 24633 6975 24636
rect 6917 24627 6975 24633
rect 7300 24596 7328 24636
rect 14001 24633 14013 24636
rect 14047 24633 14059 24667
rect 14001 24627 14059 24633
rect 14200 24664 14228 24763
rect 14384 24732 14412 24763
rect 14550 24760 14556 24812
rect 14608 24760 14614 24812
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14936 24809 14964 24840
rect 15197 24837 15209 24871
rect 15243 24868 15255 24871
rect 16945 24871 17003 24877
rect 16945 24868 16957 24871
rect 15243 24840 16957 24868
rect 15243 24837 15255 24840
rect 15197 24831 15255 24837
rect 16945 24837 16957 24840
rect 16991 24837 17003 24871
rect 16945 24831 17003 24837
rect 14921 24803 14979 24809
rect 14921 24769 14933 24803
rect 14967 24769 14979 24803
rect 14921 24763 14979 24769
rect 15013 24803 15071 24809
rect 15013 24769 15025 24803
rect 15059 24800 15071 24803
rect 15102 24800 15108 24812
rect 15059 24772 15108 24800
rect 15059 24769 15071 24772
rect 15013 24763 15071 24769
rect 15102 24760 15108 24772
rect 15160 24760 15166 24812
rect 15212 24732 15240 24831
rect 17034 24828 17040 24880
rect 17092 24828 17098 24880
rect 17144 24840 19288 24868
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15381 24803 15439 24809
rect 15381 24769 15393 24803
rect 15427 24769 15439 24803
rect 15381 24763 15439 24769
rect 14384 24704 15240 24732
rect 15396 24664 15424 24763
rect 16758 24760 16764 24812
rect 16816 24760 16822 24812
rect 17144 24809 17172 24840
rect 17129 24803 17187 24809
rect 17129 24800 17141 24803
rect 17057 24772 17141 24800
rect 17057 24664 17085 24772
rect 17129 24769 17141 24772
rect 17175 24769 17187 24803
rect 17129 24763 17187 24769
rect 18874 24760 18880 24812
rect 18932 24760 18938 24812
rect 19058 24760 19064 24812
rect 19116 24760 19122 24812
rect 19150 24760 19156 24812
rect 19208 24760 19214 24812
rect 19260 24809 19288 24840
rect 20088 24840 21404 24868
rect 20088 24809 20116 24840
rect 21192 24812 21220 24840
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24769 19303 24803
rect 19245 24763 19303 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 19260 24732 19288 24763
rect 20254 24760 20260 24812
rect 20312 24800 20318 24812
rect 20714 24800 20720 24812
rect 20312 24772 20720 24800
rect 20312 24760 20318 24772
rect 20714 24760 20720 24772
rect 20772 24800 20778 24812
rect 20901 24803 20959 24809
rect 20901 24800 20913 24803
rect 20772 24772 20913 24800
rect 20772 24760 20778 24772
rect 20901 24769 20913 24772
rect 20947 24769 20959 24803
rect 20901 24763 20959 24769
rect 21174 24760 21180 24812
rect 21232 24760 21238 24812
rect 21266 24760 21272 24812
rect 21324 24760 21330 24812
rect 21376 24809 21404 24840
rect 21450 24828 21456 24880
rect 21508 24868 21514 24880
rect 22097 24871 22155 24877
rect 22097 24868 22109 24871
rect 21508 24840 22109 24868
rect 21508 24828 21514 24840
rect 22097 24837 22109 24840
rect 22143 24837 22155 24871
rect 22278 24868 22284 24880
rect 22097 24831 22155 24837
rect 22204 24840 22284 24868
rect 21361 24803 21419 24809
rect 21361 24769 21373 24803
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24800 22063 24803
rect 22204 24800 22232 24840
rect 22278 24828 22284 24840
rect 22336 24828 22342 24880
rect 30009 24871 30067 24877
rect 27908 24840 28488 24868
rect 22051 24772 22232 24800
rect 23201 24803 23259 24809
rect 22051 24769 22063 24772
rect 22005 24763 22063 24769
rect 23201 24769 23213 24803
rect 23247 24769 23259 24803
rect 23201 24763 23259 24769
rect 22094 24732 22100 24744
rect 19260 24704 22100 24732
rect 22094 24692 22100 24704
rect 22152 24692 22158 24744
rect 23216 24732 23244 24763
rect 23382 24760 23388 24812
rect 23440 24800 23446 24812
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 23440 24772 25053 24800
rect 23440 24760 23446 24772
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25041 24763 25099 24769
rect 25409 24803 25467 24809
rect 25409 24769 25421 24803
rect 25455 24769 25467 24803
rect 25409 24763 25467 24769
rect 22296 24704 23244 24732
rect 25424 24732 25452 24763
rect 26142 24760 26148 24812
rect 26200 24760 26206 24812
rect 26329 24803 26387 24809
rect 26329 24769 26341 24803
rect 26375 24800 26387 24803
rect 27908 24800 27936 24840
rect 26375 24772 27936 24800
rect 27985 24803 28043 24809
rect 26375 24769 26387 24772
rect 26329 24763 26387 24769
rect 27985 24769 27997 24803
rect 28031 24800 28043 24803
rect 28074 24800 28080 24812
rect 28031 24772 28080 24800
rect 28031 24769 28043 24772
rect 27985 24763 28043 24769
rect 26344 24732 26372 24763
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 28258 24760 28264 24812
rect 28316 24760 28322 24812
rect 28353 24803 28411 24809
rect 28353 24769 28365 24803
rect 28399 24769 28411 24803
rect 28460 24800 28488 24840
rect 30009 24837 30021 24871
rect 30055 24868 30067 24871
rect 30558 24868 30564 24880
rect 30055 24840 30564 24868
rect 30055 24837 30067 24840
rect 30009 24831 30067 24837
rect 30558 24828 30564 24840
rect 30616 24828 30622 24880
rect 28460 24772 28856 24800
rect 28353 24763 28411 24769
rect 25424 24704 26372 24732
rect 14200 24636 17085 24664
rect 6012 24568 7328 24596
rect 5813 24559 5871 24565
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 7745 24599 7803 24605
rect 7745 24596 7757 24599
rect 7432 24568 7757 24596
rect 7432 24556 7438 24568
rect 7745 24565 7757 24568
rect 7791 24565 7803 24599
rect 7745 24559 7803 24565
rect 10686 24556 10692 24608
rect 10744 24556 10750 24608
rect 10962 24556 10968 24608
rect 11020 24556 11026 24608
rect 11054 24556 11060 24608
rect 11112 24605 11118 24608
rect 11112 24599 11161 24605
rect 11112 24565 11115 24599
rect 11149 24565 11161 24599
rect 11112 24559 11161 24565
rect 11112 24556 11118 24559
rect 11238 24556 11244 24608
rect 11296 24596 11302 24608
rect 11517 24599 11575 24605
rect 11517 24596 11529 24599
rect 11296 24568 11529 24596
rect 11296 24556 11302 24568
rect 11517 24565 11529 24568
rect 11563 24565 11575 24599
rect 11517 24559 11575 24565
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 14200 24596 14228 24636
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 22296 24664 22324 24704
rect 19300 24636 22324 24664
rect 22373 24667 22431 24673
rect 19300 24624 19306 24636
rect 22373 24633 22385 24667
rect 22419 24633 22431 24667
rect 22373 24627 22431 24633
rect 13596 24568 14228 24596
rect 13596 24556 13602 24568
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 15565 24599 15623 24605
rect 15565 24596 15577 24599
rect 15528 24568 15577 24596
rect 15528 24556 15534 24568
rect 15565 24565 15577 24568
rect 15611 24565 15623 24599
rect 15565 24559 15623 24565
rect 17218 24556 17224 24608
rect 17276 24596 17282 24608
rect 17313 24599 17371 24605
rect 17313 24596 17325 24599
rect 17276 24568 17325 24596
rect 17276 24556 17282 24568
rect 17313 24565 17325 24568
rect 17359 24565 17371 24599
rect 17313 24559 17371 24565
rect 19429 24599 19487 24605
rect 19429 24565 19441 24599
rect 19475 24596 19487 24599
rect 19610 24596 19616 24608
rect 19475 24568 19616 24596
rect 19475 24565 19487 24568
rect 19429 24559 19487 24565
rect 19610 24556 19616 24568
rect 19668 24556 19674 24608
rect 21361 24599 21419 24605
rect 21361 24565 21373 24599
rect 21407 24596 21419 24599
rect 21450 24596 21456 24608
rect 21407 24568 21456 24596
rect 21407 24565 21419 24568
rect 21361 24559 21419 24565
rect 21450 24556 21456 24568
rect 21508 24556 21514 24608
rect 21542 24556 21548 24608
rect 21600 24556 21606 24608
rect 21818 24556 21824 24608
rect 21876 24556 21882 24608
rect 22002 24556 22008 24608
rect 22060 24596 22066 24608
rect 22388 24596 22416 24627
rect 27154 24624 27160 24676
rect 27212 24664 27218 24676
rect 27212 24636 27752 24664
rect 27212 24624 27218 24636
rect 22060 24568 22416 24596
rect 22060 24556 22066 24568
rect 24302 24556 24308 24608
rect 24360 24596 24366 24608
rect 24489 24599 24547 24605
rect 24489 24596 24501 24599
rect 24360 24568 24501 24596
rect 24360 24556 24366 24568
rect 24489 24565 24501 24568
rect 24535 24596 24547 24599
rect 25130 24596 25136 24608
rect 24535 24568 25136 24596
rect 24535 24565 24547 24568
rect 24489 24559 24547 24565
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 25222 24556 25228 24608
rect 25280 24556 25286 24608
rect 25406 24556 25412 24608
rect 25464 24596 25470 24608
rect 25501 24599 25559 24605
rect 25501 24596 25513 24599
rect 25464 24568 25513 24596
rect 25464 24556 25470 24568
rect 25501 24565 25513 24568
rect 25547 24565 25559 24599
rect 27724 24596 27752 24636
rect 28368 24596 28396 24763
rect 28828 24664 28856 24772
rect 28902 24760 28908 24812
rect 28960 24800 28966 24812
rect 30101 24803 30159 24809
rect 30101 24800 30113 24803
rect 28960 24772 30113 24800
rect 28960 24760 28966 24772
rect 30101 24769 30113 24772
rect 30147 24800 30159 24803
rect 30466 24800 30472 24812
rect 30147 24772 30472 24800
rect 30147 24769 30159 24772
rect 30101 24763 30159 24769
rect 30466 24760 30472 24772
rect 30524 24800 30530 24812
rect 31220 24800 31248 24896
rect 30524 24772 31248 24800
rect 31404 24840 31616 24868
rect 30524 24760 30530 24772
rect 30285 24735 30343 24741
rect 30285 24701 30297 24735
rect 30331 24701 30343 24735
rect 30285 24695 30343 24701
rect 28828 24636 28948 24664
rect 27724 24568 28396 24596
rect 25501 24559 25559 24565
rect 28442 24556 28448 24608
rect 28500 24556 28506 24608
rect 28810 24556 28816 24608
rect 28868 24556 28874 24608
rect 28920 24596 28948 24636
rect 28994 24624 29000 24676
rect 29052 24664 29058 24676
rect 30300 24664 30328 24695
rect 30650 24692 30656 24744
rect 30708 24732 30714 24744
rect 31404 24732 31432 24840
rect 31588 24809 31616 24840
rect 32214 24828 32220 24880
rect 32272 24868 32278 24880
rect 32493 24871 32551 24877
rect 32493 24868 32505 24871
rect 32272 24840 32505 24868
rect 32272 24828 32278 24840
rect 32493 24837 32505 24840
rect 32539 24837 32551 24871
rect 32493 24831 32551 24837
rect 31481 24803 31539 24809
rect 31481 24769 31493 24803
rect 31527 24769 31539 24803
rect 31481 24763 31539 24769
rect 31573 24803 31631 24809
rect 31573 24769 31585 24803
rect 31619 24769 31631 24803
rect 31573 24763 31631 24769
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24800 32643 24803
rect 32631 24772 33180 24800
rect 32631 24769 32643 24772
rect 32585 24763 32643 24769
rect 30708 24704 31432 24732
rect 31496 24732 31524 24763
rect 33152 24744 33180 24772
rect 32677 24735 32735 24741
rect 31496 24704 32168 24732
rect 30708 24692 30714 24704
rect 32140 24673 32168 24704
rect 32677 24701 32689 24735
rect 32723 24701 32735 24735
rect 32677 24695 32735 24701
rect 32125 24667 32183 24673
rect 29052 24636 32076 24664
rect 29052 24624 29058 24636
rect 30650 24596 30656 24608
rect 28920 24568 30656 24596
rect 30650 24556 30656 24568
rect 30708 24556 30714 24608
rect 31110 24556 31116 24608
rect 31168 24596 31174 24608
rect 31297 24599 31355 24605
rect 31297 24596 31309 24599
rect 31168 24568 31309 24596
rect 31168 24556 31174 24568
rect 31297 24565 31309 24568
rect 31343 24565 31355 24599
rect 31297 24559 31355 24565
rect 31662 24556 31668 24608
rect 31720 24556 31726 24608
rect 32048 24596 32076 24636
rect 32125 24633 32137 24667
rect 32171 24633 32183 24667
rect 32125 24627 32183 24633
rect 32692 24596 32720 24695
rect 33134 24692 33140 24744
rect 33192 24692 33198 24744
rect 32048 24568 32720 24596
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 3053 24395 3111 24401
rect 3053 24361 3065 24395
rect 3099 24392 3111 24395
rect 3234 24392 3240 24404
rect 3099 24364 3240 24392
rect 3099 24361 3111 24364
rect 3053 24355 3111 24361
rect 3234 24352 3240 24364
rect 3292 24352 3298 24404
rect 5261 24395 5319 24401
rect 5261 24361 5273 24395
rect 5307 24392 5319 24395
rect 5442 24392 5448 24404
rect 5307 24364 5448 24392
rect 5307 24361 5319 24364
rect 5261 24355 5319 24361
rect 5442 24352 5448 24364
rect 5500 24352 5506 24404
rect 5721 24395 5779 24401
rect 5721 24361 5733 24395
rect 5767 24392 5779 24395
rect 6178 24392 6184 24404
rect 5767 24364 6184 24392
rect 5767 24361 5779 24364
rect 5721 24355 5779 24361
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 5736 24324 5764 24355
rect 6178 24352 6184 24364
rect 6236 24352 6242 24404
rect 7374 24392 7380 24404
rect 7116 24364 7380 24392
rect 4856 24296 5764 24324
rect 4856 24284 4862 24296
rect 3786 24256 3792 24268
rect 2746 24228 3792 24256
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24188 1731 24191
rect 2746 24188 2774 24228
rect 3786 24216 3792 24228
rect 3844 24216 3850 24268
rect 7116 24256 7144 24364
rect 7374 24352 7380 24364
rect 7432 24352 7438 24404
rect 9585 24395 9643 24401
rect 9585 24361 9597 24395
rect 9631 24392 9643 24395
rect 10042 24392 10048 24404
rect 9631 24364 10048 24392
rect 9631 24361 9643 24364
rect 9585 24355 9643 24361
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 18874 24352 18880 24404
rect 18932 24392 18938 24404
rect 19061 24395 19119 24401
rect 19061 24392 19073 24395
rect 18932 24364 19073 24392
rect 18932 24352 18938 24364
rect 19061 24361 19073 24364
rect 19107 24392 19119 24395
rect 19107 24364 19840 24392
rect 19107 24361 19119 24364
rect 19061 24355 19119 24361
rect 12805 24327 12863 24333
rect 12805 24293 12817 24327
rect 12851 24324 12863 24327
rect 13906 24324 13912 24336
rect 12851 24296 13912 24324
rect 12851 24293 12863 24296
rect 12805 24287 12863 24293
rect 13906 24284 13912 24296
rect 13964 24284 13970 24336
rect 5460 24228 5672 24256
rect 1719 24160 2774 24188
rect 3145 24191 3203 24197
rect 1719 24157 1731 24160
rect 1673 24151 1731 24157
rect 3145 24157 3157 24191
rect 3191 24188 3203 24191
rect 3234 24188 3240 24200
rect 3191 24160 3240 24188
rect 3191 24157 3203 24160
rect 3145 24151 3203 24157
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 3326 24148 3332 24200
rect 3384 24188 3390 24200
rect 3421 24191 3479 24197
rect 3421 24188 3433 24191
rect 3384 24160 3433 24188
rect 3384 24148 3390 24160
rect 3421 24157 3433 24160
rect 3467 24157 3479 24191
rect 3421 24151 3479 24157
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24188 3663 24191
rect 3694 24188 3700 24200
rect 3651 24160 3700 24188
rect 3651 24157 3663 24160
rect 3605 24151 3663 24157
rect 1940 24123 1998 24129
rect 1940 24089 1952 24123
rect 1986 24120 1998 24123
rect 2038 24120 2044 24132
rect 1986 24092 2044 24120
rect 1986 24089 1998 24092
rect 1940 24083 1998 24089
rect 2038 24080 2044 24092
rect 2096 24080 2102 24132
rect 3234 24012 3240 24064
rect 3292 24012 3298 24064
rect 3436 24052 3464 24151
rect 3694 24148 3700 24160
rect 3752 24148 3758 24200
rect 5350 24148 5356 24200
rect 5408 24188 5414 24200
rect 5460 24197 5488 24228
rect 5445 24191 5503 24197
rect 5445 24188 5457 24191
rect 5408 24160 5457 24188
rect 5408 24148 5414 24160
rect 5445 24157 5457 24160
rect 5491 24157 5503 24191
rect 5445 24151 5503 24157
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 3513 24123 3571 24129
rect 3513 24089 3525 24123
rect 3559 24120 3571 24123
rect 4034 24123 4092 24129
rect 4034 24120 4046 24123
rect 3559 24092 4046 24120
rect 3559 24089 3571 24092
rect 3513 24083 3571 24089
rect 4034 24089 4046 24092
rect 4080 24089 4092 24123
rect 5552 24120 5580 24148
rect 4034 24083 4092 24089
rect 4724 24092 5580 24120
rect 4724 24064 4752 24092
rect 4154 24052 4160 24064
rect 3436 24024 4160 24052
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 4706 24012 4712 24064
rect 4764 24012 4770 24064
rect 5169 24055 5227 24061
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5442 24052 5448 24064
rect 5215 24024 5448 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 5644 24052 5672 24228
rect 7024 24228 7144 24256
rect 6845 24191 6903 24197
rect 6845 24157 6857 24191
rect 6891 24188 6903 24191
rect 7024 24188 7052 24228
rect 8294 24216 8300 24268
rect 8352 24216 8358 24268
rect 9950 24216 9956 24268
rect 10008 24216 10014 24268
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 17589 24259 17647 24265
rect 13596 24228 14872 24256
rect 13596 24216 13602 24228
rect 6891 24160 7052 24188
rect 7101 24191 7159 24197
rect 6891 24157 6903 24160
rect 6845 24151 6903 24157
rect 7101 24157 7113 24191
rect 7147 24188 7159 24191
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 7147 24160 7205 24188
rect 7147 24157 7159 24160
rect 7101 24151 7159 24157
rect 7193 24157 7205 24160
rect 7239 24188 7251 24191
rect 8312 24188 8340 24216
rect 7239 24160 8340 24188
rect 9968 24188 9996 24216
rect 10965 24191 11023 24197
rect 10965 24188 10977 24191
rect 9968 24160 10977 24188
rect 7239 24157 7251 24160
rect 7193 24151 7251 24157
rect 10965 24157 10977 24160
rect 11011 24188 11023 24191
rect 11054 24188 11060 24200
rect 11011 24160 11060 24188
rect 11011 24157 11023 24160
rect 10965 24151 11023 24157
rect 11054 24148 11060 24160
rect 11112 24148 11118 24200
rect 7460 24123 7518 24129
rect 7460 24089 7472 24123
rect 7506 24120 7518 24123
rect 7650 24120 7656 24132
rect 7506 24092 7656 24120
rect 7506 24089 7518 24092
rect 7460 24083 7518 24089
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 10720 24123 10778 24129
rect 10720 24089 10732 24123
rect 10766 24120 10778 24123
rect 11238 24120 11244 24132
rect 10766 24092 11244 24120
rect 10766 24089 10778 24092
rect 10720 24083 10778 24089
rect 11238 24080 11244 24092
rect 11296 24080 11302 24132
rect 11333 24123 11391 24129
rect 11333 24089 11345 24123
rect 11379 24120 11391 24123
rect 11606 24120 11612 24132
rect 11379 24092 11612 24120
rect 11379 24089 11391 24092
rect 11333 24083 11391 24089
rect 11606 24080 11612 24092
rect 11664 24080 11670 24132
rect 12342 24080 12348 24132
rect 12400 24080 12406 24132
rect 13357 24123 13415 24129
rect 13357 24120 13369 24123
rect 13188 24092 13369 24120
rect 13188 24064 13216 24092
rect 13357 24089 13369 24092
rect 13403 24089 13415 24123
rect 13357 24083 13415 24089
rect 14844 24064 14872 24228
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 17954 24256 17960 24268
rect 17635 24228 17960 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 17954 24216 17960 24228
rect 18012 24216 18018 24268
rect 19812 24265 19840 24364
rect 21818 24352 21824 24404
rect 21876 24352 21882 24404
rect 23017 24395 23075 24401
rect 23017 24361 23029 24395
rect 23063 24392 23075 24395
rect 23382 24392 23388 24404
rect 23063 24364 23388 24392
rect 23063 24361 23075 24364
rect 23017 24355 23075 24361
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24225 19855 24259
rect 19797 24219 19855 24225
rect 17310 24148 17316 24200
rect 17368 24148 17374 24200
rect 21453 24191 21511 24197
rect 21453 24157 21465 24191
rect 21499 24188 21511 24191
rect 21836 24188 21864 24352
rect 21499 24160 21864 24188
rect 21499 24157 21511 24160
rect 21453 24151 21511 24157
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22925 24191 22983 24197
rect 22925 24188 22937 24191
rect 21968 24160 22937 24188
rect 21968 24148 21974 24160
rect 22925 24157 22937 24160
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 23032 24132 23060 24355
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 26142 24352 26148 24404
rect 26200 24392 26206 24404
rect 26605 24395 26663 24401
rect 26605 24392 26617 24395
rect 26200 24364 26617 24392
rect 26200 24352 26206 24364
rect 26605 24361 26617 24364
rect 26651 24361 26663 24395
rect 27154 24392 27160 24404
rect 26605 24355 26663 24361
rect 27080 24364 27160 24392
rect 25130 24216 25136 24268
rect 25188 24256 25194 24268
rect 26970 24256 26976 24268
rect 25188 24228 26976 24256
rect 25188 24216 25194 24228
rect 26970 24216 26976 24228
rect 27028 24216 27034 24268
rect 27080 24265 27108 24364
rect 27154 24352 27160 24364
rect 27212 24392 27218 24404
rect 27617 24395 27675 24401
rect 27617 24392 27629 24395
rect 27212 24364 27629 24392
rect 27212 24352 27218 24364
rect 27617 24361 27629 24364
rect 27663 24361 27675 24395
rect 27617 24355 27675 24361
rect 28994 24352 29000 24404
rect 29052 24352 29058 24404
rect 33594 24352 33600 24404
rect 33652 24392 33658 24404
rect 35342 24392 35348 24404
rect 33652 24364 35348 24392
rect 33652 24352 33658 24364
rect 35342 24352 35348 24364
rect 35400 24352 35406 24404
rect 29012 24324 29040 24352
rect 27264 24296 29040 24324
rect 27264 24268 27292 24296
rect 27065 24259 27123 24265
rect 27065 24225 27077 24259
rect 27111 24225 27123 24259
rect 27065 24219 27123 24225
rect 27246 24216 27252 24268
rect 27304 24216 27310 24268
rect 28562 24259 28620 24265
rect 28562 24225 28574 24259
rect 28608 24256 28620 24259
rect 28810 24256 28816 24268
rect 28608 24228 28816 24256
rect 28608 24225 28620 24228
rect 28562 24219 28620 24225
rect 28810 24216 28816 24228
rect 28868 24216 28874 24268
rect 29454 24256 29460 24268
rect 29012 24228 29460 24256
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24397 24191 24455 24197
rect 24397 24188 24409 24191
rect 24360 24160 24409 24188
rect 24360 24148 24366 24160
rect 24397 24157 24409 24160
rect 24443 24157 24455 24191
rect 24397 24151 24455 24157
rect 27522 24148 27528 24200
rect 27580 24148 27586 24200
rect 28074 24148 28080 24200
rect 28132 24188 28138 24200
rect 28902 24188 28908 24200
rect 28132 24160 28908 24188
rect 28132 24148 28138 24160
rect 28902 24148 28908 24160
rect 28960 24148 28966 24200
rect 29012 24197 29040 24228
rect 29454 24216 29460 24228
rect 29512 24256 29518 24268
rect 29825 24259 29883 24265
rect 29825 24256 29837 24259
rect 29512 24228 29837 24256
rect 29512 24216 29518 24228
rect 29825 24225 29837 24228
rect 29871 24225 29883 24259
rect 29825 24219 29883 24225
rect 30374 24216 30380 24268
rect 30432 24256 30438 24268
rect 30745 24259 30803 24265
rect 30745 24256 30757 24259
rect 30432 24228 30757 24256
rect 30432 24216 30438 24228
rect 30745 24225 30757 24228
rect 30791 24225 30803 24259
rect 30745 24219 30803 24225
rect 31021 24259 31079 24265
rect 31021 24225 31033 24259
rect 31067 24256 31079 24259
rect 31110 24256 31116 24268
rect 31067 24228 31116 24256
rect 31067 24225 31079 24228
rect 31021 24219 31079 24225
rect 31110 24216 31116 24228
rect 31168 24216 31174 24268
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24157 29055 24191
rect 28997 24151 29055 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24188 29975 24191
rect 30466 24188 30472 24200
rect 29963 24160 30472 24188
rect 29963 24157 29975 24160
rect 29917 24151 29975 24157
rect 18874 24120 18880 24132
rect 18814 24092 18880 24120
rect 18874 24080 18880 24092
rect 18932 24080 18938 24132
rect 22649 24123 22707 24129
rect 22649 24089 22661 24123
rect 22695 24120 22707 24123
rect 23014 24120 23020 24132
rect 22695 24092 23020 24120
rect 22695 24089 22707 24092
rect 22649 24083 22707 24089
rect 23014 24080 23020 24092
rect 23072 24080 23078 24132
rect 24670 24080 24676 24132
rect 24728 24080 24734 24132
rect 25406 24080 25412 24132
rect 25464 24080 25470 24132
rect 26973 24123 27031 24129
rect 26973 24089 26985 24123
rect 27019 24120 27031 24123
rect 28166 24120 28172 24132
rect 27019 24092 28172 24120
rect 27019 24089 27031 24092
rect 26973 24083 27031 24089
rect 28166 24080 28172 24092
rect 28224 24080 28230 24132
rect 28445 24123 28503 24129
rect 28445 24120 28457 24123
rect 28276 24092 28457 24120
rect 6822 24052 6828 24064
rect 5644 24024 6828 24052
rect 6822 24012 6828 24024
rect 6880 24012 6886 24064
rect 8570 24012 8576 24064
rect 8628 24012 8634 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 10962 24052 10968 24064
rect 9732 24024 10968 24052
rect 9732 24012 9738 24024
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 12894 24012 12900 24064
rect 12952 24012 12958 24064
rect 13170 24012 13176 24064
rect 13228 24012 13234 24064
rect 13262 24012 13268 24064
rect 13320 24012 13326 24064
rect 14826 24012 14832 24064
rect 14884 24012 14890 24064
rect 19150 24012 19156 24064
rect 19208 24052 19214 24064
rect 19245 24055 19303 24061
rect 19245 24052 19257 24055
rect 19208 24024 19257 24052
rect 19208 24012 19214 24024
rect 19245 24021 19257 24024
rect 19291 24021 19303 24055
rect 19245 24015 19303 24021
rect 20070 24012 20076 24064
rect 20128 24052 20134 24064
rect 21269 24055 21327 24061
rect 21269 24052 21281 24055
rect 20128 24024 21281 24052
rect 20128 24012 20134 24024
rect 21269 24021 21281 24024
rect 21315 24021 21327 24055
rect 21269 24015 21327 24021
rect 22370 24012 22376 24064
rect 22428 24052 22434 24064
rect 22557 24055 22615 24061
rect 22557 24052 22569 24055
rect 22428 24024 22569 24052
rect 22428 24012 22434 24024
rect 22557 24021 22569 24024
rect 22603 24021 22615 24055
rect 22557 24015 22615 24021
rect 26050 24012 26056 24064
rect 26108 24052 26114 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 26108 24024 26157 24052
rect 26108 24012 26114 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 27982 24012 27988 24064
rect 28040 24052 28046 24064
rect 28276 24052 28304 24092
rect 28445 24089 28457 24092
rect 28491 24089 28503 24123
rect 29012 24120 29040 24151
rect 30466 24148 30472 24160
rect 30524 24148 30530 24200
rect 32582 24148 32588 24200
rect 32640 24148 32646 24200
rect 32861 24191 32919 24197
rect 32861 24157 32873 24191
rect 32907 24188 32919 24191
rect 32907 24160 33180 24188
rect 32907 24157 32919 24160
rect 32861 24151 32919 24157
rect 28445 24083 28503 24089
rect 28552 24092 29040 24120
rect 28040 24024 28304 24052
rect 28040 24012 28046 24024
rect 28350 24012 28356 24064
rect 28408 24052 28414 24064
rect 28552 24052 28580 24092
rect 31662 24080 31668 24132
rect 31720 24080 31726 24132
rect 33152 24064 33180 24160
rect 28408 24024 28580 24052
rect 28408 24012 28414 24024
rect 28626 24012 28632 24064
rect 28684 24052 28690 24064
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28684 24024 28733 24052
rect 28684 24012 28690 24024
rect 28721 24021 28733 24024
rect 28767 24021 28779 24055
rect 28721 24015 28779 24021
rect 28902 24012 28908 24064
rect 28960 24012 28966 24064
rect 30282 24012 30288 24064
rect 30340 24012 30346 24064
rect 30466 24012 30472 24064
rect 30524 24052 30530 24064
rect 30650 24052 30656 24064
rect 30524 24024 30656 24052
rect 30524 24012 30530 24024
rect 30650 24012 30656 24024
rect 30708 24012 30714 24064
rect 32493 24055 32551 24061
rect 32493 24021 32505 24055
rect 32539 24052 32551 24055
rect 33134 24052 33140 24064
rect 32539 24024 33140 24052
rect 32539 24021 32551 24024
rect 32493 24015 32551 24021
rect 33134 24012 33140 24024
rect 33192 24012 33198 24064
rect 1104 23962 38824 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 38824 23962
rect 1104 23888 38824 23910
rect 2038 23808 2044 23860
rect 2096 23808 2102 23860
rect 2130 23808 2136 23860
rect 2188 23808 2194 23860
rect 3234 23808 3240 23860
rect 3292 23808 3298 23860
rect 3878 23808 3884 23860
rect 3936 23808 3942 23860
rect 4062 23808 4068 23860
rect 4120 23848 4126 23860
rect 4433 23851 4491 23857
rect 4433 23848 4445 23851
rect 4120 23820 4445 23848
rect 4120 23808 4126 23820
rect 4433 23817 4445 23820
rect 4479 23817 4491 23851
rect 4433 23811 4491 23817
rect 5350 23808 5356 23860
rect 5408 23808 5414 23860
rect 5442 23808 5448 23860
rect 5500 23808 5506 23860
rect 7650 23808 7656 23860
rect 7708 23808 7714 23860
rect 8849 23851 8907 23857
rect 8849 23817 8861 23851
rect 8895 23848 8907 23851
rect 8895 23820 10824 23848
rect 8895 23817 8907 23820
rect 8849 23811 8907 23817
rect 2041 23715 2099 23721
rect 2041 23681 2053 23715
rect 2087 23712 2099 23715
rect 2148 23712 2176 23808
rect 2087 23684 2176 23712
rect 2225 23715 2283 23721
rect 2087 23681 2099 23684
rect 2041 23675 2099 23681
rect 2225 23681 2237 23715
rect 2271 23712 2283 23715
rect 2777 23715 2835 23721
rect 2777 23712 2789 23715
rect 2271 23684 2789 23712
rect 2271 23681 2283 23684
rect 2225 23675 2283 23681
rect 2777 23681 2789 23684
rect 2823 23681 2835 23715
rect 3252 23712 3280 23808
rect 5169 23783 5227 23789
rect 5169 23780 5181 23783
rect 3804 23752 5181 23780
rect 3804 23721 3832 23752
rect 4908 23721 4936 23752
rect 5169 23749 5181 23752
rect 5215 23749 5227 23783
rect 5169 23743 5227 23749
rect 3329 23715 3387 23721
rect 3329 23712 3341 23715
rect 3252 23684 3341 23712
rect 2777 23675 2835 23681
rect 3329 23681 3341 23684
rect 3375 23681 3387 23715
rect 3329 23675 3387 23681
rect 3789 23715 3847 23721
rect 3789 23681 3801 23715
rect 3835 23681 3847 23715
rect 3789 23675 3847 23681
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23681 4307 23715
rect 4908 23715 4988 23721
rect 4908 23684 4942 23715
rect 4249 23675 4307 23681
rect 4930 23681 4942 23684
rect 4976 23681 4988 23715
rect 4930 23675 4988 23681
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5368 23712 5396 23808
rect 5123 23684 5396 23712
rect 5460 23712 5488 23808
rect 6822 23740 6828 23792
rect 6880 23780 6886 23792
rect 8864 23780 8892 23811
rect 10686 23780 10692 23792
rect 6880 23752 8892 23780
rect 9361 23752 10692 23780
rect 6880 23740 6886 23752
rect 5721 23715 5779 23721
rect 5721 23712 5733 23715
rect 5460 23684 5733 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5721 23681 5733 23684
rect 5767 23681 5779 23715
rect 5721 23675 5779 23681
rect 4264 23644 4292 23675
rect 4706 23644 4712 23656
rect 4264 23616 4712 23644
rect 4706 23604 4712 23616
rect 4764 23604 4770 23656
rect 4111 23579 4169 23585
rect 4111 23545 4123 23579
rect 4157 23576 4169 23579
rect 4798 23576 4804 23588
rect 4157 23548 4804 23576
rect 4157 23545 4169 23548
rect 4111 23539 4169 23545
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 3973 23511 4031 23517
rect 3973 23477 3985 23511
rect 4019 23508 4031 23511
rect 5092 23508 5120 23675
rect 7834 23672 7840 23724
rect 7892 23672 7898 23724
rect 8018 23672 8024 23724
rect 8076 23712 8082 23724
rect 8113 23715 8171 23721
rect 8113 23712 8125 23715
rect 8076 23684 8125 23712
rect 8076 23672 8082 23684
rect 8113 23681 8125 23684
rect 8159 23681 8171 23715
rect 8113 23675 8171 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23712 8539 23715
rect 9214 23712 9220 23724
rect 8527 23684 9220 23712
rect 8527 23681 8539 23684
rect 8481 23675 8539 23681
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 8570 23604 8576 23656
rect 8628 23644 8634 23656
rect 8665 23647 8723 23653
rect 8665 23644 8677 23647
rect 8628 23616 8677 23644
rect 8628 23604 8634 23616
rect 8665 23613 8677 23616
rect 8711 23644 8723 23647
rect 9030 23644 9036 23656
rect 8711 23616 9036 23644
rect 8711 23613 8723 23616
rect 8665 23607 8723 23613
rect 9030 23604 9036 23616
rect 9088 23644 9094 23656
rect 9127 23647 9185 23653
rect 9127 23644 9139 23647
rect 9088 23616 9139 23644
rect 9088 23604 9094 23616
rect 9127 23613 9139 23616
rect 9173 23613 9185 23647
rect 9127 23607 9185 23613
rect 9361 23585 9389 23752
rect 10686 23740 10692 23752
rect 10744 23740 10750 23792
rect 10796 23780 10824 23820
rect 11606 23808 11612 23860
rect 11664 23808 11670 23860
rect 11698 23808 11704 23860
rect 11756 23808 11762 23860
rect 12342 23808 12348 23860
rect 12400 23808 12406 23860
rect 12894 23808 12900 23860
rect 12952 23808 12958 23860
rect 13081 23851 13139 23857
rect 13081 23817 13093 23851
rect 13127 23848 13139 23851
rect 13262 23848 13268 23860
rect 13127 23820 13268 23848
rect 13127 23817 13139 23820
rect 13081 23811 13139 23817
rect 13262 23808 13268 23820
rect 13320 23808 13326 23860
rect 13906 23808 13912 23860
rect 13964 23808 13970 23860
rect 14185 23851 14243 23857
rect 14185 23817 14197 23851
rect 14231 23817 14243 23851
rect 14185 23811 14243 23817
rect 16669 23851 16727 23857
rect 16669 23817 16681 23851
rect 16715 23817 16727 23851
rect 16669 23811 16727 23817
rect 11716 23780 11744 23808
rect 12912 23780 12940 23808
rect 10796 23752 11744 23780
rect 11808 23752 12940 23780
rect 9490 23672 9496 23724
rect 9548 23712 9554 23724
rect 9585 23715 9643 23721
rect 9585 23712 9597 23715
rect 9548 23684 9597 23712
rect 9548 23672 9554 23684
rect 9585 23681 9597 23684
rect 9631 23712 9643 23715
rect 9674 23712 9680 23724
rect 9631 23684 9680 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 9674 23672 9680 23684
rect 9732 23672 9738 23724
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23712 9827 23715
rect 10870 23712 10876 23724
rect 9815 23684 10876 23712
rect 9815 23681 9827 23684
rect 9769 23675 9827 23681
rect 9784 23644 9812 23675
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 11808 23721 11836 23752
rect 11793 23715 11851 23721
rect 11793 23681 11805 23715
rect 11839 23681 11851 23715
rect 11793 23675 11851 23681
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 12526 23712 12532 23724
rect 12483 23684 12532 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23712 13783 23715
rect 13924 23712 13952 23808
rect 13771 23684 13952 23712
rect 14093 23715 14151 23721
rect 13771 23681 13783 23684
rect 13725 23675 13783 23681
rect 14093 23681 14105 23715
rect 14139 23712 14151 23715
rect 14200 23712 14228 23811
rect 14139 23684 14228 23712
rect 14553 23715 14611 23721
rect 14139 23681 14151 23684
rect 14093 23675 14151 23681
rect 14553 23681 14565 23715
rect 14599 23712 14611 23715
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 14599 23684 15025 23712
rect 14599 23681 14611 23684
rect 14553 23675 14611 23681
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15565 23715 15623 23721
rect 15565 23712 15577 23715
rect 15252 23684 15577 23712
rect 15252 23672 15258 23684
rect 15565 23681 15577 23684
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 16025 23715 16083 23721
rect 16025 23681 16037 23715
rect 16071 23712 16083 23715
rect 16684 23712 16712 23811
rect 17126 23808 17132 23860
rect 17184 23808 17190 23860
rect 18601 23851 18659 23857
rect 18601 23817 18613 23851
rect 18647 23848 18659 23851
rect 19150 23848 19156 23860
rect 18647 23820 19156 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 19150 23808 19156 23820
rect 19208 23808 19214 23860
rect 21542 23808 21548 23860
rect 21600 23808 21606 23860
rect 23477 23851 23535 23857
rect 23477 23817 23489 23851
rect 23523 23848 23535 23851
rect 23750 23848 23756 23860
rect 23523 23820 23756 23848
rect 23523 23817 23535 23820
rect 23477 23811 23535 23817
rect 23750 23808 23756 23820
rect 23808 23808 23814 23860
rect 24670 23808 24676 23860
rect 24728 23808 24734 23860
rect 26053 23851 26111 23857
rect 26053 23817 26065 23851
rect 26099 23817 26111 23851
rect 26053 23811 26111 23817
rect 28629 23851 28687 23857
rect 28629 23817 28641 23851
rect 28675 23848 28687 23851
rect 28810 23848 28816 23860
rect 28675 23820 28816 23848
rect 28675 23817 28687 23820
rect 28629 23811 28687 23817
rect 18874 23740 18880 23792
rect 18932 23740 18938 23792
rect 18966 23740 18972 23792
rect 19024 23780 19030 23792
rect 21453 23783 21511 23789
rect 19024 23752 19288 23780
rect 19024 23740 19030 23752
rect 16071 23684 16712 23712
rect 17037 23715 17095 23721
rect 16071 23681 16083 23684
rect 16025 23675 16083 23681
rect 17037 23681 17049 23715
rect 17083 23712 17095 23715
rect 17497 23715 17555 23721
rect 17497 23712 17509 23715
rect 17083 23684 17509 23712
rect 17083 23681 17095 23684
rect 17037 23675 17095 23681
rect 17497 23681 17509 23684
rect 17543 23681 17555 23715
rect 18892 23712 18920 23740
rect 19260 23721 19288 23752
rect 21453 23749 21465 23783
rect 21499 23780 21511 23783
rect 21560 23780 21588 23808
rect 21499 23752 21588 23780
rect 22480 23752 23612 23780
rect 21499 23749 21511 23752
rect 21453 23743 21511 23749
rect 19153 23715 19211 23721
rect 19153 23712 19165 23715
rect 17497 23675 17555 23681
rect 17604 23684 18828 23712
rect 18892 23684 19165 23712
rect 9508 23616 9812 23644
rect 14645 23647 14703 23653
rect 9508 23588 9536 23616
rect 14645 23613 14657 23647
rect 14691 23613 14703 23647
rect 14645 23607 14703 23613
rect 9346 23579 9404 23585
rect 9346 23545 9358 23579
rect 9392 23545 9404 23579
rect 9346 23539 9404 23545
rect 9490 23536 9496 23588
rect 9548 23536 9554 23588
rect 9582 23536 9588 23588
rect 9640 23536 9646 23588
rect 9858 23536 9864 23588
rect 9916 23536 9922 23588
rect 14660 23576 14688 23607
rect 14826 23604 14832 23656
rect 14884 23644 14890 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 14884 23616 17325 23644
rect 14884 23604 14890 23616
rect 17313 23613 17325 23616
rect 17359 23644 17371 23647
rect 17604 23644 17632 23684
rect 17359 23616 17632 23644
rect 18049 23647 18107 23653
rect 17359 23613 17371 23616
rect 17313 23607 17371 23613
rect 18049 23613 18061 23647
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 14734 23576 14740 23588
rect 14660 23548 14740 23576
rect 14734 23536 14740 23548
rect 14792 23576 14798 23588
rect 15010 23576 15016 23588
rect 14792 23548 15016 23576
rect 14792 23536 14798 23548
rect 15010 23536 15016 23548
rect 15068 23536 15074 23588
rect 16758 23536 16764 23588
rect 16816 23576 16822 23588
rect 18064 23576 18092 23607
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 18693 23647 18751 23653
rect 18693 23644 18705 23647
rect 18472 23616 18705 23644
rect 18472 23604 18478 23616
rect 18693 23613 18705 23616
rect 18739 23613 18751 23647
rect 18800 23644 18828 23684
rect 19153 23681 19165 23684
rect 19199 23681 19211 23715
rect 19153 23675 19211 23681
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 18877 23647 18935 23653
rect 18877 23644 18889 23647
rect 18800 23616 18889 23644
rect 18693 23607 18751 23613
rect 18877 23613 18889 23616
rect 18923 23644 18935 23647
rect 20070 23644 20076 23656
rect 18923 23616 20076 23644
rect 18923 23613 18935 23616
rect 18877 23607 18935 23613
rect 16816 23548 18092 23576
rect 18708 23576 18736 23607
rect 20070 23604 20076 23616
rect 20128 23604 20134 23656
rect 22370 23604 22376 23656
rect 22428 23644 22434 23656
rect 22480 23653 22508 23752
rect 22646 23672 22652 23724
rect 22704 23712 22710 23724
rect 23584 23721 23612 23752
rect 22741 23715 22799 23721
rect 22741 23712 22753 23715
rect 22704 23684 22753 23712
rect 22704 23672 22710 23684
rect 22741 23681 22753 23684
rect 22787 23681 22799 23715
rect 22741 23675 22799 23681
rect 23569 23715 23627 23721
rect 23569 23681 23581 23715
rect 23615 23681 23627 23715
rect 23768 23712 23796 23808
rect 26068 23780 26096 23811
rect 28810 23808 28816 23820
rect 28868 23808 28874 23860
rect 28902 23808 28908 23860
rect 28960 23808 28966 23860
rect 30282 23808 30288 23860
rect 30340 23808 30346 23860
rect 32582 23808 32588 23860
rect 32640 23848 32646 23860
rect 32640 23820 34100 23848
rect 32640 23808 32646 23820
rect 28920 23780 28948 23808
rect 24872 23752 26096 23780
rect 28276 23752 28948 23780
rect 30300 23780 30328 23808
rect 32309 23783 32367 23789
rect 30300 23752 30788 23780
rect 24872 23721 24900 23752
rect 23845 23715 23903 23721
rect 23845 23712 23857 23715
rect 23768 23684 23857 23712
rect 23569 23675 23627 23681
rect 23845 23681 23857 23684
rect 23891 23681 23903 23715
rect 23845 23675 23903 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23712 25007 23715
rect 25130 23712 25136 23724
rect 24995 23684 25136 23712
rect 24995 23681 25007 23684
rect 24949 23675 25007 23681
rect 25130 23672 25136 23684
rect 25188 23672 25194 23724
rect 25225 23715 25283 23721
rect 25225 23681 25237 23715
rect 25271 23712 25283 23715
rect 25271 23684 26096 23712
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 26068 23656 26096 23684
rect 26418 23672 26424 23724
rect 26476 23672 26482 23724
rect 28074 23672 28080 23724
rect 28132 23672 28138 23724
rect 28276 23721 28304 23752
rect 28261 23715 28319 23721
rect 28261 23681 28273 23715
rect 28307 23681 28319 23715
rect 28632 23715 28690 23721
rect 28632 23712 28644 23715
rect 28261 23675 28319 23681
rect 28368 23684 28644 23712
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22428 23616 22477 23644
rect 22428 23604 22434 23616
rect 22465 23613 22477 23616
rect 22511 23613 22523 23647
rect 22465 23607 22523 23613
rect 26050 23604 26056 23656
rect 26108 23644 26114 23656
rect 26513 23647 26571 23653
rect 26513 23644 26525 23647
rect 26108 23616 26525 23644
rect 26108 23604 26114 23616
rect 26513 23613 26525 23616
rect 26559 23613 26571 23647
rect 26513 23607 26571 23613
rect 26697 23647 26755 23653
rect 26697 23613 26709 23647
rect 26743 23644 26755 23647
rect 27246 23644 27252 23656
rect 26743 23616 27252 23644
rect 26743 23613 26755 23616
rect 26697 23607 26755 23613
rect 27246 23604 27252 23616
rect 27304 23604 27310 23656
rect 28092 23644 28120 23672
rect 28169 23647 28227 23653
rect 28169 23644 28181 23647
rect 28092 23616 28181 23644
rect 28169 23613 28181 23616
rect 28215 23613 28227 23647
rect 28169 23607 28227 23613
rect 18708 23548 19104 23576
rect 16816 23536 16822 23548
rect 4019 23480 5120 23508
rect 8021 23511 8079 23517
rect 4019 23477 4031 23480
rect 3973 23471 4031 23477
rect 8021 23477 8033 23511
rect 8067 23508 8079 23511
rect 8297 23511 8355 23517
rect 8297 23508 8309 23511
rect 8067 23480 8309 23508
rect 8067 23477 8079 23480
rect 8021 23471 8079 23477
rect 8297 23477 8309 23480
rect 8343 23477 8355 23511
rect 8297 23471 8355 23477
rect 9217 23511 9275 23517
rect 9217 23477 9229 23511
rect 9263 23508 9275 23511
rect 9876 23508 9904 23536
rect 19076 23520 19104 23548
rect 25866 23536 25872 23588
rect 25924 23576 25930 23588
rect 25924 23548 26372 23576
rect 25924 23536 25930 23548
rect 9263 23480 9904 23508
rect 9263 23477 9275 23480
rect 9217 23471 9275 23477
rect 13906 23468 13912 23520
rect 13964 23468 13970 23520
rect 15746 23468 15752 23520
rect 15804 23508 15810 23520
rect 15841 23511 15899 23517
rect 15841 23508 15853 23511
rect 15804 23480 15853 23508
rect 15804 23468 15810 23480
rect 15841 23477 15853 23480
rect 15887 23477 15899 23511
rect 15841 23471 15899 23477
rect 18230 23468 18236 23520
rect 18288 23468 18294 23520
rect 19058 23468 19064 23520
rect 19116 23468 19122 23520
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 20622 23468 20628 23520
rect 20680 23508 20686 23520
rect 21177 23511 21235 23517
rect 21177 23508 21189 23511
rect 20680 23480 21189 23508
rect 20680 23468 20686 23480
rect 21177 23477 21189 23480
rect 21223 23477 21235 23511
rect 21177 23471 21235 23477
rect 24578 23468 24584 23520
rect 24636 23468 24642 23520
rect 25961 23511 26019 23517
rect 25961 23477 25973 23511
rect 26007 23508 26019 23511
rect 26142 23508 26148 23520
rect 26007 23480 26148 23508
rect 26007 23477 26019 23480
rect 25961 23471 26019 23477
rect 26142 23468 26148 23480
rect 26200 23468 26206 23520
rect 26344 23508 26372 23548
rect 27982 23536 27988 23588
rect 28040 23576 28046 23588
rect 28368 23576 28396 23684
rect 28632 23681 28644 23684
rect 28678 23681 28690 23715
rect 30300 23712 30328 23752
rect 30760 23721 30788 23752
rect 32309 23749 32321 23783
rect 32355 23780 32367 23783
rect 33134 23780 33140 23792
rect 32355 23752 33140 23780
rect 32355 23749 32367 23752
rect 32309 23743 32367 23749
rect 33134 23740 33140 23752
rect 33192 23740 33198 23792
rect 30469 23715 30527 23721
rect 30469 23712 30481 23715
rect 30300 23684 30481 23712
rect 28632 23675 28690 23681
rect 30469 23681 30481 23684
rect 30515 23681 30527 23715
rect 30469 23675 30527 23681
rect 30653 23715 30711 23721
rect 30653 23681 30665 23715
rect 30699 23681 30711 23715
rect 30653 23675 30711 23681
rect 30745 23715 30803 23721
rect 30745 23681 30757 23715
rect 30791 23681 30803 23715
rect 30745 23675 30803 23681
rect 30929 23715 30987 23721
rect 30929 23681 30941 23715
rect 30975 23712 30987 23715
rect 30975 23684 32812 23712
rect 30975 23681 30987 23684
rect 30929 23675 30987 23681
rect 30668 23644 30696 23675
rect 30944 23644 30972 23675
rect 30668 23616 30972 23644
rect 32582 23576 32588 23588
rect 28040 23548 28396 23576
rect 28460 23548 32588 23576
rect 28040 23536 28046 23548
rect 28460 23508 28488 23548
rect 32582 23536 32588 23548
rect 32640 23536 32646 23588
rect 32784 23585 32812 23684
rect 33594 23672 33600 23724
rect 33652 23672 33658 23724
rect 33686 23672 33692 23724
rect 33744 23712 33750 23724
rect 33965 23715 34023 23721
rect 33965 23712 33977 23715
rect 33744 23684 33977 23712
rect 33744 23672 33750 23684
rect 33965 23681 33977 23684
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 33873 23647 33931 23653
rect 33873 23613 33885 23647
rect 33919 23644 33931 23647
rect 34072 23644 34100 23820
rect 34149 23715 34207 23721
rect 34149 23681 34161 23715
rect 34195 23681 34207 23715
rect 34149 23675 34207 23681
rect 33919 23616 34100 23644
rect 33919 23613 33931 23616
rect 33873 23607 33931 23613
rect 32677 23579 32735 23585
rect 32677 23545 32689 23579
rect 32723 23545 32735 23579
rect 32677 23539 32735 23545
rect 32769 23579 32827 23585
rect 32769 23545 32781 23579
rect 32815 23576 32827 23579
rect 34164 23576 34192 23675
rect 32815 23548 32996 23576
rect 32815 23545 32827 23548
rect 32769 23539 32827 23545
rect 26344 23480 28488 23508
rect 28810 23468 28816 23520
rect 28868 23468 28874 23520
rect 30650 23468 30656 23520
rect 30708 23468 30714 23520
rect 30834 23468 30840 23520
rect 30892 23468 30898 23520
rect 32692 23508 32720 23539
rect 32858 23508 32864 23520
rect 32692 23480 32864 23508
rect 32858 23468 32864 23480
rect 32916 23468 32922 23520
rect 32968 23508 32996 23548
rect 33796 23548 34192 23576
rect 33796 23508 33824 23548
rect 32968 23480 33824 23508
rect 33870 23468 33876 23520
rect 33928 23508 33934 23520
rect 33965 23511 34023 23517
rect 33965 23508 33977 23511
rect 33928 23480 33977 23508
rect 33928 23468 33934 23480
rect 33965 23477 33977 23480
rect 34011 23477 34023 23511
rect 33965 23471 34023 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 8018 23264 8024 23316
rect 8076 23304 8082 23316
rect 9582 23304 9588 23316
rect 8076 23276 9588 23304
rect 8076 23264 8082 23276
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 9674 23264 9680 23316
rect 9732 23264 9738 23316
rect 16758 23264 16764 23316
rect 16816 23304 16822 23316
rect 17129 23307 17187 23313
rect 17129 23304 17141 23307
rect 16816 23276 17141 23304
rect 16816 23264 16822 23276
rect 17129 23273 17141 23276
rect 17175 23273 17187 23307
rect 17129 23267 17187 23273
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 18233 23307 18291 23313
rect 18233 23304 18245 23307
rect 18012 23276 18245 23304
rect 18012 23264 18018 23276
rect 18233 23273 18245 23276
rect 18279 23273 18291 23307
rect 18233 23267 18291 23273
rect 21174 23264 21180 23316
rect 21232 23264 21238 23316
rect 25222 23304 25228 23316
rect 25056 23276 25228 23304
rect 2961 23171 3019 23177
rect 2961 23137 2973 23171
rect 3007 23168 3019 23171
rect 3881 23171 3939 23177
rect 3881 23168 3893 23171
rect 3007 23140 3893 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3881 23137 3893 23140
rect 3927 23137 3939 23171
rect 9692 23168 9720 23264
rect 12161 23239 12219 23245
rect 12161 23205 12173 23239
rect 12207 23205 12219 23239
rect 12161 23199 12219 23205
rect 9692 23140 9996 23168
rect 3881 23131 3939 23137
rect 2866 23060 2872 23112
rect 2924 23060 2930 23112
rect 4522 23060 4528 23112
rect 4580 23060 4586 23112
rect 6362 23060 6368 23112
rect 6420 23060 6426 23112
rect 9030 23060 9036 23112
rect 9088 23060 9094 23112
rect 9968 23109 9996 23140
rect 9677 23103 9735 23109
rect 9677 23069 9689 23103
rect 9723 23100 9735 23103
rect 9769 23103 9827 23109
rect 9769 23100 9781 23103
rect 9723 23072 9781 23100
rect 9723 23069 9735 23072
rect 9677 23063 9735 23069
rect 9769 23069 9781 23072
rect 9815 23069 9827 23103
rect 9769 23063 9827 23069
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23069 10011 23103
rect 9953 23063 10011 23069
rect 11885 23103 11943 23109
rect 11885 23069 11897 23103
rect 11931 23100 11943 23103
rect 12176 23100 12204 23199
rect 12526 23128 12532 23180
rect 12584 23128 12590 23180
rect 12805 23171 12863 23177
rect 12805 23137 12817 23171
rect 12851 23168 12863 23171
rect 13538 23168 13544 23180
rect 12851 23140 13544 23168
rect 12851 23137 12863 23140
rect 12805 23131 12863 23137
rect 13538 23128 13544 23140
rect 13596 23128 13602 23180
rect 13633 23171 13691 23177
rect 13633 23137 13645 23171
rect 13679 23168 13691 23171
rect 13814 23168 13820 23180
rect 13679 23140 13820 23168
rect 13679 23137 13691 23140
rect 13633 23131 13691 23137
rect 13814 23128 13820 23140
rect 13872 23168 13878 23180
rect 14550 23168 14556 23180
rect 13872 23140 14556 23168
rect 13872 23128 13878 23140
rect 14550 23128 14556 23140
rect 14608 23128 14614 23180
rect 15381 23171 15439 23177
rect 15381 23137 15393 23171
rect 15427 23168 15439 23171
rect 17310 23168 17316 23180
rect 15427 23140 17316 23168
rect 15427 23137 15439 23140
rect 15381 23131 15439 23137
rect 17310 23128 17316 23140
rect 17368 23168 17374 23180
rect 19426 23168 19432 23180
rect 17368 23140 19432 23168
rect 17368 23128 17374 23140
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 19705 23171 19763 23177
rect 19705 23137 19717 23171
rect 19751 23168 19763 23171
rect 19794 23168 19800 23180
rect 19751 23140 19800 23168
rect 19751 23137 19763 23140
rect 19705 23131 19763 23137
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 24302 23168 24308 23180
rect 21560 23140 24308 23168
rect 11931 23072 12204 23100
rect 12544 23100 12572 23128
rect 21560 23112 21588 23140
rect 24302 23128 24308 23140
rect 24360 23128 24366 23180
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 12544 23072 14381 23100
rect 11931 23069 11943 23072
rect 11885 23063 11943 23069
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 17405 23103 17463 23109
rect 17405 23069 17417 23103
rect 17451 23069 17463 23103
rect 17405 23063 17463 23069
rect 12529 23035 12587 23041
rect 12529 23001 12541 23035
rect 12575 23032 12587 23035
rect 12989 23035 13047 23041
rect 12989 23032 13001 23035
rect 12575 23004 13001 23032
rect 12575 23001 12587 23004
rect 12529 22995 12587 23001
rect 12989 23001 13001 23004
rect 13035 23001 13047 23035
rect 14384 23032 14412 23063
rect 15657 23035 15715 23041
rect 14384 23004 15608 23032
rect 12989 22995 13047 23001
rect 3237 22967 3295 22973
rect 3237 22933 3249 22967
rect 3283 22964 3295 22967
rect 3602 22964 3608 22976
rect 3283 22936 3608 22964
rect 3283 22933 3295 22936
rect 3237 22927 3295 22933
rect 3602 22924 3608 22936
rect 3660 22924 3666 22976
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7190 22964 7196 22976
rect 6963 22936 7196 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7190 22924 7196 22936
rect 7248 22924 7254 22976
rect 9858 22924 9864 22976
rect 9916 22924 9922 22976
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22964 11759 22967
rect 11790 22964 11796 22976
rect 11747 22936 11796 22964
rect 11747 22933 11759 22936
rect 11701 22927 11759 22933
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 12618 22924 12624 22976
rect 12676 22924 12682 22976
rect 14458 22924 14464 22976
rect 14516 22924 14522 22976
rect 15580 22964 15608 23004
rect 15657 23001 15669 23035
rect 15703 23032 15715 23035
rect 15746 23032 15752 23044
rect 15703 23004 15752 23032
rect 15703 23001 15715 23004
rect 15657 22995 15715 23001
rect 15746 22992 15752 23004
rect 15804 22992 15810 23044
rect 17313 23035 17371 23041
rect 17313 23032 17325 23035
rect 16882 23004 17325 23032
rect 17313 23001 17325 23004
rect 17359 23001 17371 23035
rect 17313 22995 17371 23001
rect 17420 23032 17448 23063
rect 18138 23060 18144 23112
rect 18196 23060 18202 23112
rect 18230 23060 18236 23112
rect 18288 23100 18294 23112
rect 18417 23103 18475 23109
rect 18417 23100 18429 23103
rect 18288 23072 18429 23100
rect 18288 23060 18294 23072
rect 18417 23069 18429 23072
rect 18463 23069 18475 23103
rect 18417 23063 18475 23069
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 18966 23100 18972 23112
rect 18555 23072 18972 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 18524 23032 18552 23063
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 21453 23103 21511 23109
rect 21453 23069 21465 23103
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 17420 23004 18552 23032
rect 17420 22964 17448 23004
rect 15580 22936 17448 22964
rect 17954 22924 17960 22976
rect 18012 22924 18018 22976
rect 18598 22924 18604 22976
rect 18656 22924 18662 22976
rect 18984 22964 19012 23060
rect 21361 23035 21419 23041
rect 21361 23032 21373 23035
rect 20930 23004 21373 23032
rect 21361 23001 21373 23004
rect 21407 23001 21419 23035
rect 21361 22995 21419 23001
rect 21468 22976 21496 23063
rect 21542 23060 21548 23112
rect 21600 23060 21606 23112
rect 25056 23109 25084 23276
rect 25222 23264 25228 23276
rect 25280 23304 25286 23316
rect 25866 23304 25872 23316
rect 25280 23276 25872 23304
rect 25280 23264 25286 23276
rect 25866 23264 25872 23276
rect 25924 23264 25930 23316
rect 27522 23264 27528 23316
rect 27580 23304 27586 23316
rect 27893 23307 27951 23313
rect 27893 23304 27905 23307
rect 27580 23276 27905 23304
rect 27580 23264 27586 23276
rect 27893 23273 27905 23276
rect 27939 23273 27951 23307
rect 27893 23267 27951 23273
rect 28166 23264 28172 23316
rect 28224 23304 28230 23316
rect 28261 23307 28319 23313
rect 28261 23304 28273 23307
rect 28224 23276 28273 23304
rect 28224 23264 28230 23276
rect 28261 23273 28273 23276
rect 28307 23273 28319 23307
rect 35434 23304 35440 23316
rect 28261 23267 28319 23273
rect 31726 23276 35440 23304
rect 26142 23196 26148 23248
rect 26200 23236 26206 23248
rect 31726 23236 31754 23276
rect 35434 23264 35440 23276
rect 35492 23264 35498 23316
rect 26200 23208 31754 23236
rect 26200 23196 26206 23208
rect 33134 23196 33140 23248
rect 33192 23196 33198 23248
rect 33321 23239 33379 23245
rect 33321 23205 33333 23239
rect 33367 23236 33379 23239
rect 33686 23236 33692 23248
rect 33367 23208 33692 23236
rect 33367 23205 33379 23208
rect 33321 23199 33379 23205
rect 33686 23196 33692 23208
rect 33744 23196 33750 23248
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23069 25099 23103
rect 25501 23103 25559 23109
rect 25501 23100 25513 23103
rect 25041 23063 25099 23069
rect 25240 23072 25513 23100
rect 21821 23035 21879 23041
rect 21821 23001 21833 23035
rect 21867 23032 21879 23035
rect 22094 23032 22100 23044
rect 21867 23004 22100 23032
rect 21867 23001 21879 23004
rect 21821 22995 21879 23001
rect 22094 22992 22100 23004
rect 22152 22992 22158 23044
rect 22278 22992 22284 23044
rect 22336 22992 22342 23044
rect 23382 22992 23388 23044
rect 23440 23032 23446 23044
rect 23569 23035 23627 23041
rect 23569 23032 23581 23035
rect 23440 23004 23581 23032
rect 23440 22992 23446 23004
rect 23569 23001 23581 23004
rect 23615 23001 23627 23035
rect 23569 22995 23627 23001
rect 25240 22976 25268 23072
rect 25501 23069 25513 23072
rect 25547 23069 25559 23103
rect 25501 23063 25559 23069
rect 25777 23103 25835 23109
rect 25777 23069 25789 23103
rect 25823 23100 25835 23103
rect 26160 23100 26188 23196
rect 25823 23072 26188 23100
rect 27264 23140 28120 23168
rect 25823 23069 25835 23072
rect 25777 23063 25835 23069
rect 27264 23032 27292 23140
rect 27341 23103 27399 23109
rect 27341 23069 27353 23103
rect 27387 23100 27399 23103
rect 27522 23100 27528 23112
rect 27387 23072 27528 23100
rect 27387 23069 27399 23072
rect 27341 23063 27399 23069
rect 27522 23060 27528 23072
rect 27580 23060 27586 23112
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 27663 23072 27920 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 27264 23004 27568 23032
rect 21450 22964 21456 22976
rect 18984 22936 21456 22964
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 25222 22924 25228 22976
rect 25280 22924 25286 22976
rect 26510 22924 26516 22976
rect 26568 22924 26574 22976
rect 27430 22924 27436 22976
rect 27488 22973 27494 22976
rect 27540 22973 27568 23004
rect 27488 22927 27497 22973
rect 27525 22967 27583 22973
rect 27525 22933 27537 22967
rect 27571 22933 27583 22967
rect 27525 22927 27583 22933
rect 27488 22924 27494 22927
rect 27614 22924 27620 22976
rect 27672 22964 27678 22976
rect 27892 22973 27920 23072
rect 28092 23041 28120 23140
rect 28166 23128 28172 23180
rect 28224 23128 28230 23180
rect 28902 23128 28908 23180
rect 28960 23168 28966 23180
rect 29730 23168 29736 23180
rect 28960 23140 29736 23168
rect 28960 23128 28966 23140
rect 29730 23128 29736 23140
rect 29788 23128 29794 23180
rect 32858 23128 32864 23180
rect 32916 23128 32922 23180
rect 28350 23060 28356 23112
rect 28408 23060 28414 23112
rect 28442 23060 28448 23112
rect 28500 23060 28506 23112
rect 28721 23103 28779 23109
rect 28721 23069 28733 23103
rect 28767 23100 28779 23103
rect 28810 23100 28816 23112
rect 28767 23072 28816 23100
rect 28767 23069 28779 23072
rect 28721 23063 28779 23069
rect 28810 23060 28816 23072
rect 28868 23100 28874 23112
rect 28997 23103 29055 23109
rect 28997 23100 29009 23103
rect 28868 23072 29009 23100
rect 28868 23060 28874 23072
rect 28997 23069 29009 23072
rect 29043 23069 29055 23103
rect 28997 23063 29055 23069
rect 30650 23060 30656 23112
rect 30708 23060 30714 23112
rect 28077 23035 28135 23041
rect 28077 23001 28089 23035
rect 28123 23032 28135 23035
rect 28258 23032 28264 23044
rect 28123 23004 28264 23032
rect 28123 23001 28135 23004
rect 28077 22995 28135 23001
rect 28258 22992 28264 23004
rect 28316 22992 28322 23044
rect 28537 23035 28595 23041
rect 28537 23001 28549 23035
rect 28583 23032 28595 23035
rect 28626 23032 28632 23044
rect 28583 23004 28632 23032
rect 28583 23001 28595 23004
rect 28537 22995 28595 23001
rect 28626 22992 28632 23004
rect 28684 22992 28690 23044
rect 29018 23004 29408 23032
rect 27709 22967 27767 22973
rect 27709 22964 27721 22967
rect 27672 22936 27721 22964
rect 27672 22924 27678 22936
rect 27709 22933 27721 22936
rect 27755 22933 27767 22967
rect 27709 22927 27767 22933
rect 27877 22967 27935 22973
rect 27877 22933 27889 22967
rect 27923 22964 27935 22967
rect 29018 22964 29046 23004
rect 29380 22976 29408 23004
rect 27923 22936 29046 22964
rect 27923 22933 27935 22936
rect 27877 22927 27935 22933
rect 29086 22924 29092 22976
rect 29144 22924 29150 22976
rect 29362 22924 29368 22976
rect 29420 22924 29426 22976
rect 29546 22924 29552 22976
rect 29604 22964 29610 22976
rect 30742 22964 30748 22976
rect 29604 22936 30748 22964
rect 29604 22924 29610 22936
rect 30742 22924 30748 22936
rect 30800 22924 30806 22976
rect 1104 22874 38824 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 38824 22874
rect 1104 22800 38824 22822
rect 2777 22763 2835 22769
rect 2777 22729 2789 22763
rect 2823 22760 2835 22763
rect 2866 22760 2872 22772
rect 2823 22732 2872 22760
rect 2823 22729 2835 22732
rect 2777 22723 2835 22729
rect 2866 22720 2872 22732
rect 2924 22720 2930 22772
rect 3786 22720 3792 22772
rect 3844 22720 3850 22772
rect 4522 22720 4528 22772
rect 4580 22760 4586 22772
rect 4709 22763 4767 22769
rect 4709 22760 4721 22763
rect 4580 22732 4721 22760
rect 4580 22720 4586 22732
rect 4709 22729 4721 22732
rect 4755 22729 4767 22763
rect 4709 22723 4767 22729
rect 6362 22720 6368 22772
rect 6420 22720 6426 22772
rect 9125 22763 9183 22769
rect 9125 22729 9137 22763
rect 9171 22760 9183 22763
rect 9674 22760 9680 22772
rect 9171 22732 9680 22760
rect 9171 22729 9183 22732
rect 9125 22723 9183 22729
rect 9674 22720 9680 22732
rect 9732 22720 9738 22772
rect 9858 22720 9864 22772
rect 9916 22720 9922 22772
rect 13265 22763 13323 22769
rect 13265 22729 13277 22763
rect 13311 22760 13323 22763
rect 13630 22760 13636 22772
rect 13311 22732 13636 22760
rect 13311 22729 13323 22732
rect 13265 22723 13323 22729
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 13906 22760 13912 22772
rect 13740 22732 13912 22760
rect 3804 22692 3832 22720
rect 3344 22664 3832 22692
rect 3344 22633 3372 22664
rect 3602 22633 3608 22636
rect 3329 22627 3387 22633
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 3596 22624 3608 22633
rect 3563 22596 3608 22624
rect 3329 22587 3387 22593
rect 3596 22587 3608 22596
rect 3602 22584 3608 22587
rect 3660 22584 3666 22636
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22624 5043 22627
rect 5258 22624 5264 22636
rect 5031 22596 5264 22624
rect 5031 22593 5043 22596
rect 4985 22587 5043 22593
rect 5258 22584 5264 22596
rect 5316 22584 5322 22636
rect 5810 22584 5816 22636
rect 5868 22624 5874 22636
rect 6365 22627 6423 22633
rect 6365 22624 6377 22627
rect 5868 22596 6377 22624
rect 5868 22584 5874 22596
rect 6365 22593 6377 22596
rect 6411 22593 6423 22627
rect 6365 22587 6423 22593
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22624 7711 22627
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7699 22596 7757 22624
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 3237 22559 3295 22565
rect 3237 22525 3249 22559
rect 3283 22525 3295 22559
rect 3237 22519 3295 22525
rect 5077 22559 5135 22565
rect 5077 22525 5089 22559
rect 5123 22525 5135 22559
rect 5077 22519 5135 22525
rect 3252 22420 3280 22519
rect 5092 22488 5120 22519
rect 5442 22516 5448 22568
rect 5500 22516 5506 22568
rect 4264 22460 5120 22488
rect 5353 22491 5411 22497
rect 4062 22420 4068 22432
rect 3252 22392 4068 22420
rect 4062 22380 4068 22392
rect 4120 22420 4126 22432
rect 4264 22420 4292 22460
rect 5353 22457 5365 22491
rect 5399 22488 5411 22491
rect 5534 22488 5540 22500
rect 5399 22460 5540 22488
rect 5399 22457 5411 22460
rect 5353 22451 5411 22457
rect 5534 22448 5540 22460
rect 5592 22488 5598 22500
rect 6564 22488 6592 22587
rect 7282 22516 7288 22568
rect 7340 22516 7346 22568
rect 7484 22556 7512 22587
rect 8478 22584 8484 22636
rect 8536 22584 8542 22636
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22624 9551 22627
rect 9876 22624 9904 22720
rect 11882 22692 11888 22704
rect 11532 22664 11888 22692
rect 9539 22596 9904 22624
rect 9539 22593 9551 22596
rect 9493 22587 9551 22593
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 11532 22633 11560 22664
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 12434 22652 12440 22704
rect 12492 22652 12498 22704
rect 13740 22701 13768 22732
rect 13906 22720 13912 22732
rect 13964 22720 13970 22772
rect 15194 22720 15200 22772
rect 15252 22720 15258 22772
rect 17954 22760 17960 22772
rect 17880 22732 17960 22760
rect 13725 22695 13783 22701
rect 13725 22661 13737 22695
rect 13771 22661 13783 22695
rect 13725 22655 13783 22661
rect 14458 22652 14464 22704
rect 14516 22652 14522 22704
rect 17880 22701 17908 22732
rect 17954 22720 17960 22732
rect 18012 22720 18018 22772
rect 19429 22763 19487 22769
rect 19429 22729 19441 22763
rect 19475 22760 19487 22763
rect 19610 22760 19616 22772
rect 19475 22732 19616 22760
rect 19475 22729 19487 22732
rect 19429 22723 19487 22729
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 19797 22763 19855 22769
rect 19797 22729 19809 22763
rect 19843 22760 19855 22763
rect 20441 22763 20499 22769
rect 20441 22760 20453 22763
rect 19843 22732 20453 22760
rect 19843 22729 19855 22732
rect 19797 22723 19855 22729
rect 20441 22729 20453 22732
rect 20487 22760 20499 22763
rect 20530 22760 20536 22772
rect 20487 22732 20536 22760
rect 20487 22729 20499 22732
rect 20441 22723 20499 22729
rect 20530 22720 20536 22732
rect 20588 22760 20594 22772
rect 21174 22760 21180 22772
rect 20588 22732 21180 22760
rect 20588 22720 20594 22732
rect 21174 22720 21180 22732
rect 21232 22720 21238 22772
rect 21450 22720 21456 22772
rect 21508 22720 21514 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 22278 22760 22284 22772
rect 21591 22732 22284 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 22646 22720 22652 22772
rect 22704 22760 22710 22772
rect 22925 22763 22983 22769
rect 22925 22760 22937 22763
rect 22704 22732 22937 22760
rect 22704 22720 22710 22732
rect 22925 22729 22937 22732
rect 22971 22729 22983 22763
rect 22925 22723 22983 22729
rect 17865 22695 17923 22701
rect 17865 22661 17877 22695
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 18598 22652 18604 22704
rect 18656 22652 18662 22704
rect 20806 22692 20812 22704
rect 20548 22664 20812 22692
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 11112 22596 11529 22624
rect 11112 22584 11118 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 20346 22624 20352 22636
rect 11517 22587 11575 22593
rect 19352 22596 20352 22624
rect 8110 22556 8116 22568
rect 7484 22528 8116 22556
rect 8110 22516 8116 22528
rect 8168 22516 8174 22568
rect 8386 22516 8392 22568
rect 8444 22516 8450 22568
rect 8754 22516 8760 22568
rect 8812 22556 8818 22568
rect 8849 22559 8907 22565
rect 8849 22556 8861 22559
rect 8812 22528 8861 22556
rect 8812 22516 8818 22528
rect 8849 22525 8861 22528
rect 8895 22525 8907 22559
rect 8849 22519 8907 22525
rect 10134 22516 10140 22568
rect 10192 22516 10198 22568
rect 11790 22516 11796 22568
rect 11848 22516 11854 22568
rect 11882 22516 11888 22568
rect 11940 22556 11946 22568
rect 13449 22559 13507 22565
rect 13449 22556 13461 22559
rect 11940 22528 13461 22556
rect 11940 22516 11946 22528
rect 13449 22525 13461 22528
rect 13495 22556 13507 22559
rect 13495 22528 13584 22556
rect 13495 22525 13507 22528
rect 13449 22519 13507 22525
rect 5592 22460 6592 22488
rect 5592 22448 5598 22460
rect 13556 22432 13584 22528
rect 16850 22516 16856 22568
rect 16908 22556 16914 22568
rect 17310 22556 17316 22568
rect 16908 22528 17316 22556
rect 16908 22516 16914 22528
rect 17310 22516 17316 22528
rect 17368 22556 17374 22568
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 17368 22528 17601 22556
rect 17368 22516 17374 22528
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17589 22519 17647 22525
rect 19352 22432 19380 22596
rect 20346 22584 20352 22596
rect 20404 22584 20410 22636
rect 20548 22633 20576 22664
rect 20806 22652 20812 22664
rect 20864 22652 20870 22704
rect 21468 22633 21496 22720
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22593 20591 22627
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20533 22587 20591 22593
rect 20732 22596 21097 22624
rect 20732 22568 20760 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 19886 22516 19892 22568
rect 19944 22516 19950 22568
rect 20070 22516 20076 22568
rect 20128 22516 20134 22568
rect 20714 22516 20720 22568
rect 20772 22516 20778 22568
rect 20898 22516 20904 22568
rect 20956 22516 20962 22568
rect 21468 22556 21496 22587
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21784 22596 21833 22624
rect 21784 22584 21790 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 22830 22584 22836 22636
rect 22888 22584 22894 22636
rect 22940 22624 22968 22723
rect 24578 22720 24584 22772
rect 24636 22720 24642 22772
rect 25501 22763 25559 22769
rect 25501 22729 25513 22763
rect 25547 22760 25559 22763
rect 26418 22760 26424 22772
rect 25547 22732 26424 22760
rect 25547 22729 25559 22732
rect 25501 22723 25559 22729
rect 26418 22720 26424 22732
rect 26476 22720 26482 22772
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 27985 22763 28043 22769
rect 27488 22732 27844 22760
rect 27488 22720 27494 22732
rect 23382 22624 23388 22636
rect 22940 22596 23388 22624
rect 23382 22584 23388 22596
rect 23440 22624 23446 22636
rect 23477 22627 23535 22633
rect 23477 22624 23489 22627
rect 23440 22596 23489 22624
rect 23440 22584 23446 22596
rect 23477 22593 23489 22596
rect 23523 22593 23535 22627
rect 24121 22627 24179 22633
rect 24121 22624 24133 22627
rect 23477 22587 23535 22593
rect 23584 22596 24133 22624
rect 22097 22559 22155 22565
rect 22097 22556 22109 22559
rect 21468 22528 22109 22556
rect 22097 22525 22109 22528
rect 22143 22556 22155 22559
rect 22646 22556 22652 22568
rect 22143 22528 22652 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 22646 22516 22652 22528
rect 22704 22516 22710 22568
rect 23584 22565 23612 22596
rect 24121 22593 24133 22596
rect 24167 22624 24179 22627
rect 24596 22624 24624 22720
rect 25593 22695 25651 22701
rect 25593 22661 25605 22695
rect 25639 22661 25651 22695
rect 25593 22655 25651 22661
rect 25700 22664 26372 22692
rect 24167 22596 24624 22624
rect 24167 22593 24179 22596
rect 24121 22587 24179 22593
rect 25314 22584 25320 22636
rect 25372 22584 25378 22636
rect 25501 22627 25559 22633
rect 25501 22593 25513 22627
rect 25547 22624 25559 22627
rect 25608 22624 25636 22655
rect 25547 22596 25636 22624
rect 25547 22593 25559 22596
rect 25501 22587 25559 22593
rect 23017 22559 23075 22565
rect 23017 22525 23029 22559
rect 23063 22525 23075 22559
rect 23017 22519 23075 22525
rect 23569 22559 23627 22565
rect 23569 22525 23581 22559
rect 23615 22525 23627 22559
rect 25593 22559 25651 22565
rect 25593 22556 25605 22559
rect 23569 22519 23627 22525
rect 24412 22528 25605 22556
rect 22186 22448 22192 22500
rect 22244 22488 22250 22500
rect 23032 22488 23060 22519
rect 24412 22488 24440 22528
rect 25593 22525 25605 22528
rect 25639 22556 25651 22559
rect 25700 22556 25728 22664
rect 25869 22627 25927 22633
rect 25869 22624 25881 22627
rect 25792 22596 25881 22624
rect 25792 22568 25820 22596
rect 25869 22593 25881 22596
rect 25915 22624 25927 22627
rect 26237 22627 26295 22633
rect 26237 22624 26249 22627
rect 25915 22596 26249 22624
rect 25915 22593 25927 22596
rect 25869 22587 25927 22593
rect 26237 22593 26249 22596
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 25639 22528 25728 22556
rect 25639 22525 25651 22528
rect 25593 22519 25651 22525
rect 25774 22516 25780 22568
rect 25832 22516 25838 22568
rect 25958 22516 25964 22568
rect 26016 22516 26022 22568
rect 26344 22556 26372 22664
rect 26510 22584 26516 22636
rect 26568 22624 26574 22636
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 26568 22596 26985 22624
rect 26568 22584 26574 22596
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 27120 22596 27169 22624
rect 27120 22584 27126 22596
rect 27157 22593 27169 22596
rect 27203 22624 27215 22627
rect 27522 22624 27528 22636
rect 27203 22596 27528 22624
rect 27203 22593 27215 22596
rect 27157 22587 27215 22593
rect 27522 22584 27528 22596
rect 27580 22624 27586 22636
rect 27816 22633 27844 22732
rect 27985 22729 27997 22763
rect 28031 22760 28043 22763
rect 28166 22760 28172 22772
rect 28031 22732 28172 22760
rect 28031 22729 28043 22732
rect 27985 22723 28043 22729
rect 28166 22720 28172 22732
rect 28224 22720 28230 22772
rect 28261 22763 28319 22769
rect 28261 22729 28273 22763
rect 28307 22760 28319 22763
rect 28350 22760 28356 22772
rect 28307 22732 28356 22760
rect 28307 22729 28319 22732
rect 28261 22723 28319 22729
rect 28350 22720 28356 22732
rect 28408 22720 28414 22772
rect 28442 22720 28448 22772
rect 28500 22760 28506 22772
rect 29003 22763 29061 22769
rect 29003 22760 29015 22763
rect 28500 22732 29015 22760
rect 28500 22720 28506 22732
rect 29003 22729 29015 22732
rect 29049 22729 29061 22763
rect 29003 22723 29061 22729
rect 29089 22763 29147 22769
rect 29089 22729 29101 22763
rect 29135 22760 29147 22763
rect 29546 22760 29552 22772
rect 29135 22732 29552 22760
rect 29135 22729 29147 22732
rect 29089 22723 29147 22729
rect 28460 22664 29224 22692
rect 28460 22633 28488 22664
rect 29196 22636 29224 22664
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 27580 22596 27721 22624
rect 27580 22584 27586 22596
rect 27709 22593 27721 22596
rect 27755 22593 27767 22627
rect 27709 22587 27767 22593
rect 27801 22627 27859 22633
rect 27801 22593 27813 22627
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 28445 22627 28503 22633
rect 28445 22593 28457 22627
rect 28491 22593 28503 22627
rect 28445 22587 28503 22593
rect 28629 22627 28687 22633
rect 28629 22593 28641 22627
rect 28675 22624 28687 22627
rect 28902 22624 28908 22636
rect 28675 22596 28908 22624
rect 28675 22593 28687 22596
rect 28629 22587 28687 22593
rect 28902 22584 28908 22596
rect 28960 22584 28966 22636
rect 29178 22584 29184 22636
rect 29236 22584 29242 22636
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 26344 22528 27997 22556
rect 27985 22525 27997 22528
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 28537 22559 28595 22565
rect 28537 22525 28549 22559
rect 28583 22525 28595 22559
rect 28537 22519 28595 22525
rect 22244 22460 23060 22488
rect 23308 22460 24440 22488
rect 22244 22448 22250 22460
rect 23308 22432 23336 22460
rect 4120 22392 4292 22420
rect 4120 22380 4126 22392
rect 4522 22380 4528 22432
rect 4580 22420 4586 22432
rect 4985 22423 5043 22429
rect 4985 22420 4997 22423
rect 4580 22392 4997 22420
rect 4580 22380 4586 22392
rect 4985 22389 4997 22392
rect 5031 22389 5043 22423
rect 4985 22383 5043 22389
rect 6086 22380 6092 22432
rect 6144 22380 6150 22432
rect 6733 22423 6791 22429
rect 6733 22389 6745 22423
rect 6779 22420 6791 22423
rect 6914 22420 6920 22432
rect 6779 22392 6920 22420
rect 6779 22389 6791 22392
rect 6733 22383 6791 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 7558 22380 7564 22432
rect 7616 22380 7622 22432
rect 8662 22429 8668 22432
rect 8646 22423 8668 22429
rect 8646 22389 8658 22423
rect 8646 22383 8668 22389
rect 8662 22380 8668 22383
rect 8720 22380 8726 22432
rect 8757 22423 8815 22429
rect 8757 22389 8769 22423
rect 8803 22420 8815 22423
rect 9030 22420 9036 22432
rect 8803 22392 9036 22420
rect 8803 22389 8815 22392
rect 8757 22383 8815 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 10042 22380 10048 22432
rect 10100 22380 10106 22432
rect 10778 22380 10784 22432
rect 10836 22380 10842 22432
rect 13538 22380 13544 22432
rect 13596 22380 13602 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 19058 22420 19064 22432
rect 15620 22392 19064 22420
rect 15620 22380 15626 22392
rect 19058 22380 19064 22392
rect 19116 22380 19122 22432
rect 19334 22380 19340 22432
rect 19392 22380 19398 22432
rect 22462 22380 22468 22432
rect 22520 22380 22526 22432
rect 23290 22380 23296 22432
rect 23348 22380 23354 22432
rect 23750 22380 23756 22432
rect 23808 22380 23814 22432
rect 24026 22380 24032 22432
rect 24084 22380 24090 22432
rect 25777 22423 25835 22429
rect 25777 22389 25789 22423
rect 25823 22420 25835 22423
rect 27157 22423 27215 22429
rect 27157 22420 27169 22423
rect 25823 22392 27169 22420
rect 25823 22389 25835 22392
rect 25777 22383 25835 22389
rect 27157 22389 27169 22392
rect 27203 22389 27215 22423
rect 28000 22420 28028 22519
rect 28552 22488 28580 22519
rect 28718 22516 28724 22568
rect 28776 22516 28782 22568
rect 28902 22488 28908 22500
rect 28552 22460 28908 22488
rect 28902 22448 28908 22460
rect 28960 22488 28966 22500
rect 29288 22488 29316 22732
rect 29546 22720 29552 22732
rect 29604 22720 29610 22772
rect 29825 22763 29883 22769
rect 29825 22729 29837 22763
rect 29871 22729 29883 22763
rect 29825 22723 29883 22729
rect 29840 22692 29868 22723
rect 30558 22720 30564 22772
rect 30616 22720 30622 22772
rect 30834 22720 30840 22772
rect 30892 22720 30898 22772
rect 32861 22763 32919 22769
rect 32861 22729 32873 22763
rect 32907 22729 32919 22763
rect 32861 22723 32919 22729
rect 30055 22695 30113 22701
rect 30055 22692 30067 22695
rect 29840 22664 30067 22692
rect 30055 22661 30067 22664
rect 30101 22661 30113 22695
rect 30055 22655 30113 22661
rect 30742 22652 30748 22704
rect 30800 22652 30806 22704
rect 29454 22584 29460 22636
rect 29512 22584 29518 22636
rect 30190 22584 30196 22636
rect 30248 22584 30254 22636
rect 30282 22584 30288 22636
rect 30340 22584 30346 22636
rect 30374 22584 30380 22636
rect 30432 22584 30438 22636
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22624 30711 22627
rect 30760 22624 30788 22652
rect 30852 22633 30880 22720
rect 32876 22692 32904 22723
rect 32950 22720 32956 22772
rect 33008 22760 33014 22772
rect 33008 22732 33180 22760
rect 33008 22720 33014 22732
rect 32784 22664 32904 22692
rect 32784 22633 32812 22664
rect 32999 22661 33057 22667
rect 30699 22596 30788 22624
rect 30837 22627 30895 22633
rect 30699 22593 30711 22596
rect 30653 22587 30711 22593
rect 30837 22593 30849 22627
rect 30883 22593 30895 22627
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 30837 22587 30895 22593
rect 30944 22596 32781 22624
rect 29362 22516 29368 22568
rect 29420 22516 29426 22568
rect 29914 22516 29920 22568
rect 29972 22516 29978 22568
rect 28960 22460 29316 22488
rect 29380 22488 29408 22516
rect 30944 22488 30972 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32999 22627 33011 22661
rect 33045 22658 33057 22661
rect 33045 22627 33072 22658
rect 32999 22621 33072 22627
rect 32769 22587 32827 22593
rect 31294 22516 31300 22568
rect 31352 22556 31358 22568
rect 32493 22559 32551 22565
rect 32493 22556 32505 22559
rect 31352 22528 32505 22556
rect 31352 22516 31358 22528
rect 32493 22525 32505 22528
rect 32539 22525 32551 22559
rect 32493 22519 32551 22525
rect 32950 22516 32956 22568
rect 33008 22556 33014 22568
rect 33044 22556 33072 22621
rect 33152 22624 33180 22732
rect 33229 22695 33287 22701
rect 33229 22661 33241 22695
rect 33275 22692 33287 22695
rect 33505 22695 33563 22701
rect 33505 22692 33517 22695
rect 33275 22664 33517 22692
rect 33275 22661 33287 22664
rect 33229 22655 33287 22661
rect 33505 22661 33517 22664
rect 33551 22692 33563 22695
rect 33551 22664 33732 22692
rect 33551 22661 33563 22664
rect 33505 22655 33563 22661
rect 33704 22636 33732 22664
rect 33321 22627 33379 22633
rect 33321 22624 33333 22627
rect 33152 22596 33333 22624
rect 33321 22593 33333 22596
rect 33367 22593 33379 22627
rect 33321 22587 33379 22593
rect 33597 22627 33655 22633
rect 33597 22593 33609 22627
rect 33643 22593 33655 22627
rect 33597 22587 33655 22593
rect 33612 22556 33640 22587
rect 33686 22584 33692 22636
rect 33744 22584 33750 22636
rect 33008 22528 33640 22556
rect 33008 22516 33014 22528
rect 29380 22460 30972 22488
rect 32677 22491 32735 22497
rect 28960 22448 28966 22460
rect 32677 22457 32689 22491
rect 32723 22488 32735 22491
rect 33321 22491 33379 22497
rect 33321 22488 33333 22491
rect 32723 22460 33333 22488
rect 32723 22457 32735 22460
rect 32677 22451 32735 22457
rect 33321 22457 33333 22460
rect 33367 22457 33379 22491
rect 33321 22451 33379 22457
rect 29914 22420 29920 22432
rect 28000 22392 29920 22420
rect 27157 22383 27215 22389
rect 29914 22380 29920 22392
rect 29972 22380 29978 22432
rect 30742 22380 30748 22432
rect 30800 22380 30806 22432
rect 32582 22380 32588 22432
rect 32640 22380 32646 22432
rect 32858 22380 32864 22432
rect 32916 22420 32922 22432
rect 33045 22423 33103 22429
rect 33045 22420 33057 22423
rect 32916 22392 33057 22420
rect 32916 22380 32922 22392
rect 33045 22389 33057 22392
rect 33091 22389 33103 22423
rect 33045 22383 33103 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 3786 22176 3792 22228
rect 3844 22176 3850 22228
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 4028 22188 5304 22216
rect 4028 22176 4034 22188
rect 3804 22148 3832 22176
rect 3620 22120 3832 22148
rect 5276 22148 5304 22188
rect 5810 22176 5816 22228
rect 5868 22176 5874 22228
rect 5920 22188 12388 22216
rect 5920 22148 5948 22188
rect 5276 22120 5948 22148
rect 3620 22089 3648 22120
rect 8478 22108 8484 22160
rect 8536 22148 8542 22160
rect 8754 22148 8760 22160
rect 8536 22120 8760 22148
rect 8536 22108 8542 22120
rect 8754 22108 8760 22120
rect 8812 22108 8818 22160
rect 12360 22148 12388 22188
rect 12434 22176 12440 22228
rect 12492 22176 12498 22228
rect 13909 22219 13967 22225
rect 13909 22216 13921 22219
rect 12636 22188 13921 22216
rect 12636 22148 12664 22188
rect 13909 22185 13921 22188
rect 13955 22185 13967 22219
rect 17494 22216 17500 22228
rect 13909 22179 13967 22185
rect 16408 22188 17500 22216
rect 12360 22120 12664 22148
rect 3605 22083 3663 22089
rect 3605 22080 3617 22083
rect 3563 22052 3617 22080
rect 3605 22049 3617 22052
rect 3651 22080 3663 22083
rect 4341 22083 4399 22089
rect 4341 22080 4353 22083
rect 3651 22052 4353 22080
rect 3651 22049 3663 22052
rect 3605 22043 3663 22049
rect 4341 22049 4353 22052
rect 4387 22049 4399 22083
rect 12897 22083 12955 22089
rect 12897 22080 12909 22083
rect 4341 22043 4399 22049
rect 10980 22052 12909 22080
rect 10980 22024 11008 22052
rect 12897 22049 12909 22052
rect 12943 22049 12955 22083
rect 12897 22043 12955 22049
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 3360 21947 3418 21953
rect 3360 21913 3372 21947
rect 3406 21944 3418 21947
rect 3881 21947 3939 21953
rect 3881 21944 3893 21947
rect 3406 21916 3893 21944
rect 3406 21913 3418 21916
rect 3360 21907 3418 21913
rect 3881 21913 3893 21916
rect 3927 21913 3939 21947
rect 3881 21907 3939 21913
rect 3988 21888 4016 21975
rect 6914 21972 6920 22024
rect 6972 22021 6978 22024
rect 6972 21975 6984 22021
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 7285 22015 7343 22021
rect 7285 22012 7297 22015
rect 7239 21984 7297 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 7285 21981 7297 21984
rect 7331 22012 7343 22015
rect 8294 22012 8300 22024
rect 7331 21984 8300 22012
rect 7331 21981 7343 21984
rect 7285 21975 7343 21981
rect 6972 21972 6978 21975
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 4608 21947 4666 21953
rect 4608 21913 4620 21947
rect 4654 21944 4666 21947
rect 4798 21944 4804 21956
rect 4654 21916 4804 21944
rect 4654 21913 4666 21916
rect 4608 21907 4666 21913
rect 4798 21904 4804 21916
rect 4856 21904 4862 21956
rect 7558 21953 7564 21956
rect 7552 21907 7564 21953
rect 7558 21904 7564 21907
rect 7616 21904 7622 21956
rect 8478 21904 8484 21956
rect 8536 21944 8542 21956
rect 9508 21944 9536 21975
rect 10778 21972 10784 22024
rect 10836 22021 10842 22024
rect 10836 21975 10848 22021
rect 10836 21972 10842 21975
rect 10962 21972 10968 22024
rect 11020 21972 11026 22024
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 22012 11115 22015
rect 11514 22012 11520 22024
rect 11103 21984 11520 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 11514 21972 11520 21984
rect 11572 21972 11578 22024
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 8536 21916 9536 21944
rect 8536 21904 8542 21916
rect 2225 21879 2283 21885
rect 2225 21845 2237 21879
rect 2271 21876 2283 21879
rect 3234 21876 3240 21888
rect 2271 21848 3240 21876
rect 2271 21845 2283 21848
rect 2225 21839 2283 21845
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 3970 21836 3976 21888
rect 4028 21836 4034 21888
rect 5718 21836 5724 21888
rect 5776 21836 5782 21888
rect 8680 21885 8708 21916
rect 8665 21879 8723 21885
rect 8665 21845 8677 21879
rect 8711 21845 8723 21879
rect 8665 21839 8723 21845
rect 8938 21836 8944 21888
rect 8996 21836 9002 21888
rect 9030 21836 9036 21888
rect 9088 21876 9094 21888
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9088 21848 9689 21876
rect 9088 21836 9094 21848
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 12912 21876 12940 22043
rect 13173 22015 13231 22021
rect 13173 21981 13185 22015
rect 13219 22012 13231 22015
rect 13219 21984 13308 22012
rect 13219 21981 13231 21984
rect 13173 21975 13231 21981
rect 13280 21956 13308 21984
rect 13262 21904 13268 21956
rect 13320 21904 13326 21956
rect 13924 21944 13952 22179
rect 13998 22040 14004 22092
rect 14056 22080 14062 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 14056 22052 14105 22080
rect 14056 22040 14062 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 16408 22021 16436 22188
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 18049 22219 18107 22225
rect 18049 22185 18061 22219
rect 18095 22216 18107 22219
rect 18138 22216 18144 22228
rect 18095 22188 18144 22216
rect 18095 22185 18107 22188
rect 18049 22179 18107 22185
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 20901 22219 20959 22225
rect 20901 22216 20913 22219
rect 20864 22188 20913 22216
rect 20864 22176 20870 22188
rect 20901 22185 20913 22188
rect 20947 22185 20959 22219
rect 20901 22179 20959 22185
rect 22094 22176 22100 22228
rect 22152 22176 22158 22228
rect 25958 22176 25964 22228
rect 26016 22216 26022 22228
rect 26053 22219 26111 22225
rect 26053 22216 26065 22219
rect 26016 22188 26065 22216
rect 26016 22176 26022 22188
rect 26053 22185 26065 22188
rect 26099 22185 26111 22219
rect 26053 22179 26111 22185
rect 29178 22176 29184 22228
rect 29236 22216 29242 22228
rect 30009 22219 30067 22225
rect 30009 22216 30021 22219
rect 29236 22188 30021 22216
rect 29236 22176 29242 22188
rect 30009 22185 30021 22188
rect 30055 22216 30067 22219
rect 30282 22216 30288 22228
rect 30055 22188 30288 22216
rect 30055 22185 30067 22188
rect 30009 22179 30067 22185
rect 30282 22176 30288 22188
rect 30340 22176 30346 22228
rect 30374 22176 30380 22228
rect 30432 22216 30438 22228
rect 30561 22219 30619 22225
rect 30561 22216 30573 22219
rect 30432 22188 30573 22216
rect 30432 22176 30438 22188
rect 30561 22185 30573 22188
rect 30607 22185 30619 22219
rect 30561 22179 30619 22185
rect 32582 22176 32588 22228
rect 32640 22176 32646 22228
rect 33594 22216 33600 22228
rect 33152 22188 33600 22216
rect 17126 22108 17132 22160
rect 17184 22148 17190 22160
rect 17681 22151 17739 22157
rect 17681 22148 17693 22151
rect 17184 22120 17693 22148
rect 17184 22108 17190 22120
rect 17681 22117 17693 22120
rect 17727 22117 17739 22151
rect 17681 22111 17739 22117
rect 18708 22120 20116 22148
rect 18708 22089 18736 22120
rect 20088 22092 20116 22120
rect 20530 22108 20536 22160
rect 20588 22108 20594 22160
rect 20622 22108 20628 22160
rect 20680 22148 20686 22160
rect 24394 22148 24400 22160
rect 20680 22120 24400 22148
rect 20680 22108 20686 22120
rect 24394 22108 24400 22120
rect 24452 22108 24458 22160
rect 29914 22108 29920 22160
rect 29972 22148 29978 22160
rect 31294 22148 31300 22160
rect 29972 22120 31300 22148
rect 29972 22108 29978 22120
rect 31294 22108 31300 22120
rect 31352 22108 31358 22160
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 18739 22052 18773 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 20070 22040 20076 22092
rect 20128 22040 20134 22092
rect 23014 22080 23020 22092
rect 20180 22052 23020 22080
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 16393 22015 16451 22021
rect 16393 22012 16405 22015
rect 14369 21975 14427 21981
rect 14568 21984 16405 22012
rect 14384 21944 14412 21975
rect 13924 21916 14412 21944
rect 13998 21876 14004 21888
rect 12912 21848 14004 21876
rect 9677 21839 9735 21845
rect 13998 21836 14004 21848
rect 14056 21876 14062 21888
rect 14568 21876 14596 21984
rect 16393 21981 16405 21984
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 16574 21972 16580 22024
rect 16632 22012 16638 22024
rect 16669 22015 16727 22021
rect 16669 22012 16681 22015
rect 16632 21984 16681 22012
rect 16632 21972 16638 21984
rect 16669 21981 16681 21984
rect 16715 21981 16727 22015
rect 17497 22015 17555 22021
rect 17497 22012 17509 22015
rect 16669 21975 16727 21981
rect 17420 21984 17509 22012
rect 14642 21904 14648 21956
rect 14700 21944 14706 21956
rect 15197 21947 15255 21953
rect 15197 21944 15209 21947
rect 14700 21916 15209 21944
rect 14700 21904 14706 21916
rect 15197 21913 15209 21916
rect 15243 21913 15255 21947
rect 15197 21907 15255 21913
rect 15473 21947 15531 21953
rect 15473 21913 15485 21947
rect 15519 21944 15531 21947
rect 17420 21944 17448 21984
rect 17497 21981 17509 21984
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 19334 22012 19340 22024
rect 18463 21984 19340 22012
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 15519 21916 17448 21944
rect 15519 21913 15531 21916
rect 15473 21907 15531 21913
rect 14056 21848 14596 21876
rect 14056 21836 14062 21848
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15381 21879 15439 21885
rect 15381 21876 15393 21879
rect 15160 21848 15393 21876
rect 15160 21836 15166 21848
rect 15381 21845 15393 21848
rect 15427 21845 15439 21879
rect 15381 21839 15439 21845
rect 15562 21836 15568 21888
rect 15620 21836 15626 21888
rect 15746 21836 15752 21888
rect 15804 21836 15810 21888
rect 17420 21885 17448 21916
rect 18690 21904 18696 21956
rect 18748 21944 18754 21956
rect 20180 21944 20208 22052
rect 23014 22040 23020 22052
rect 23072 22040 23078 22092
rect 23661 22083 23719 22089
rect 23661 22049 23673 22083
rect 23707 22080 23719 22083
rect 23750 22080 23756 22092
rect 23707 22052 23756 22080
rect 23707 22049 23719 22052
rect 23661 22043 23719 22049
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 27062 22080 27068 22092
rect 26252 22052 27068 22080
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 22012 22339 22015
rect 22462 22012 22468 22024
rect 22327 21984 22468 22012
rect 22327 21981 22339 21984
rect 22281 21975 22339 21981
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 23566 21972 23572 22024
rect 23624 21972 23630 22024
rect 26252 22021 26280 22052
rect 27062 22040 27068 22052
rect 27120 22040 27126 22092
rect 28902 22040 28908 22092
rect 28960 22040 28966 22092
rect 28997 22083 29055 22089
rect 28997 22049 29009 22083
rect 29043 22080 29055 22083
rect 30742 22080 30748 22092
rect 29043 22052 29868 22080
rect 29043 22049 29055 22052
rect 28997 22043 29055 22049
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 22012 26479 22015
rect 26510 22012 26516 22024
rect 26467 21984 26516 22012
rect 26467 21981 26479 21984
rect 26421 21975 26479 21981
rect 26510 21972 26516 21984
rect 26568 21972 26574 22024
rect 28718 21972 28724 22024
rect 28776 21972 28782 22024
rect 29089 22015 29147 22021
rect 29089 21981 29101 22015
rect 29135 21981 29147 22015
rect 29089 21975 29147 21981
rect 18748 21916 20208 21944
rect 29104 21944 29132 21975
rect 29270 21972 29276 22024
rect 29328 21972 29334 22024
rect 29730 21972 29736 22024
rect 29788 21972 29794 22024
rect 29840 21944 29868 22052
rect 30208 22052 30748 22080
rect 30208 22021 30236 22052
rect 30742 22040 30748 22052
rect 30800 22040 30806 22092
rect 32033 22083 32091 22089
rect 32033 22049 32045 22083
rect 32079 22080 32091 22083
rect 32600 22080 32628 22176
rect 32079 22052 32628 22080
rect 32079 22049 32091 22052
rect 32033 22043 32091 22049
rect 29917 22015 29975 22021
rect 29917 21981 29929 22015
rect 29963 22012 29975 22015
rect 30193 22015 30251 22021
rect 30193 22012 30205 22015
rect 29963 21984 30205 22012
rect 29963 21981 29975 21984
rect 29917 21975 29975 21981
rect 30193 21981 30205 21984
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 30469 22015 30527 22021
rect 30469 21981 30481 22015
rect 30515 21981 30527 22015
rect 30469 21975 30527 21981
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30760 22012 30788 22040
rect 30607 21984 30788 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 30484 21944 30512 21975
rect 31754 21972 31760 22024
rect 31812 21972 31818 22024
rect 31849 22015 31907 22021
rect 31849 21981 31861 22015
rect 31895 22012 31907 22015
rect 32122 22012 32128 22024
rect 31895 21984 32128 22012
rect 31895 21981 31907 21984
rect 31849 21975 31907 21981
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 32493 22015 32551 22021
rect 32493 21981 32505 22015
rect 32539 21981 32551 22015
rect 32493 21975 32551 21981
rect 29104 21916 29316 21944
rect 29840 21916 30512 21944
rect 18748 21904 18754 21916
rect 29288 21888 29316 21916
rect 17405 21879 17463 21885
rect 17405 21845 17417 21879
rect 17451 21845 17463 21879
rect 17405 21839 17463 21845
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 18874 21876 18880 21888
rect 18555 21848 18880 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 18874 21836 18880 21848
rect 18932 21836 18938 21888
rect 20714 21836 20720 21888
rect 20772 21876 20778 21888
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20772 21848 20913 21876
rect 20772 21836 20778 21848
rect 20901 21845 20913 21848
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21876 21143 21879
rect 21910 21876 21916 21888
rect 21131 21848 21916 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 23934 21836 23940 21888
rect 23992 21876 23998 21888
rect 24486 21876 24492 21888
rect 23992 21848 24492 21876
rect 23992 21836 23998 21848
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 28534 21836 28540 21888
rect 28592 21836 28598 21888
rect 29270 21836 29276 21888
rect 29328 21876 29334 21888
rect 29549 21879 29607 21885
rect 29549 21876 29561 21879
rect 29328 21848 29561 21876
rect 29328 21836 29334 21848
rect 29549 21845 29561 21848
rect 29595 21845 29607 21879
rect 29549 21839 29607 21845
rect 30374 21836 30380 21888
rect 30432 21836 30438 21888
rect 30484 21876 30512 21916
rect 30650 21904 30656 21956
rect 30708 21953 30714 21956
rect 30708 21947 30730 21953
rect 30718 21913 30730 21947
rect 30708 21907 30730 21913
rect 30837 21947 30895 21953
rect 30837 21913 30849 21947
rect 30883 21944 30895 21947
rect 32309 21947 32367 21953
rect 32309 21944 32321 21947
rect 30883 21916 32321 21944
rect 30883 21913 30895 21916
rect 30837 21907 30895 21913
rect 32309 21913 32321 21916
rect 32355 21913 32367 21947
rect 32508 21944 32536 21975
rect 32582 21972 32588 22024
rect 32640 22012 32646 22024
rect 32769 22015 32827 22021
rect 32769 22012 32781 22015
rect 32640 21984 32781 22012
rect 32640 21972 32646 21984
rect 32769 21981 32781 21984
rect 32815 21981 32827 22015
rect 32769 21975 32827 21981
rect 32858 21972 32864 22024
rect 32916 21972 32922 22024
rect 33152 22021 33180 22188
rect 33594 22176 33600 22188
rect 33652 22176 33658 22228
rect 33689 22219 33747 22225
rect 33689 22185 33701 22219
rect 33735 22185 33747 22219
rect 33689 22179 33747 22185
rect 33704 22148 33732 22179
rect 33688 22120 33732 22148
rect 33688 22080 33716 22120
rect 33688 22052 33732 22080
rect 33704 22024 33732 22052
rect 33137 22015 33195 22021
rect 33137 21981 33149 22015
rect 33183 21981 33195 22015
rect 33137 21975 33195 21981
rect 33413 22015 33471 22021
rect 33413 21981 33425 22015
rect 33459 22006 33471 22015
rect 33686 22012 33692 22024
rect 33612 22006 33692 22012
rect 33459 21984 33692 22006
rect 33459 21981 33640 21984
rect 33413 21978 33640 21981
rect 33413 21975 33471 21978
rect 33686 21972 33692 21984
rect 33744 21972 33750 22024
rect 32876 21944 32904 21972
rect 33873 21947 33931 21953
rect 33873 21944 33885 21947
rect 32508 21916 32904 21944
rect 33336 21916 33885 21944
rect 32309 21907 32367 21913
rect 30708 21904 30714 21907
rect 30852 21876 30880 21907
rect 30484 21848 30880 21876
rect 32033 21879 32091 21885
rect 32033 21845 32045 21879
rect 32079 21876 32091 21879
rect 32214 21876 32220 21888
rect 32079 21848 32220 21876
rect 32079 21845 32091 21848
rect 32033 21839 32091 21845
rect 32214 21836 32220 21848
rect 32272 21836 32278 21888
rect 32677 21879 32735 21885
rect 32677 21845 32689 21879
rect 32723 21876 32735 21879
rect 32953 21879 33011 21885
rect 32953 21876 32965 21879
rect 32723 21848 32965 21876
rect 32723 21845 32735 21848
rect 32677 21839 32735 21845
rect 32953 21845 32965 21848
rect 32999 21876 33011 21879
rect 33042 21876 33048 21888
rect 32999 21848 33048 21876
rect 32999 21845 33011 21848
rect 32953 21839 33011 21845
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 33134 21836 33140 21888
rect 33192 21876 33198 21888
rect 33336 21885 33364 21916
rect 33873 21913 33885 21916
rect 33919 21913 33931 21947
rect 33873 21907 33931 21913
rect 33321 21879 33379 21885
rect 33321 21876 33333 21879
rect 33192 21848 33333 21876
rect 33192 21836 33198 21848
rect 33321 21845 33333 21848
rect 33367 21845 33379 21879
rect 33321 21839 33379 21845
rect 33502 21836 33508 21888
rect 33560 21836 33566 21888
rect 33668 21879 33726 21885
rect 33668 21845 33680 21879
rect 33714 21876 33726 21879
rect 33778 21876 33784 21888
rect 33714 21848 33784 21876
rect 33714 21845 33726 21848
rect 33668 21839 33726 21845
rect 33778 21836 33784 21848
rect 33836 21836 33842 21888
rect 1104 21786 38824 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 38824 21786
rect 1104 21712 38824 21734
rect 4798 21632 4804 21684
rect 4856 21632 4862 21684
rect 5258 21632 5264 21684
rect 5316 21672 5322 21684
rect 5537 21675 5595 21681
rect 5537 21672 5549 21675
rect 5316 21644 5549 21672
rect 5316 21632 5322 21644
rect 5537 21641 5549 21644
rect 5583 21641 5595 21675
rect 5537 21635 5595 21641
rect 5718 21632 5724 21684
rect 5776 21632 5782 21684
rect 7282 21632 7288 21684
rect 7340 21632 7346 21684
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 8386 21672 8392 21684
rect 8067 21644 8392 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8386 21632 8392 21644
rect 8444 21632 8450 21684
rect 8846 21632 8852 21684
rect 8904 21632 8910 21684
rect 8938 21632 8944 21684
rect 8996 21632 9002 21684
rect 11514 21632 11520 21684
rect 11572 21672 11578 21684
rect 13630 21672 13636 21684
rect 11572 21644 13636 21672
rect 11572 21632 11578 21644
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14553 21675 14611 21681
rect 14553 21641 14565 21675
rect 14599 21672 14611 21675
rect 15286 21672 15292 21684
rect 14599 21644 15292 21672
rect 14599 21641 14611 21644
rect 14553 21635 14611 21641
rect 15286 21632 15292 21644
rect 15344 21632 15350 21684
rect 15457 21675 15515 21681
rect 15457 21641 15469 21675
rect 15503 21672 15515 21675
rect 15562 21672 15568 21684
rect 15503 21644 15568 21672
rect 15503 21641 15515 21644
rect 15457 21635 15515 21641
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 15746 21632 15752 21684
rect 15804 21632 15810 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 16669 21675 16727 21681
rect 16669 21672 16681 21675
rect 16632 21644 16681 21672
rect 16632 21632 16638 21644
rect 16669 21641 16681 21644
rect 16715 21641 16727 21675
rect 22002 21672 22008 21684
rect 16669 21635 16727 21641
rect 20824 21644 22008 21672
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 4062 21536 4068 21548
rect 3292 21508 4068 21536
rect 3292 21496 3298 21508
rect 4062 21496 4068 21508
rect 4120 21536 4126 21548
rect 5736 21536 5764 21632
rect 5810 21564 5816 21616
rect 5868 21604 5874 21616
rect 6365 21607 6423 21613
rect 6365 21604 6377 21607
rect 5868 21576 6377 21604
rect 5868 21564 5874 21576
rect 6365 21573 6377 21576
rect 6411 21573 6423 21607
rect 6365 21567 6423 21573
rect 7101 21607 7159 21613
rect 7101 21573 7113 21607
rect 7147 21604 7159 21607
rect 8956 21604 8984 21632
rect 7147 21576 7420 21604
rect 7147 21573 7159 21576
rect 7101 21567 7159 21573
rect 6089 21539 6147 21545
rect 6089 21536 6101 21539
rect 4120 21508 5672 21536
rect 5736 21508 6101 21536
rect 4120 21496 4126 21508
rect 4706 21428 4712 21480
rect 4764 21428 4770 21480
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 5534 21468 5540 21480
rect 5491 21440 5540 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 5534 21428 5540 21440
rect 5592 21428 5598 21480
rect 5644 21468 5672 21508
rect 6089 21505 6101 21508
rect 6135 21536 6147 21539
rect 6512 21539 6570 21545
rect 6512 21536 6524 21539
rect 6135 21508 6524 21536
rect 6135 21505 6147 21508
rect 6089 21499 6147 21505
rect 6512 21505 6524 21508
rect 6558 21505 6570 21539
rect 6512 21499 6570 21505
rect 7190 21496 7196 21548
rect 7248 21496 7254 21548
rect 7392 21545 7420 21576
rect 8036 21576 8984 21604
rect 8036 21545 8064 21576
rect 9030 21564 9036 21616
rect 9088 21564 9094 21616
rect 10042 21564 10048 21616
rect 10100 21613 10106 21616
rect 10100 21604 10112 21613
rect 10100 21576 10145 21604
rect 10100 21567 10112 21576
rect 10100 21564 10106 21567
rect 7377 21539 7435 21545
rect 7377 21505 7389 21539
rect 7423 21536 7435 21539
rect 7837 21539 7895 21545
rect 7837 21536 7849 21539
rect 7423 21508 7849 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7837 21505 7849 21508
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 8021 21539 8079 21545
rect 8021 21505 8033 21539
rect 8067 21505 8079 21539
rect 8021 21499 8079 21505
rect 6733 21471 6791 21477
rect 6733 21468 6745 21471
rect 5644 21440 6745 21468
rect 6733 21437 6745 21440
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 4724 21400 4752 21428
rect 6641 21403 6699 21409
rect 6641 21400 6653 21403
rect 4724 21372 6653 21400
rect 6641 21369 6653 21372
rect 6687 21369 6699 21403
rect 7852 21400 7880 21499
rect 8110 21496 8116 21548
rect 8168 21496 8174 21548
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21536 8355 21539
rect 8386 21536 8392 21548
rect 8343 21508 8392 21536
rect 8343 21505 8355 21508
rect 8297 21499 8355 21505
rect 8386 21496 8392 21508
rect 8444 21496 8450 21548
rect 8481 21539 8539 21545
rect 8481 21505 8493 21539
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 8573 21539 8631 21545
rect 8573 21505 8585 21539
rect 8619 21536 8631 21539
rect 9048 21536 9076 21564
rect 11532 21545 11560 21632
rect 12066 21564 12072 21616
rect 12124 21604 12130 21616
rect 14737 21607 14795 21613
rect 14737 21604 14749 21607
rect 12124 21576 12282 21604
rect 14384 21576 14749 21604
rect 12124 21564 12130 21576
rect 8619 21508 9076 21536
rect 10321 21539 10379 21545
rect 8619 21505 8631 21508
rect 8573 21499 8631 21505
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 10367 21508 11529 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 8496 21468 8524 21499
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14384 21545 14412 21576
rect 14737 21573 14749 21576
rect 14783 21604 14795 21607
rect 15010 21604 15016 21616
rect 14783 21576 15016 21604
rect 14783 21573 14795 21576
rect 14737 21567 14795 21573
rect 15010 21564 15016 21576
rect 15068 21604 15074 21616
rect 15657 21607 15715 21613
rect 15657 21604 15669 21607
rect 15068 21576 15669 21604
rect 15068 21564 15074 21576
rect 15657 21573 15669 21576
rect 15703 21573 15715 21607
rect 15764 21604 15792 21632
rect 15933 21607 15991 21613
rect 15933 21604 15945 21607
rect 15764 21576 15945 21604
rect 15657 21567 15715 21573
rect 15933 21573 15945 21576
rect 15979 21573 15991 21607
rect 15933 21567 15991 21573
rect 17052 21576 18000 21604
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 14240 21508 14381 21536
rect 14240 21496 14246 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21505 14703 21539
rect 14645 21499 14703 21505
rect 8404 21440 8524 21468
rect 8404 21400 8432 21440
rect 8662 21428 8668 21480
rect 8720 21468 8726 21480
rect 8849 21471 8907 21477
rect 8849 21468 8861 21471
rect 8720 21440 8861 21468
rect 8720 21428 8726 21440
rect 8849 21437 8861 21440
rect 8895 21437 8907 21471
rect 8849 21431 8907 21437
rect 8570 21400 8576 21412
rect 7852 21372 8576 21400
rect 6641 21363 6699 21369
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 8864 21400 8892 21431
rect 11790 21428 11796 21480
rect 11848 21428 11854 21480
rect 14660 21468 14688 21499
rect 15102 21496 15108 21548
rect 15160 21496 15166 21548
rect 15562 21496 15568 21548
rect 15620 21496 15626 21548
rect 15580 21468 15608 21496
rect 14660 21440 15608 21468
rect 15654 21428 15660 21480
rect 15712 21468 15718 21480
rect 17052 21468 17080 21576
rect 17402 21496 17408 21548
rect 17460 21496 17466 21548
rect 17494 21496 17500 21548
rect 17552 21536 17558 21548
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17552 21508 17693 21536
rect 17552 21496 17558 21508
rect 17681 21505 17693 21508
rect 17727 21536 17739 21539
rect 17770 21536 17776 21548
rect 17727 21508 17776 21536
rect 17727 21505 17739 21508
rect 17681 21499 17739 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 17972 21545 18000 21576
rect 17957 21539 18015 21545
rect 17957 21505 17969 21539
rect 18003 21536 18015 21539
rect 18782 21536 18788 21548
rect 18003 21508 18788 21536
rect 18003 21505 18015 21508
rect 17957 21499 18015 21505
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20714 21536 20720 21548
rect 20119 21508 20720 21536
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 20824 21545 20852 21644
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23293 21675 23351 21681
rect 23293 21672 23305 21675
rect 22888 21644 23305 21672
rect 22888 21632 22894 21644
rect 23293 21641 23305 21644
rect 23339 21641 23351 21675
rect 24679 21675 24737 21681
rect 24679 21672 24691 21675
rect 23293 21635 23351 21641
rect 23777 21644 24691 21672
rect 21910 21564 21916 21616
rect 21968 21564 21974 21616
rect 23658 21604 23664 21616
rect 23308 21576 23664 21604
rect 20809 21539 20867 21545
rect 20809 21505 20821 21539
rect 20855 21505 20867 21539
rect 20809 21499 20867 21505
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 20956 21508 21097 21536
rect 20956 21496 20962 21508
rect 21085 21505 21097 21508
rect 21131 21505 21143 21539
rect 21085 21499 21143 21505
rect 15712 21440 17080 21468
rect 15712 21428 15718 21440
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 8941 21403 8999 21409
rect 8941 21400 8953 21403
rect 8864 21372 8953 21400
rect 8941 21369 8953 21372
rect 8987 21369 8999 21403
rect 8941 21363 8999 21369
rect 14369 21403 14427 21409
rect 14369 21369 14381 21403
rect 14415 21400 14427 21403
rect 15194 21400 15200 21412
rect 14415 21372 15200 21400
rect 14415 21369 14427 21372
rect 14369 21363 14427 21369
rect 15194 21360 15200 21372
rect 15252 21360 15258 21412
rect 15286 21360 15292 21412
rect 15344 21360 15350 21412
rect 15749 21403 15807 21409
rect 15749 21400 15761 21403
rect 15396 21372 15761 21400
rect 3789 21335 3847 21341
rect 3789 21301 3801 21335
rect 3835 21332 3847 21335
rect 3970 21332 3976 21344
rect 3835 21304 3976 21332
rect 3835 21301 3847 21304
rect 3789 21295 3847 21301
rect 3970 21292 3976 21304
rect 4028 21332 4034 21344
rect 5074 21332 5080 21344
rect 4028 21304 5080 21332
rect 4028 21292 4034 21304
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 8110 21292 8116 21344
rect 8168 21332 8174 21344
rect 8665 21335 8723 21341
rect 8665 21332 8677 21335
rect 8168 21304 8677 21332
rect 8168 21292 8174 21304
rect 8665 21301 8677 21304
rect 8711 21301 8723 21335
rect 8665 21295 8723 21301
rect 12802 21292 12808 21344
rect 12860 21332 12866 21344
rect 13262 21332 13268 21344
rect 12860 21304 13268 21332
rect 12860 21292 12866 21304
rect 13262 21292 13268 21304
rect 13320 21292 13326 21344
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14918 21332 14924 21344
rect 14516 21304 14924 21332
rect 14516 21292 14522 21304
rect 14918 21292 14924 21304
rect 14976 21332 14982 21344
rect 15396 21332 15424 21372
rect 15749 21369 15761 21372
rect 15795 21369 15807 21403
rect 15749 21363 15807 21369
rect 20070 21360 20076 21412
rect 20128 21400 20134 21412
rect 20272 21400 20300 21431
rect 20990 21428 20996 21480
rect 21048 21468 21054 21480
rect 23308 21477 23336 21576
rect 23658 21564 23664 21576
rect 23716 21564 23722 21616
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21536 23627 21539
rect 23777 21536 23805 21644
rect 24679 21641 24691 21644
rect 24725 21641 24737 21675
rect 24679 21635 24737 21641
rect 30374 21632 30380 21684
rect 30432 21672 30438 21684
rect 30650 21672 30656 21684
rect 30432 21644 30656 21672
rect 30432 21632 30438 21644
rect 30650 21632 30656 21644
rect 30708 21632 30714 21684
rect 31754 21632 31760 21684
rect 31812 21681 31818 21684
rect 31812 21672 31821 21681
rect 31812 21644 31857 21672
rect 31812 21635 31821 21644
rect 31812 21632 31818 21635
rect 32122 21632 32128 21684
rect 32180 21632 32186 21684
rect 32858 21632 32864 21684
rect 32916 21672 32922 21684
rect 33502 21672 33508 21684
rect 32916 21644 33508 21672
rect 32916 21632 32922 21644
rect 33502 21632 33508 21644
rect 33560 21632 33566 21684
rect 28626 21604 28632 21616
rect 24688 21576 28632 21604
rect 23615 21508 23805 21536
rect 23615 21505 23627 21508
rect 23569 21499 23627 21505
rect 23934 21496 23940 21548
rect 23992 21536 23998 21548
rect 24121 21539 24179 21545
rect 24121 21536 24133 21539
rect 23992 21508 24133 21536
rect 23992 21496 23998 21508
rect 24121 21505 24133 21508
rect 24167 21505 24179 21539
rect 24121 21499 24179 21505
rect 24213 21539 24271 21545
rect 24213 21505 24225 21539
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21048 21440 21557 21468
rect 21048 21428 21054 21440
rect 21545 21437 21557 21440
rect 21591 21468 21603 21471
rect 23293 21471 23351 21477
rect 21591 21440 22094 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 20128 21372 20300 21400
rect 20809 21403 20867 21409
rect 20128 21360 20134 21372
rect 20809 21369 20821 21403
rect 20855 21400 20867 21403
rect 21174 21400 21180 21412
rect 20855 21372 21180 21400
rect 20855 21369 20867 21372
rect 20809 21363 20867 21369
rect 21174 21360 21180 21372
rect 21232 21360 21238 21412
rect 14976 21304 15424 21332
rect 14976 21292 14982 21304
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 16758 21332 16764 21344
rect 15528 21304 16764 21332
rect 15528 21292 15534 21304
rect 16758 21292 16764 21304
rect 16816 21332 16822 21344
rect 17034 21332 17040 21344
rect 16816 21304 17040 21332
rect 16816 21292 16822 21304
rect 17034 21292 17040 21304
rect 17092 21292 17098 21344
rect 17865 21335 17923 21341
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 17954 21332 17960 21344
rect 17911 21304 17960 21332
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 19702 21292 19708 21344
rect 19760 21292 19766 21344
rect 22066 21332 22094 21440
rect 23293 21437 23305 21471
rect 23339 21437 23351 21471
rect 24228 21468 24256 21499
rect 24486 21496 24492 21548
rect 24544 21536 24550 21548
rect 24581 21539 24639 21545
rect 24581 21536 24593 21539
rect 24544 21508 24593 21536
rect 24544 21496 24550 21508
rect 24581 21505 24593 21508
rect 24627 21505 24639 21539
rect 24581 21499 24639 21505
rect 23293 21431 23351 21437
rect 24136 21440 24256 21468
rect 24305 21471 24363 21477
rect 24136 21344 24164 21440
rect 24305 21437 24317 21471
rect 24351 21437 24363 21471
rect 24305 21431 24363 21437
rect 24320 21400 24348 21431
rect 24394 21428 24400 21480
rect 24452 21468 24458 21480
rect 24688 21468 24716 21576
rect 28626 21564 28632 21576
rect 28684 21564 28690 21616
rect 24762 21496 24768 21548
rect 24820 21496 24826 21548
rect 24857 21539 24915 21545
rect 24857 21505 24869 21539
rect 24903 21505 24915 21539
rect 24857 21499 24915 21505
rect 25961 21539 26019 21545
rect 25961 21505 25973 21539
rect 26007 21505 26019 21539
rect 25961 21499 26019 21505
rect 24452 21440 24716 21468
rect 24452 21428 24458 21440
rect 24780 21400 24808 21496
rect 24320 21372 24808 21400
rect 22189 21335 22247 21341
rect 22189 21332 22201 21335
rect 22066 21304 22201 21332
rect 22189 21301 22201 21304
rect 22235 21332 22247 21335
rect 23382 21332 23388 21344
rect 22235 21304 23388 21332
rect 22235 21301 22247 21304
rect 22189 21295 22247 21301
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23937 21335 23995 21341
rect 23937 21332 23949 21335
rect 23523 21304 23949 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23937 21301 23949 21304
rect 23983 21301 23995 21335
rect 23937 21295 23995 21301
rect 24118 21292 24124 21344
rect 24176 21332 24182 21344
rect 24872 21332 24900 21499
rect 25976 21468 26004 21499
rect 26050 21496 26056 21548
rect 26108 21536 26114 21548
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 26108 21508 26249 21536
rect 26108 21496 26114 21508
rect 26237 21505 26249 21508
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 31849 21539 31907 21545
rect 31849 21505 31861 21539
rect 31895 21505 31907 21539
rect 31849 21499 31907 21505
rect 26329 21471 26387 21477
rect 26329 21468 26341 21471
rect 25976 21440 26341 21468
rect 26329 21437 26341 21440
rect 26375 21468 26387 21471
rect 26510 21468 26516 21480
rect 26375 21440 26516 21468
rect 26375 21437 26387 21440
rect 26329 21431 26387 21437
rect 26510 21428 26516 21440
rect 26568 21428 26574 21480
rect 31680 21400 31708 21499
rect 31864 21468 31892 21499
rect 31938 21496 31944 21548
rect 31996 21536 32002 21548
rect 32876 21545 32904 21632
rect 32953 21607 33011 21613
rect 32953 21573 32965 21607
rect 32999 21604 33011 21607
rect 32999 21576 33364 21604
rect 32999 21573 33011 21576
rect 32953 21567 33011 21573
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 31996 21508 32321 21536
rect 31996 21496 32002 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 32493 21539 32551 21545
rect 32493 21505 32505 21539
rect 32539 21536 32551 21539
rect 32861 21539 32919 21545
rect 32539 21508 32720 21536
rect 32539 21505 32551 21508
rect 32493 21499 32551 21505
rect 32398 21468 32404 21480
rect 31864 21440 32404 21468
rect 32398 21428 32404 21440
rect 32456 21428 32462 21480
rect 32508 21400 32536 21499
rect 32585 21471 32643 21477
rect 32585 21437 32597 21471
rect 32631 21437 32643 21471
rect 32692 21468 32720 21508
rect 32861 21505 32873 21539
rect 32907 21505 32919 21539
rect 32861 21499 32919 21505
rect 33042 21496 33048 21548
rect 33100 21536 33106 21548
rect 33336 21545 33364 21576
rect 33137 21539 33195 21545
rect 33137 21536 33149 21539
rect 33100 21508 33149 21536
rect 33100 21496 33106 21508
rect 33137 21505 33149 21508
rect 33183 21505 33195 21539
rect 33137 21499 33195 21505
rect 33321 21539 33379 21545
rect 33321 21505 33333 21539
rect 33367 21505 33379 21539
rect 33321 21499 33379 21505
rect 33229 21471 33287 21477
rect 33229 21468 33241 21471
rect 32692 21440 33241 21468
rect 32585 21431 32643 21437
rect 33229 21437 33241 21440
rect 33275 21437 33287 21471
rect 33229 21431 33287 21437
rect 31496 21372 32536 21400
rect 31496 21344 31524 21372
rect 24176 21304 24900 21332
rect 24176 21292 24182 21304
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 26605 21335 26663 21341
rect 26605 21301 26617 21335
rect 26651 21332 26663 21335
rect 27614 21332 27620 21344
rect 26651 21304 27620 21332
rect 26651 21301 26663 21304
rect 26605 21295 26663 21301
rect 27614 21292 27620 21304
rect 27672 21292 27678 21344
rect 31478 21292 31484 21344
rect 31536 21292 31542 21344
rect 31570 21292 31576 21344
rect 31628 21332 31634 21344
rect 32600 21332 32628 21431
rect 31628 21304 32628 21332
rect 31628 21292 31634 21304
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 4706 21088 4712 21140
rect 4764 21128 4770 21140
rect 5169 21131 5227 21137
rect 5169 21128 5181 21131
rect 4764 21100 5181 21128
rect 4764 21088 4770 21100
rect 5169 21097 5181 21100
rect 5215 21097 5227 21131
rect 5169 21091 5227 21097
rect 5261 21131 5319 21137
rect 5261 21097 5273 21131
rect 5307 21128 5319 21131
rect 5350 21128 5356 21140
rect 5307 21100 5356 21128
rect 5307 21097 5319 21100
rect 5261 21091 5319 21097
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 5534 21088 5540 21140
rect 5592 21088 5598 21140
rect 9030 21088 9036 21140
rect 9088 21088 9094 21140
rect 9401 21131 9459 21137
rect 9401 21097 9413 21131
rect 9447 21128 9459 21131
rect 10134 21128 10140 21140
rect 9447 21100 10140 21128
rect 9447 21097 9459 21100
rect 9401 21091 9459 21097
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 11790 21088 11796 21140
rect 11848 21088 11854 21140
rect 12066 21088 12072 21140
rect 12124 21088 12130 21140
rect 17678 21088 17684 21140
rect 17736 21128 17742 21140
rect 18601 21131 18659 21137
rect 18601 21128 18613 21131
rect 17736 21100 18613 21128
rect 17736 21088 17742 21100
rect 18601 21097 18613 21100
rect 18647 21097 18659 21131
rect 18601 21091 18659 21097
rect 19702 21088 19708 21140
rect 19760 21088 19766 21140
rect 19996 21100 22692 21128
rect 9048 21060 9076 21088
rect 14829 21063 14887 21069
rect 9048 21032 9168 21060
rect 5258 20952 5264 21004
rect 5316 20992 5322 21004
rect 5353 20995 5411 21001
rect 5353 20992 5365 20995
rect 5316 20964 5365 20992
rect 5316 20952 5322 20964
rect 5353 20961 5365 20964
rect 5399 20961 5411 20995
rect 5353 20955 5411 20961
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 9033 20995 9091 21001
rect 9033 20992 9045 20995
rect 8168 20964 9045 20992
rect 8168 20952 8174 20964
rect 9033 20961 9045 20964
rect 9079 20961 9091 20995
rect 9033 20955 9091 20961
rect 5074 20884 5080 20936
rect 5132 20884 5138 20936
rect 5442 20884 5448 20936
rect 5500 20884 5506 20936
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20924 5687 20927
rect 6086 20924 6092 20936
rect 5675 20896 6092 20924
rect 5675 20893 5687 20896
rect 5629 20887 5687 20893
rect 6086 20884 6092 20896
rect 6144 20884 6150 20936
rect 9140 20933 9168 21032
rect 14829 21029 14841 21063
rect 14875 21060 14887 21063
rect 15013 21063 15071 21069
rect 15013 21060 15025 21063
rect 14875 21032 15025 21060
rect 14875 21029 14887 21032
rect 14829 21023 14887 21029
rect 15013 21029 15025 21032
rect 15059 21029 15071 21063
rect 15013 21023 15071 21029
rect 15102 21020 15108 21072
rect 15160 21020 15166 21072
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 15243 20964 19334 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 11977 20927 12035 20933
rect 11977 20893 11989 20927
rect 12023 20893 12035 20927
rect 11977 20887 12035 20893
rect 11992 20856 12020 20887
rect 14090 20884 14096 20936
rect 14148 20924 14154 20936
rect 14642 20924 14648 20936
rect 14148 20896 14648 20924
rect 14148 20884 14154 20896
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 11072 20828 12020 20856
rect 14844 20856 14872 20887
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 14976 20896 15021 20924
rect 15286 20900 15292 20936
rect 14976 20884 14982 20896
rect 15120 20884 15292 20900
rect 15344 20924 15350 20936
rect 15565 20927 15623 20933
rect 15565 20924 15577 20927
rect 15344 20896 15577 20924
rect 15344 20884 15350 20896
rect 15565 20893 15577 20896
rect 15611 20893 15623 20927
rect 15565 20887 15623 20893
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20924 16451 20927
rect 16574 20924 16580 20936
rect 16439 20896 16580 20924
rect 16439 20893 16451 20896
rect 16393 20887 16451 20893
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20893 16727 20927
rect 16669 20887 16727 20893
rect 15120 20872 15332 20884
rect 15120 20856 15148 20872
rect 14844 20828 15148 20856
rect 11072 20800 11100 20828
rect 11054 20748 11060 20800
rect 11112 20748 11118 20800
rect 11992 20788 12020 20828
rect 15378 20816 15384 20868
rect 15436 20816 15442 20868
rect 16684 20856 16712 20887
rect 17954 20884 17960 20936
rect 18012 20924 18018 20936
rect 18012 20896 18078 20924
rect 18012 20884 18018 20896
rect 16850 20856 16856 20868
rect 16684 20828 16856 20856
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 16945 20859 17003 20865
rect 16945 20825 16957 20859
rect 16991 20825 17003 20859
rect 16945 20819 17003 20825
rect 15654 20788 15660 20800
rect 11992 20760 15660 20788
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 15749 20791 15807 20797
rect 15749 20757 15761 20791
rect 15795 20788 15807 20791
rect 15838 20788 15844 20800
rect 15795 20760 15844 20788
rect 15795 20757 15807 20760
rect 15749 20751 15807 20757
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 16577 20791 16635 20797
rect 16577 20757 16589 20791
rect 16623 20788 16635 20791
rect 16960 20788 16988 20819
rect 18690 20816 18696 20868
rect 18748 20816 18754 20868
rect 19306 20856 19334 20964
rect 19720 20933 19748 21088
rect 19996 20933 20024 21100
rect 22557 21063 22615 21069
rect 22557 21029 22569 21063
rect 22603 21029 22615 21063
rect 22557 21023 22615 21029
rect 20809 20995 20867 21001
rect 20809 20961 20821 20995
rect 20855 20992 20867 20995
rect 21542 20992 21548 21004
rect 20855 20964 21548 20992
rect 20855 20961 20867 20964
rect 20809 20955 20867 20961
rect 21542 20952 21548 20964
rect 21600 20952 21606 21004
rect 22572 20936 22600 21023
rect 22664 20936 22692 21100
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 25866 21128 25872 21140
rect 25556 21100 25872 21128
rect 25556 21088 25562 21100
rect 25866 21088 25872 21100
rect 25924 21128 25930 21140
rect 25961 21131 26019 21137
rect 25961 21128 25973 21131
rect 25924 21100 25973 21128
rect 25924 21088 25930 21100
rect 25961 21097 25973 21100
rect 26007 21097 26019 21131
rect 27893 21131 27951 21137
rect 27893 21128 27905 21131
rect 25961 21091 26019 21097
rect 26620 21100 27905 21128
rect 25332 21060 25360 21088
rect 26620 21060 26648 21100
rect 27893 21097 27905 21100
rect 27939 21097 27951 21131
rect 27893 21091 27951 21097
rect 28442 21088 28448 21140
rect 28500 21128 28506 21140
rect 28500 21100 28764 21128
rect 28500 21088 28506 21100
rect 25332 21032 26648 21060
rect 27614 21020 27620 21072
rect 27672 21020 27678 21072
rect 28534 21020 28540 21072
rect 28592 21020 28598 21072
rect 28736 21069 28764 21100
rect 30374 21088 30380 21140
rect 30432 21128 30438 21140
rect 30469 21131 30527 21137
rect 30469 21128 30481 21131
rect 30432 21100 30481 21128
rect 30432 21088 30438 21100
rect 30469 21097 30481 21100
rect 30515 21097 30527 21131
rect 30469 21091 30527 21097
rect 33134 21088 33140 21140
rect 33192 21088 33198 21140
rect 28721 21063 28779 21069
rect 28721 21029 28733 21063
rect 28767 21029 28779 21063
rect 28721 21023 28779 21029
rect 28810 21020 28816 21072
rect 28868 21060 28874 21072
rect 31570 21060 31576 21072
rect 28868 21032 31576 21060
rect 28868 21020 28874 21032
rect 31570 21020 31576 21032
rect 31628 21020 31634 21072
rect 26050 20992 26056 21004
rect 25332 20964 26056 20992
rect 25332 20936 25360 20964
rect 26050 20952 26056 20964
rect 26108 20952 26114 21004
rect 27433 20995 27491 21001
rect 27433 20961 27445 20995
rect 27479 20992 27491 20995
rect 27632 20992 27660 21020
rect 28552 20992 28580 21020
rect 29181 20995 29239 21001
rect 29181 20992 29193 20995
rect 27479 20964 27660 20992
rect 28092 20964 29193 20992
rect 27479 20961 27491 20964
rect 27433 20955 27491 20961
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19981 20927 20039 20933
rect 19981 20893 19993 20927
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 22554 20884 22560 20936
rect 22612 20884 22618 20936
rect 22646 20884 22652 20936
rect 22704 20884 22710 20936
rect 25314 20884 25320 20936
rect 25372 20884 25378 20936
rect 25682 20884 25688 20936
rect 25740 20924 25746 20936
rect 25961 20927 26019 20933
rect 25961 20924 25973 20927
rect 25740 20896 25973 20924
rect 25740 20884 25746 20896
rect 25961 20893 25973 20896
rect 26007 20893 26019 20927
rect 25961 20887 26019 20893
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20924 27675 20927
rect 27982 20924 27988 20936
rect 27663 20896 27988 20924
rect 27663 20893 27675 20896
rect 27617 20887 27675 20893
rect 27982 20884 27988 20896
rect 28040 20884 28046 20936
rect 28092 20933 28120 20964
rect 29181 20961 29193 20964
rect 29227 20961 29239 20995
rect 29181 20955 29239 20961
rect 28077 20927 28135 20933
rect 28077 20893 28089 20927
rect 28123 20893 28135 20927
rect 28077 20887 28135 20893
rect 28442 20884 28448 20936
rect 28500 20884 28506 20936
rect 28534 20884 28540 20936
rect 28592 20884 28598 20936
rect 28629 20927 28687 20933
rect 28629 20893 28641 20927
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 20806 20856 20812 20868
rect 19306 20828 20812 20856
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 21082 20816 21088 20868
rect 21140 20816 21146 20868
rect 22741 20859 22799 20865
rect 22741 20856 22753 20859
rect 22310 20828 22753 20856
rect 22741 20825 22753 20828
rect 22787 20825 22799 20859
rect 22741 20819 22799 20825
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 23440 20828 25544 20856
rect 23440 20816 23446 20828
rect 16623 20760 16988 20788
rect 16623 20757 16635 20760
rect 16577 20751 16635 20757
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 18417 20791 18475 20797
rect 18417 20788 18429 20791
rect 17368 20760 18429 20788
rect 17368 20748 17374 20760
rect 18417 20757 18429 20760
rect 18463 20757 18475 20791
rect 18417 20751 18475 20757
rect 19518 20748 19524 20800
rect 19576 20748 19582 20800
rect 19978 20748 19984 20800
rect 20036 20788 20042 20800
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 20036 20760 20085 20788
rect 20036 20748 20042 20760
rect 20073 20757 20085 20760
rect 20119 20757 20131 20791
rect 20073 20751 20131 20757
rect 20162 20748 20168 20800
rect 20220 20788 20226 20800
rect 23750 20788 23756 20800
rect 20220 20760 23756 20788
rect 20220 20748 20226 20760
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 25406 20748 25412 20800
rect 25464 20748 25470 20800
rect 25516 20788 25544 20828
rect 25590 20816 25596 20868
rect 25648 20816 25654 20868
rect 25774 20816 25780 20868
rect 25832 20816 25838 20868
rect 28169 20859 28227 20865
rect 28169 20825 28181 20859
rect 28215 20825 28227 20859
rect 28169 20819 28227 20825
rect 28261 20859 28319 20865
rect 28261 20825 28273 20859
rect 28307 20856 28319 20859
rect 28350 20856 28356 20868
rect 28307 20828 28356 20856
rect 28307 20825 28319 20828
rect 28261 20819 28319 20825
rect 26050 20788 26056 20800
rect 25516 20760 26056 20788
rect 26050 20748 26056 20760
rect 26108 20748 26114 20800
rect 26326 20748 26332 20800
rect 26384 20748 26390 20800
rect 27706 20748 27712 20800
rect 27764 20788 27770 20800
rect 27801 20791 27859 20797
rect 27801 20788 27813 20791
rect 27764 20760 27813 20788
rect 27764 20748 27770 20760
rect 27801 20757 27813 20760
rect 27847 20757 27859 20791
rect 28184 20788 28212 20819
rect 28350 20816 28356 20828
rect 28408 20856 28414 20868
rect 28644 20856 28672 20887
rect 28718 20884 28724 20936
rect 28776 20924 28782 20936
rect 28997 20927 29055 20933
rect 28997 20924 29009 20927
rect 28776 20896 29009 20924
rect 28776 20884 28782 20896
rect 28997 20893 29009 20896
rect 29043 20893 29055 20927
rect 28997 20887 29055 20893
rect 30098 20884 30104 20936
rect 30156 20924 30162 20936
rect 31297 20927 31355 20933
rect 31297 20924 31309 20927
rect 30156 20896 31309 20924
rect 30156 20884 30162 20896
rect 31297 20893 31309 20896
rect 31343 20893 31355 20927
rect 31297 20887 31355 20893
rect 31478 20884 31484 20936
rect 31536 20884 31542 20936
rect 33045 20927 33103 20933
rect 33045 20893 33057 20927
rect 33091 20893 33103 20927
rect 33045 20887 33103 20893
rect 28408 20828 28672 20856
rect 28408 20816 28414 20828
rect 30282 20816 30288 20868
rect 30340 20816 30346 20868
rect 31386 20816 31392 20868
rect 31444 20856 31450 20868
rect 31665 20859 31723 20865
rect 31665 20856 31677 20859
rect 31444 20828 31677 20856
rect 31444 20816 31450 20828
rect 31665 20825 31677 20828
rect 31711 20825 31723 20859
rect 31665 20819 31723 20825
rect 33060 20800 33088 20887
rect 28626 20788 28632 20800
rect 28184 20760 28632 20788
rect 27801 20751 27859 20757
rect 28626 20748 28632 20760
rect 28684 20748 28690 20800
rect 33042 20748 33048 20800
rect 33100 20748 33106 20800
rect 1104 20698 38824 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 38824 20698
rect 1104 20624 38824 20646
rect 4062 20544 4068 20596
rect 4120 20584 4126 20596
rect 15194 20584 15200 20596
rect 4120 20556 15200 20584
rect 4120 20544 4126 20556
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 16574 20544 16580 20596
rect 16632 20584 16638 20596
rect 16945 20587 17003 20593
rect 16945 20584 16957 20587
rect 16632 20556 16957 20584
rect 16632 20544 16638 20556
rect 16945 20553 16957 20556
rect 16991 20553 17003 20587
rect 20622 20584 20628 20596
rect 16945 20547 17003 20553
rect 17052 20556 20628 20584
rect 13078 20516 13084 20528
rect 12406 20488 13084 20516
rect 9677 20451 9735 20457
rect 9677 20417 9689 20451
rect 9723 20417 9735 20451
rect 9677 20411 9735 20417
rect 9692 20380 9720 20411
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 11054 20448 11060 20460
rect 9824 20420 11060 20448
rect 9824 20408 9830 20420
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 11609 20451 11667 20457
rect 11609 20417 11621 20451
rect 11655 20448 11667 20451
rect 11698 20448 11704 20460
rect 11655 20420 11704 20448
rect 11655 20417 11667 20420
rect 11609 20411 11667 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 11974 20380 11980 20392
rect 9692 20352 11980 20380
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 12069 20383 12127 20389
rect 12069 20349 12081 20383
rect 12115 20380 12127 20383
rect 12406 20380 12434 20488
rect 13078 20476 13084 20488
rect 13136 20516 13142 20528
rect 13383 20519 13441 20525
rect 13383 20516 13395 20519
rect 13136 20488 13395 20516
rect 13136 20476 13142 20488
rect 13383 20485 13395 20488
rect 13429 20485 13441 20519
rect 13383 20479 13441 20485
rect 13538 20457 13544 20460
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 13508 20451 13544 20457
rect 12575 20420 13400 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 12115 20352 12434 20380
rect 12621 20383 12679 20389
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12621 20349 12633 20383
rect 12667 20380 12679 20383
rect 12710 20380 12716 20392
rect 12667 20352 12716 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 12805 20383 12863 20389
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13262 20380 13268 20392
rect 13035 20352 13268 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 11606 20272 11612 20324
rect 11664 20312 11670 20324
rect 12161 20315 12219 20321
rect 12161 20312 12173 20315
rect 11664 20284 12173 20312
rect 11664 20272 11670 20284
rect 12161 20281 12173 20284
rect 12207 20281 12219 20315
rect 12161 20275 12219 20281
rect 12526 20272 12532 20324
rect 12584 20312 12590 20324
rect 12820 20312 12848 20343
rect 13262 20340 13268 20352
rect 13320 20340 13326 20392
rect 13372 20380 13400 20420
rect 13508 20417 13520 20451
rect 13508 20411 13544 20417
rect 13538 20408 13544 20411
rect 13596 20408 13602 20460
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20448 14795 20451
rect 15010 20448 15016 20460
rect 14783 20420 15016 20448
rect 14783 20417 14795 20420
rect 14737 20411 14795 20417
rect 15010 20408 15016 20420
rect 15068 20448 15074 20460
rect 17052 20448 17080 20556
rect 20622 20544 20628 20556
rect 20680 20544 20686 20596
rect 20714 20544 20720 20596
rect 20772 20544 20778 20596
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 21140 20556 21373 20584
rect 21140 20544 21146 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 21821 20587 21879 20593
rect 21821 20553 21833 20587
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 22189 20587 22247 20593
rect 22189 20553 22201 20587
rect 22235 20584 22247 20587
rect 24397 20587 24455 20593
rect 24397 20584 24409 20587
rect 22235 20556 24409 20584
rect 22235 20553 22247 20556
rect 22189 20547 22247 20553
rect 24397 20553 24409 20556
rect 24443 20553 24455 20587
rect 25406 20584 25412 20596
rect 24397 20547 24455 20553
rect 24596 20556 25412 20584
rect 19245 20519 19303 20525
rect 15068 20420 17080 20448
rect 17236 20488 19012 20516
rect 15068 20408 15074 20420
rect 13998 20380 14004 20392
rect 13372 20352 14004 20380
rect 13998 20340 14004 20352
rect 14056 20340 14062 20392
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 15102 20380 15108 20392
rect 14507 20352 15108 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 16850 20340 16856 20392
rect 16908 20380 16914 20392
rect 17236 20380 17264 20488
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20448 17371 20451
rect 17954 20448 17960 20460
rect 17359 20420 17960 20448
rect 17359 20417 17371 20420
rect 17313 20411 17371 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 18046 20408 18052 20460
rect 18104 20408 18110 20460
rect 18984 20457 19012 20488
rect 19245 20485 19257 20519
rect 19291 20516 19303 20519
rect 19518 20516 19524 20528
rect 19291 20488 19524 20516
rect 19291 20485 19303 20488
rect 19245 20479 19303 20485
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 19978 20476 19984 20528
rect 20036 20476 20042 20528
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 16908 20352 17264 20380
rect 16908 20340 16914 20352
rect 17402 20340 17408 20392
rect 17460 20340 17466 20392
rect 17494 20340 17500 20392
rect 17552 20340 17558 20392
rect 17770 20340 17776 20392
rect 17828 20340 17834 20392
rect 18892 20380 18920 20411
rect 20806 20408 20812 20460
rect 20864 20408 20870 20460
rect 21545 20451 21603 20457
rect 21545 20417 21557 20451
rect 21591 20448 21603 20451
rect 21836 20448 21864 20547
rect 23290 20516 23296 20528
rect 21591 20420 21864 20448
rect 22020 20488 23296 20516
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 20824 20380 20852 20408
rect 22020 20380 22048 20488
rect 23290 20476 23296 20488
rect 23348 20516 23354 20528
rect 23348 20488 23796 20516
rect 23348 20476 23354 20488
rect 22554 20448 22560 20460
rect 22296 20420 22560 20448
rect 18892 20352 19104 20380
rect 20824 20352 22048 20380
rect 12584 20284 12848 20312
rect 13633 20315 13691 20321
rect 12584 20272 12590 20284
rect 13633 20281 13645 20315
rect 13679 20312 13691 20315
rect 14734 20312 14740 20324
rect 13679 20284 14740 20312
rect 13679 20281 13691 20284
rect 13633 20275 13691 20281
rect 14734 20272 14740 20284
rect 14792 20272 14798 20324
rect 19076 20256 19104 20352
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 22296 20389 22324 20420
rect 22554 20408 22560 20420
rect 22612 20448 22618 20460
rect 22833 20451 22891 20457
rect 22833 20448 22845 20451
rect 22612 20420 22845 20448
rect 22612 20408 22618 20420
rect 22833 20417 22845 20420
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 23474 20408 23480 20460
rect 23532 20408 23538 20460
rect 23566 20408 23572 20460
rect 23624 20448 23630 20460
rect 23768 20457 23796 20488
rect 24118 20476 24124 20528
rect 24176 20476 24182 20528
rect 24596 20516 24624 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 25869 20587 25927 20593
rect 25869 20584 25881 20587
rect 25832 20556 25881 20584
rect 25832 20544 25838 20556
rect 25869 20553 25881 20556
rect 25915 20553 25927 20587
rect 25869 20547 25927 20553
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 27764 20556 28212 20584
rect 27764 20544 27770 20556
rect 28184 20525 28212 20556
rect 28350 20544 28356 20596
rect 28408 20544 28414 20596
rect 28629 20587 28687 20593
rect 28629 20553 28641 20587
rect 28675 20584 28687 20587
rect 28718 20584 28724 20596
rect 28675 20556 28724 20584
rect 28675 20553 28687 20556
rect 28629 20547 28687 20553
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 31757 20587 31815 20593
rect 31757 20584 31769 20587
rect 30944 20556 31769 20584
rect 30944 20525 30972 20556
rect 31757 20553 31769 20556
rect 31803 20584 31815 20587
rect 31938 20584 31944 20596
rect 31803 20556 31944 20584
rect 31803 20553 31815 20556
rect 31757 20547 31815 20553
rect 31938 20544 31944 20556
rect 31996 20544 32002 20596
rect 32585 20587 32643 20593
rect 32585 20553 32597 20587
rect 32631 20553 32643 20587
rect 32585 20547 32643 20553
rect 27801 20519 27859 20525
rect 24320 20488 24624 20516
rect 26068 20488 27476 20516
rect 24212 20473 24270 20479
rect 23661 20451 23719 20457
rect 23661 20448 23673 20451
rect 23624 20420 23673 20448
rect 23624 20408 23630 20420
rect 23661 20417 23673 20420
rect 23707 20417 23719 20451
rect 23661 20411 23719 20417
rect 23753 20451 23811 20457
rect 23753 20417 23765 20451
rect 23799 20417 23811 20451
rect 23753 20411 23811 20417
rect 23842 20408 23848 20460
rect 23900 20457 23906 20460
rect 23900 20451 23949 20457
rect 23900 20417 23903 20451
rect 23937 20417 23949 20451
rect 23900 20411 23949 20417
rect 24029 20451 24087 20457
rect 24029 20417 24041 20451
rect 24075 20417 24087 20451
rect 24212 20439 24224 20473
rect 24258 20472 24270 20473
rect 24320 20472 24348 20488
rect 24258 20444 24348 20472
rect 24673 20451 24731 20457
rect 24258 20439 24270 20444
rect 24212 20433 24270 20439
rect 24029 20411 24087 20417
rect 24673 20417 24685 20451
rect 24719 20417 24731 20451
rect 24673 20411 24731 20417
rect 23900 20408 23906 20411
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 22152 20352 22293 20380
rect 22152 20340 22158 20352
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 22281 20343 22339 20349
rect 22462 20340 22468 20392
rect 22520 20340 22526 20392
rect 23293 20383 23351 20389
rect 23293 20349 23305 20383
rect 23339 20380 23351 20383
rect 23584 20380 23612 20408
rect 24044 20380 24072 20411
rect 23339 20352 23612 20380
rect 23952 20352 24072 20380
rect 24688 20380 24716 20411
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 24949 20451 25007 20457
rect 24949 20448 24961 20451
rect 24912 20420 24961 20448
rect 24912 20408 24918 20420
rect 24949 20417 24961 20420
rect 24995 20417 25007 20451
rect 24949 20411 25007 20417
rect 25133 20451 25191 20457
rect 25133 20417 25145 20451
rect 25179 20417 25191 20451
rect 25133 20411 25191 20417
rect 25148 20380 25176 20411
rect 25314 20408 25320 20460
rect 25372 20408 25378 20460
rect 25409 20451 25467 20457
rect 25409 20417 25421 20451
rect 25455 20448 25467 20451
rect 25498 20448 25504 20460
rect 25455 20420 25504 20448
rect 25455 20417 25467 20420
rect 25409 20411 25467 20417
rect 25498 20408 25504 20420
rect 25556 20408 25562 20460
rect 25593 20451 25651 20457
rect 25593 20417 25605 20451
rect 25639 20448 25651 20451
rect 25682 20448 25688 20460
rect 25639 20420 25688 20448
rect 25639 20417 25651 20420
rect 25593 20411 25651 20417
rect 25682 20408 25688 20420
rect 25740 20408 25746 20460
rect 26068 20457 26096 20488
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20448 25835 20451
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 25823 20420 26065 20448
rect 25823 20417 25835 20420
rect 25777 20411 25835 20417
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 26326 20408 26332 20460
rect 26384 20408 26390 20460
rect 24688 20352 25176 20380
rect 23339 20349 23351 20352
rect 23293 20343 23351 20349
rect 22186 20272 22192 20324
rect 22244 20312 22250 20324
rect 22480 20312 22508 20340
rect 22244 20284 22508 20312
rect 22244 20272 22250 20284
rect 22830 20272 22836 20324
rect 22888 20312 22894 20324
rect 23109 20315 23167 20321
rect 23109 20312 23121 20315
rect 22888 20284 23121 20312
rect 22888 20272 22894 20284
rect 23109 20281 23121 20284
rect 23155 20281 23167 20315
rect 23109 20275 23167 20281
rect 23382 20272 23388 20324
rect 23440 20312 23446 20324
rect 23477 20315 23535 20321
rect 23477 20312 23489 20315
rect 23440 20284 23489 20312
rect 23440 20272 23446 20284
rect 23477 20281 23489 20284
rect 23523 20281 23535 20315
rect 23477 20275 23535 20281
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 9493 20247 9551 20253
rect 9493 20244 9505 20247
rect 9364 20216 9505 20244
rect 9364 20204 9370 20216
rect 9493 20213 9505 20216
rect 9539 20213 9551 20247
rect 9493 20207 9551 20213
rect 9858 20204 9864 20256
rect 9916 20204 9922 20256
rect 11882 20204 11888 20256
rect 11940 20204 11946 20256
rect 12710 20204 12716 20256
rect 12768 20244 12774 20256
rect 13081 20247 13139 20253
rect 13081 20244 13093 20247
rect 12768 20216 13093 20244
rect 12768 20204 12774 20216
rect 13081 20213 13093 20216
rect 13127 20213 13139 20247
rect 13081 20207 13139 20213
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 13780 20216 14565 20244
rect 13780 20204 13786 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 18046 20244 18052 20256
rect 17920 20216 18052 20244
rect 17920 20204 17926 20216
rect 18046 20204 18052 20216
rect 18104 20204 18110 20256
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 23566 20204 23572 20256
rect 23624 20244 23630 20256
rect 23952 20244 23980 20352
rect 25148 20312 25176 20352
rect 25406 20312 25412 20324
rect 25148 20284 25412 20312
rect 25406 20272 25412 20284
rect 25464 20272 25470 20324
rect 26142 20272 26148 20324
rect 26200 20272 26206 20324
rect 26237 20315 26295 20321
rect 26237 20281 26249 20315
rect 26283 20281 26295 20315
rect 26344 20312 26372 20408
rect 27448 20389 27476 20488
rect 27801 20485 27813 20519
rect 27847 20516 27859 20519
rect 27985 20519 28043 20525
rect 27985 20516 27997 20519
rect 27847 20488 27997 20516
rect 27847 20485 27859 20488
rect 27801 20479 27859 20485
rect 27985 20485 27997 20488
rect 28031 20485 28043 20519
rect 27985 20479 28043 20485
rect 28169 20519 28227 20525
rect 28169 20485 28181 20519
rect 28215 20485 28227 20519
rect 30929 20519 30987 20525
rect 28169 20479 28227 20485
rect 28828 20488 29132 20516
rect 27614 20408 27620 20460
rect 27672 20448 27678 20460
rect 28828 20457 28856 20488
rect 29104 20460 29132 20488
rect 29196 20488 30144 20516
rect 27709 20451 27767 20457
rect 27709 20448 27721 20451
rect 27672 20420 27721 20448
rect 27672 20408 27678 20420
rect 27709 20417 27721 20420
rect 27755 20417 27767 20451
rect 27709 20411 27767 20417
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20448 27951 20451
rect 28813 20451 28871 20457
rect 27939 20420 28028 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 28000 20392 28028 20420
rect 28813 20417 28825 20451
rect 28859 20417 28871 20451
rect 28813 20411 28871 20417
rect 28905 20451 28963 20457
rect 28905 20417 28917 20451
rect 28951 20417 28963 20451
rect 28905 20411 28963 20417
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20349 27491 20383
rect 27433 20343 27491 20349
rect 27065 20315 27123 20321
rect 27065 20312 27077 20315
rect 26344 20284 27077 20312
rect 26237 20275 26295 20281
rect 27065 20281 27077 20284
rect 27111 20281 27123 20315
rect 27065 20275 27123 20281
rect 23624 20216 23980 20244
rect 24489 20247 24547 20253
rect 23624 20204 23630 20216
rect 24489 20213 24501 20247
rect 24535 20244 24547 20247
rect 24762 20244 24768 20256
rect 24535 20216 24768 20244
rect 24535 20213 24547 20216
rect 24489 20207 24547 20213
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 25038 20204 25044 20256
rect 25096 20204 25102 20256
rect 26252 20244 26280 20275
rect 27448 20256 27476 20343
rect 27982 20340 27988 20392
rect 28040 20340 28046 20392
rect 28920 20380 28948 20411
rect 28994 20408 29000 20460
rect 29052 20408 29058 20460
rect 29086 20408 29092 20460
rect 29144 20408 29150 20460
rect 29196 20457 29224 20488
rect 30116 20460 30144 20488
rect 30929 20485 30941 20519
rect 30975 20485 30987 20519
rect 30929 20479 30987 20485
rect 31159 20519 31217 20525
rect 31159 20485 31171 20519
rect 31205 20516 31217 20519
rect 32600 20516 32628 20547
rect 31205 20488 32628 20516
rect 31205 20485 31217 20488
rect 31159 20479 31217 20485
rect 29181 20451 29239 20457
rect 29181 20417 29193 20451
rect 29227 20417 29239 20451
rect 29181 20411 29239 20417
rect 29270 20408 29276 20460
rect 29328 20408 29334 20460
rect 29914 20408 29920 20460
rect 29972 20408 29978 20460
rect 30006 20408 30012 20460
rect 30064 20408 30070 20460
rect 30098 20408 30104 20460
rect 30156 20408 30162 20460
rect 30834 20408 30840 20460
rect 30892 20408 30898 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 30024 20380 30052 20408
rect 31036 20380 31064 20411
rect 31294 20408 31300 20460
rect 31352 20408 31358 20460
rect 31386 20408 31392 20460
rect 31444 20408 31450 20460
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 32953 20451 33011 20457
rect 32953 20417 32965 20451
rect 32999 20448 33011 20451
rect 33134 20448 33140 20460
rect 32999 20420 33140 20448
rect 32999 20417 33011 20420
rect 32953 20411 33011 20417
rect 28920 20352 29684 20380
rect 30024 20352 31064 20380
rect 29656 20256 29684 20352
rect 30282 20272 30288 20324
rect 30340 20312 30346 20324
rect 31588 20312 31616 20411
rect 33134 20408 33140 20420
rect 33192 20448 33198 20460
rect 33686 20448 33692 20460
rect 33192 20420 33692 20448
rect 33192 20408 33198 20420
rect 33686 20408 33692 20420
rect 33744 20448 33750 20460
rect 34330 20448 34336 20460
rect 33744 20420 34336 20448
rect 33744 20408 33750 20420
rect 34330 20408 34336 20420
rect 34388 20408 34394 20460
rect 33045 20383 33103 20389
rect 33045 20349 33057 20383
rect 33091 20349 33103 20383
rect 33045 20343 33103 20349
rect 30340 20284 31616 20312
rect 30340 20272 30346 20284
rect 32950 20272 32956 20324
rect 33008 20312 33014 20324
rect 33060 20312 33088 20343
rect 33008 20284 33088 20312
rect 33008 20272 33014 20284
rect 26786 20244 26792 20256
rect 26252 20216 26792 20244
rect 26786 20204 26792 20216
rect 26844 20204 26850 20256
rect 26970 20204 26976 20256
rect 27028 20204 27034 20256
rect 27430 20204 27436 20256
rect 27488 20204 27494 20256
rect 29638 20204 29644 20256
rect 29696 20204 29702 20256
rect 29730 20204 29736 20256
rect 29788 20204 29794 20256
rect 30466 20204 30472 20256
rect 30524 20244 30530 20256
rect 30653 20247 30711 20253
rect 30653 20244 30665 20247
rect 30524 20216 30665 20244
rect 30524 20204 30530 20216
rect 30653 20213 30665 20216
rect 30699 20213 30711 20247
rect 30653 20207 30711 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 13998 20000 14004 20052
rect 14056 20000 14062 20052
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 14642 20040 14648 20052
rect 14599 20012 14648 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 17862 20040 17868 20052
rect 15252 20012 17868 20040
rect 15252 20000 15258 20012
rect 17862 20000 17868 20012
rect 17920 20040 17926 20052
rect 17957 20043 18015 20049
rect 17957 20040 17969 20043
rect 17920 20012 17969 20040
rect 17920 20000 17926 20012
rect 17957 20009 17969 20012
rect 18003 20009 18015 20043
rect 20990 20040 20996 20052
rect 17957 20003 18015 20009
rect 18064 20012 20996 20040
rect 11974 19932 11980 19984
rect 12032 19932 12038 19984
rect 12618 19972 12624 19984
rect 12452 19944 12624 19972
rect 9217 19907 9275 19913
rect 9217 19873 9229 19907
rect 9263 19904 9275 19907
rect 9306 19904 9312 19916
rect 9263 19876 9312 19904
rect 9263 19873 9275 19876
rect 9217 19867 9275 19873
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8352 19808 8953 19836
rect 8352 19796 8358 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19836 10839 19839
rect 10962 19836 10968 19848
rect 10827 19808 10968 19836
rect 10827 19805 10839 19808
rect 10781 19799 10839 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 9858 19728 9864 19780
rect 9916 19728 9922 19780
rect 11072 19768 11100 19799
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 12452 19836 12480 19944
rect 12618 19932 12624 19944
rect 12676 19972 12682 19984
rect 13906 19972 13912 19984
rect 12676 19944 13912 19972
rect 12676 19932 12682 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 14016 19972 14044 20000
rect 15381 19975 15439 19981
rect 15381 19972 15393 19975
rect 14016 19944 15393 19972
rect 15381 19941 15393 19944
rect 15427 19941 15439 19975
rect 15381 19935 15439 19941
rect 17586 19932 17592 19984
rect 17644 19972 17650 19984
rect 18064 19972 18092 20012
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 23293 20043 23351 20049
rect 23293 20009 23305 20043
rect 23339 20040 23351 20043
rect 23474 20040 23480 20052
rect 23339 20012 23480 20040
rect 23339 20009 23351 20012
rect 23293 20003 23351 20009
rect 23474 20000 23480 20012
rect 23532 20000 23538 20052
rect 25038 20000 25044 20052
rect 25096 20000 25102 20052
rect 29638 20000 29644 20052
rect 29696 20040 29702 20052
rect 29733 20043 29791 20049
rect 29733 20040 29745 20043
rect 29696 20012 29745 20040
rect 29696 20000 29702 20012
rect 29733 20009 29745 20012
rect 29779 20009 29791 20043
rect 29733 20003 29791 20009
rect 17644 19944 18092 19972
rect 17644 19932 17650 19944
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 23109 19975 23167 19981
rect 23109 19972 23121 19975
rect 22152 19944 23121 19972
rect 22152 19932 22158 19944
rect 23109 19941 23121 19944
rect 23155 19941 23167 19975
rect 23109 19935 23167 19941
rect 23382 19932 23388 19984
rect 23440 19972 23446 19984
rect 24854 19972 24860 19984
rect 23440 19944 24860 19972
rect 23440 19932 23446 19944
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 12526 19864 12532 19916
rect 12584 19864 12590 19916
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19904 13139 19907
rect 13354 19904 13360 19916
rect 13127 19876 13360 19904
rect 13127 19873 13139 19876
rect 13081 19867 13139 19873
rect 13354 19864 13360 19876
rect 13412 19904 13418 19916
rect 14182 19904 14188 19916
rect 13412 19876 14188 19904
rect 13412 19864 13418 19876
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 14369 19907 14427 19913
rect 14369 19873 14381 19907
rect 14415 19904 14427 19907
rect 14829 19907 14887 19913
rect 14829 19904 14841 19907
rect 14415 19876 14841 19904
rect 14415 19873 14427 19876
rect 14369 19867 14427 19873
rect 14829 19873 14841 19876
rect 14875 19873 14887 19907
rect 17604 19904 17632 19932
rect 14829 19867 14887 19873
rect 15764 19876 17632 19904
rect 11940 19808 12480 19836
rect 11940 19796 11946 19808
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12768 19808 13018 19836
rect 12768 19796 12774 19808
rect 13722 19796 13728 19848
rect 13780 19796 13786 19848
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 14734 19796 14740 19848
rect 14792 19796 14798 19848
rect 14918 19796 14924 19848
rect 14976 19796 14982 19848
rect 15562 19796 15568 19848
rect 15620 19796 15626 19848
rect 15764 19845 15792 19876
rect 18966 19864 18972 19916
rect 19024 19864 19030 19916
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 24762 19864 24768 19916
rect 24820 19864 24826 19916
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 15838 19796 15844 19848
rect 15896 19845 15902 19848
rect 15896 19839 15925 19845
rect 15913 19805 15925 19839
rect 15896 19799 15925 19805
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19836 16083 19839
rect 16114 19836 16120 19848
rect 16071 19808 16120 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 15896 19796 15902 19799
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 17770 19796 17776 19848
rect 17828 19836 17834 19848
rect 18414 19836 18420 19848
rect 17828 19808 18420 19836
rect 17828 19796 17834 19808
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18616 19808 18705 19836
rect 10612 19740 11100 19768
rect 12345 19771 12403 19777
rect 9950 19660 9956 19712
rect 10008 19700 10014 19712
rect 10612 19700 10640 19740
rect 12345 19737 12357 19771
rect 12391 19768 12403 19771
rect 13740 19768 13768 19796
rect 12391 19740 13768 19768
rect 13909 19771 13967 19777
rect 12391 19737 12403 19740
rect 12345 19731 12403 19737
rect 13909 19737 13921 19771
rect 13955 19768 13967 19771
rect 15378 19768 15384 19780
rect 13955 19740 15384 19768
rect 13955 19737 13967 19740
rect 13909 19731 13967 19737
rect 15378 19728 15384 19740
rect 15436 19728 15442 19780
rect 15657 19771 15715 19777
rect 15657 19737 15669 19771
rect 15703 19737 15715 19771
rect 15657 19731 15715 19737
rect 10008 19672 10640 19700
rect 10008 19660 10014 19672
rect 10686 19660 10692 19712
rect 10744 19700 10750 19712
rect 11698 19700 11704 19712
rect 10744 19672 11704 19700
rect 10744 19660 10750 19672
rect 11698 19660 11704 19672
rect 11756 19700 11762 19712
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 11756 19672 12449 19700
rect 11756 19660 11762 19672
rect 12437 19669 12449 19672
rect 12483 19700 12495 19703
rect 13722 19700 13728 19712
rect 12483 19672 13728 19700
rect 12483 19669 12495 19672
rect 12437 19663 12495 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 15672 19700 15700 19731
rect 18616 19712 18644 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25056 19836 25084 20000
rect 27522 19932 27528 19984
rect 27580 19972 27586 19984
rect 29748 19972 29776 20003
rect 29914 20000 29920 20052
rect 29972 20040 29978 20052
rect 30101 20043 30159 20049
rect 30101 20040 30113 20043
rect 29972 20012 30113 20040
rect 29972 20000 29978 20012
rect 30101 20009 30113 20012
rect 30147 20009 30159 20043
rect 30101 20003 30159 20009
rect 30742 20000 30748 20052
rect 30800 20000 30806 20052
rect 30834 20000 30840 20052
rect 30892 20040 30898 20052
rect 31113 20043 31171 20049
rect 31113 20040 31125 20043
rect 30892 20012 31125 20040
rect 30892 20000 30898 20012
rect 31113 20009 31125 20012
rect 31159 20009 31171 20043
rect 33134 20040 33140 20052
rect 31113 20003 31171 20009
rect 32692 20012 33140 20040
rect 30760 19972 30788 20000
rect 27580 19944 27936 19972
rect 29748 19944 30788 19972
rect 27580 19932 27586 19944
rect 27706 19904 27712 19916
rect 26160 19876 27712 19904
rect 26160 19848 26188 19876
rect 24995 19808 25084 19836
rect 25133 19839 25191 19845
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25590 19836 25596 19848
rect 25179 19808 25596 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 25590 19796 25596 19808
rect 25648 19836 25654 19848
rect 25777 19839 25835 19845
rect 25777 19836 25789 19839
rect 25648 19808 25789 19836
rect 25648 19796 25654 19808
rect 25777 19805 25789 19808
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 26142 19796 26148 19848
rect 26200 19796 26206 19848
rect 26326 19796 26332 19848
rect 26384 19796 26390 19848
rect 26786 19796 26792 19848
rect 26844 19796 26850 19848
rect 26896 19845 26924 19876
rect 27706 19864 27712 19876
rect 27764 19864 27770 19916
rect 27908 19904 27936 19944
rect 30653 19907 30711 19913
rect 30653 19904 30665 19907
rect 27908 19876 30665 19904
rect 30653 19873 30665 19876
rect 30699 19873 30711 19907
rect 30653 19867 30711 19873
rect 32401 19907 32459 19913
rect 32401 19873 32413 19907
rect 32447 19904 32459 19907
rect 32692 19904 32720 20012
rect 33134 20000 33140 20012
rect 33192 20000 33198 20052
rect 32447 19876 32720 19904
rect 32447 19873 32459 19876
rect 32401 19867 32459 19873
rect 32766 19864 32772 19916
rect 32824 19864 32830 19916
rect 33410 19864 33416 19916
rect 33468 19904 33474 19916
rect 33965 19907 34023 19913
rect 33965 19904 33977 19907
rect 33468 19876 33977 19904
rect 33468 19864 33474 19876
rect 33965 19873 33977 19876
rect 34011 19873 34023 19907
rect 33965 19867 34023 19873
rect 26881 19839 26939 19845
rect 26881 19805 26893 19839
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 27430 19796 27436 19848
rect 27488 19796 27494 19848
rect 27617 19839 27675 19845
rect 27617 19805 27629 19839
rect 27663 19805 27675 19839
rect 27724 19836 27752 19864
rect 27795 19839 27853 19845
rect 27795 19836 27807 19839
rect 27724 19808 27807 19836
rect 27617 19799 27675 19805
rect 27795 19805 27807 19808
rect 27841 19805 27853 19839
rect 27795 19799 27853 19805
rect 24118 19728 24124 19780
rect 24176 19768 24182 19780
rect 25685 19771 25743 19777
rect 25685 19768 25697 19771
rect 24176 19740 25697 19768
rect 24176 19728 24182 19740
rect 25685 19737 25697 19740
rect 25731 19737 25743 19771
rect 26804 19768 26832 19796
rect 27632 19768 27660 19799
rect 28442 19796 28448 19848
rect 28500 19796 28506 19848
rect 30466 19796 30472 19848
rect 30524 19796 30530 19848
rect 31021 19839 31079 19845
rect 31021 19805 31033 19839
rect 31067 19805 31079 19839
rect 31021 19799 31079 19805
rect 31205 19839 31263 19845
rect 31205 19805 31217 19839
rect 31251 19836 31263 19839
rect 31386 19836 31392 19848
rect 31251 19808 31392 19836
rect 31251 19805 31263 19808
rect 31205 19799 31263 19805
rect 28460 19768 28488 19796
rect 26804 19740 28488 19768
rect 25685 19731 25743 19737
rect 28994 19728 29000 19780
rect 29052 19768 29058 19780
rect 29549 19771 29607 19777
rect 29549 19768 29561 19771
rect 29052 19740 29561 19768
rect 29052 19728 29058 19740
rect 29549 19737 29561 19740
rect 29595 19768 29607 19771
rect 29638 19768 29644 19780
rect 29595 19740 29644 19768
rect 29595 19737 29607 19740
rect 29549 19731 29607 19737
rect 29638 19728 29644 19740
rect 29696 19728 29702 19780
rect 30282 19768 30288 19780
rect 29932 19740 30288 19768
rect 16298 19700 16304 19712
rect 15672 19672 16304 19700
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 18598 19660 18604 19712
rect 18656 19660 18662 19712
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 27062 19700 27068 19712
rect 19668 19672 27068 19700
rect 19668 19660 19674 19672
rect 27062 19660 27068 19672
rect 27120 19660 27126 19712
rect 27706 19660 27712 19712
rect 27764 19660 27770 19712
rect 29086 19660 29092 19712
rect 29144 19700 29150 19712
rect 29932 19709 29960 19740
rect 30282 19728 30288 19740
rect 30340 19768 30346 19780
rect 31036 19768 31064 19799
rect 31386 19796 31392 19808
rect 31444 19836 31450 19848
rect 31849 19839 31907 19845
rect 31444 19808 31754 19836
rect 31444 19796 31450 19808
rect 30340 19740 31064 19768
rect 30340 19728 30346 19740
rect 29749 19703 29807 19709
rect 29749 19700 29761 19703
rect 29144 19672 29761 19700
rect 29144 19660 29150 19672
rect 29749 19669 29761 19672
rect 29795 19669 29807 19703
rect 29749 19663 29807 19669
rect 29917 19703 29975 19709
rect 29917 19669 29929 19703
rect 29963 19669 29975 19703
rect 29917 19663 29975 19669
rect 30561 19703 30619 19709
rect 30561 19669 30573 19703
rect 30607 19700 30619 19703
rect 31018 19700 31024 19712
rect 30607 19672 31024 19700
rect 30607 19669 30619 19672
rect 30561 19663 30619 19669
rect 31018 19660 31024 19672
rect 31076 19660 31082 19712
rect 31726 19700 31754 19808
rect 31849 19805 31861 19839
rect 31895 19805 31907 19839
rect 31849 19799 31907 19805
rect 31864 19768 31892 19799
rect 32030 19796 32036 19848
rect 32088 19796 32094 19848
rect 32214 19796 32220 19848
rect 32272 19836 32278 19848
rect 32309 19839 32367 19845
rect 32309 19836 32321 19839
rect 32272 19808 32321 19836
rect 32272 19796 32278 19808
rect 32309 19805 32321 19808
rect 32355 19836 32367 19839
rect 33042 19836 33048 19848
rect 32355 19830 32720 19836
rect 32876 19830 33048 19836
rect 32355 19808 33048 19830
rect 32355 19805 32367 19808
rect 32309 19799 32367 19805
rect 32692 19802 32904 19808
rect 33042 19796 33048 19808
rect 33100 19796 33106 19848
rect 33873 19839 33931 19845
rect 33873 19836 33885 19839
rect 33336 19808 33885 19836
rect 32398 19768 32404 19780
rect 31864 19740 32404 19768
rect 32398 19728 32404 19740
rect 32456 19768 32462 19780
rect 32582 19768 32588 19780
rect 32456 19740 32588 19768
rect 32456 19728 32462 19740
rect 32582 19728 32588 19740
rect 32640 19728 32646 19780
rect 31849 19703 31907 19709
rect 31849 19700 31861 19703
rect 31726 19672 31861 19700
rect 31849 19669 31861 19672
rect 31895 19669 31907 19703
rect 31849 19663 31907 19669
rect 32677 19703 32735 19709
rect 32677 19669 32689 19703
rect 32723 19700 32735 19703
rect 33336 19700 33364 19808
rect 33873 19805 33885 19808
rect 33919 19805 33931 19839
rect 33873 19799 33931 19805
rect 35526 19768 35532 19780
rect 33796 19740 35532 19768
rect 33796 19712 33824 19740
rect 35526 19728 35532 19740
rect 35584 19728 35590 19780
rect 32723 19672 33364 19700
rect 32723 19669 32735 19672
rect 32677 19663 32735 19669
rect 33778 19660 33784 19712
rect 33836 19660 33842 19712
rect 1104 19610 38824 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 38824 19610
rect 1104 19536 38824 19558
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 9861 19499 9919 19505
rect 9861 19496 9873 19499
rect 4120 19468 9873 19496
rect 4120 19456 4126 19468
rect 9861 19465 9873 19468
rect 9907 19496 9919 19499
rect 9950 19496 9956 19508
rect 9907 19468 9956 19496
rect 9907 19465 9919 19468
rect 9861 19459 9919 19465
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 14737 19499 14795 19505
rect 14737 19496 14749 19499
rect 14332 19468 14749 19496
rect 14332 19456 14338 19468
rect 14737 19465 14749 19468
rect 14783 19465 14795 19499
rect 14737 19459 14795 19465
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 15160 19468 15500 19496
rect 15160 19456 15166 19468
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 12986 19428 12992 19440
rect 3476 19400 12992 19428
rect 3476 19388 3482 19400
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 15472 19428 15500 19468
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15620 19468 15761 19496
rect 15620 19456 15626 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 16206 19496 16212 19508
rect 15749 19459 15807 19465
rect 15948 19468 16212 19496
rect 15948 19428 15976 19468
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 16298 19456 16304 19508
rect 16356 19456 16362 19508
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 22370 19496 22376 19508
rect 19024 19468 22376 19496
rect 19024 19456 19030 19468
rect 15472 19400 15976 19428
rect 10597 19363 10655 19369
rect 10597 19329 10609 19363
rect 10643 19360 10655 19363
rect 10686 19360 10692 19372
rect 10643 19332 10692 19360
rect 10643 19329 10655 19332
rect 10597 19323 10655 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 10962 19360 10968 19372
rect 10919 19332 10968 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11204 19332 11897 19360
rect 11204 19320 11210 19332
rect 11885 19329 11897 19332
rect 11931 19360 11943 19363
rect 11931 19332 12434 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12406 19224 12434 19332
rect 13538 19320 13544 19372
rect 13596 19320 13602 19372
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 13817 19363 13875 19369
rect 13817 19360 13829 19363
rect 13780 19332 13829 19360
rect 13780 19320 13786 19332
rect 13817 19329 13829 19332
rect 13863 19329 13875 19363
rect 13817 19323 13875 19329
rect 14016 19332 14228 19360
rect 13556 19292 13584 19320
rect 14016 19292 14044 19332
rect 13556 19264 14044 19292
rect 14090 19252 14096 19304
rect 14148 19252 14154 19304
rect 14200 19301 14228 19332
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 15948 19369 15976 19400
rect 16666 19388 16672 19440
rect 16724 19388 16730 19440
rect 17678 19388 17684 19440
rect 17736 19428 17742 19440
rect 20809 19431 20867 19437
rect 17736 19400 20760 19428
rect 17736 19388 17742 19400
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14516 19332 14933 19360
rect 14516 19320 14522 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15194 19363 15252 19369
rect 15194 19329 15206 19363
rect 15240 19329 15252 19363
rect 15194 19323 15252 19329
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16117 19366 16175 19369
rect 16209 19366 16267 19369
rect 16117 19363 16267 19366
rect 16117 19329 16129 19363
rect 16163 19338 16221 19363
rect 16163 19329 16175 19338
rect 16117 19323 16175 19329
rect 16209 19329 16221 19338
rect 16255 19360 16267 19363
rect 16255 19332 16309 19360
rect 16255 19329 16267 19332
rect 16209 19323 16267 19329
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19261 14243 19295
rect 15212 19292 15240 19323
rect 15470 19292 15476 19304
rect 15212 19264 15476 19292
rect 14185 19255 14243 19261
rect 15470 19252 15476 19264
rect 15528 19292 15534 19304
rect 16224 19292 16252 19323
rect 16390 19320 16396 19372
rect 16448 19360 16454 19372
rect 18506 19360 18512 19372
rect 16448 19332 18512 19360
rect 16448 19320 16454 19332
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20622 19360 20628 19372
rect 19935 19332 20628 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20732 19360 20760 19400
rect 20809 19397 20821 19431
rect 20855 19428 20867 19431
rect 20898 19428 20904 19440
rect 20855 19400 20904 19428
rect 20855 19397 20867 19400
rect 20809 19391 20867 19397
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 21836 19372 21864 19468
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24213 19499 24271 19505
rect 24213 19496 24225 19499
rect 24084 19468 24225 19496
rect 24084 19456 24090 19468
rect 24213 19465 24225 19468
rect 24259 19465 24271 19499
rect 24213 19459 24271 19465
rect 25682 19456 25688 19508
rect 25740 19456 25746 19508
rect 29730 19496 29736 19508
rect 29564 19468 29736 19496
rect 24305 19431 24363 19437
rect 24305 19428 24317 19431
rect 23584 19400 24317 19428
rect 20732 19332 21220 19360
rect 21192 19304 21220 19332
rect 21818 19320 21824 19372
rect 21876 19320 21882 19372
rect 22094 19320 22100 19372
rect 22152 19320 22158 19372
rect 22830 19320 22836 19372
rect 22888 19360 22894 19372
rect 23584 19369 23612 19400
rect 24305 19397 24317 19400
rect 24351 19397 24363 19431
rect 29454 19428 29460 19440
rect 24305 19391 24363 19397
rect 29288 19400 29460 19428
rect 23569 19363 23627 19369
rect 23569 19360 23581 19363
rect 22888 19332 23581 19360
rect 22888 19320 22894 19332
rect 23569 19329 23581 19332
rect 23615 19329 23627 19363
rect 23569 19323 23627 19329
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 23934 19360 23940 19372
rect 23799 19332 23940 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 23934 19320 23940 19332
rect 23992 19320 23998 19372
rect 24118 19320 24124 19372
rect 24176 19360 24182 19372
rect 24176 19332 24624 19360
rect 24176 19320 24182 19332
rect 15528 19264 16252 19292
rect 15528 19252 15534 19264
rect 21174 19252 21180 19304
rect 21232 19252 21238 19304
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19292 23535 19295
rect 23661 19295 23719 19301
rect 23523 19264 23612 19292
rect 23523 19261 23535 19264
rect 23477 19255 23535 19261
rect 17957 19227 18015 19233
rect 17957 19224 17969 19227
rect 12406 19196 17969 19224
rect 17957 19193 17969 19196
rect 18003 19224 18015 19227
rect 19242 19224 19248 19236
rect 18003 19196 19248 19224
rect 18003 19193 18015 19196
rect 17957 19187 18015 19193
rect 19242 19184 19248 19196
rect 19300 19224 19306 19236
rect 23584 19224 23612 19264
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 24026 19292 24032 19304
rect 23707 19264 24032 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 24026 19252 24032 19264
rect 24084 19292 24090 19304
rect 24489 19295 24547 19301
rect 24489 19292 24501 19295
rect 24084 19264 24501 19292
rect 24084 19252 24090 19264
rect 24489 19261 24501 19264
rect 24535 19261 24547 19295
rect 24489 19255 24547 19261
rect 24596 19292 24624 19332
rect 25314 19320 25320 19372
rect 25372 19320 25378 19372
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 25501 19363 25559 19369
rect 25501 19360 25513 19363
rect 25464 19332 25513 19360
rect 25464 19320 25470 19332
rect 25501 19329 25513 19332
rect 25547 19329 25559 19363
rect 25501 19323 25559 19329
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 29288 19369 29316 19400
rect 29454 19388 29460 19400
rect 29512 19388 29518 19440
rect 29564 19437 29592 19468
rect 29730 19456 29736 19468
rect 29788 19456 29794 19508
rect 31018 19456 31024 19508
rect 31076 19496 31082 19508
rect 31076 19468 31754 19496
rect 31076 19456 31082 19468
rect 29549 19431 29607 19437
rect 29549 19397 29561 19431
rect 29595 19397 29607 19431
rect 29549 19391 29607 19397
rect 30558 19388 30564 19440
rect 30616 19388 30622 19440
rect 31726 19428 31754 19468
rect 32030 19456 32036 19508
rect 32088 19496 32094 19508
rect 32493 19499 32551 19505
rect 32493 19496 32505 19499
rect 32088 19468 32505 19496
rect 32088 19456 32094 19468
rect 32493 19465 32505 19468
rect 32539 19465 32551 19499
rect 32493 19459 32551 19465
rect 32582 19456 32588 19508
rect 32640 19496 32646 19508
rect 32953 19499 33011 19505
rect 32953 19496 32965 19499
rect 32640 19468 32965 19496
rect 32640 19456 32646 19468
rect 32953 19465 32965 19468
rect 32999 19465 33011 19499
rect 32953 19459 33011 19465
rect 33410 19456 33416 19508
rect 33468 19456 33474 19508
rect 33778 19456 33784 19508
rect 33836 19456 33842 19508
rect 34330 19456 34336 19508
rect 34388 19456 34394 19508
rect 32214 19428 32220 19440
rect 31726 19400 32220 19428
rect 32214 19388 32220 19400
rect 32272 19388 32278 19440
rect 32861 19431 32919 19437
rect 32861 19397 32873 19431
rect 32907 19428 32919 19431
rect 33428 19428 33456 19456
rect 32907 19400 33456 19428
rect 32907 19397 32919 19400
rect 32861 19391 32919 19397
rect 27249 19363 27307 19369
rect 27249 19360 27261 19363
rect 27028 19332 27261 19360
rect 27028 19320 27034 19332
rect 27249 19329 27261 19332
rect 27295 19329 27307 19363
rect 27249 19323 27307 19329
rect 29273 19363 29331 19369
rect 29273 19329 29285 19363
rect 29319 19329 29331 19363
rect 29273 19323 29331 19329
rect 32677 19363 32735 19369
rect 32677 19329 32689 19363
rect 32723 19360 32735 19363
rect 32950 19360 32956 19372
rect 32723 19332 32956 19360
rect 32723 19329 32735 19332
rect 32677 19323 32735 19329
rect 32950 19320 32956 19332
rect 33008 19320 33014 19372
rect 33152 19369 33180 19400
rect 33137 19363 33195 19369
rect 33137 19329 33149 19363
rect 33183 19329 33195 19363
rect 33137 19323 33195 19329
rect 33597 19363 33655 19369
rect 33597 19329 33609 19363
rect 33643 19360 33655 19363
rect 33796 19360 33824 19456
rect 33643 19332 33824 19360
rect 33643 19329 33655 19332
rect 33597 19323 33655 19329
rect 25866 19292 25872 19304
rect 24596 19264 25872 19292
rect 24596 19224 24624 19264
rect 25866 19252 25872 19264
rect 25924 19252 25930 19304
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19292 27399 19295
rect 27706 19292 27712 19304
rect 27387 19264 27712 19292
rect 27387 19261 27399 19264
rect 27341 19255 27399 19261
rect 27706 19252 27712 19264
rect 27764 19252 27770 19304
rect 33318 19252 33324 19304
rect 33376 19252 33382 19304
rect 19300 19196 21036 19224
rect 19300 19184 19306 19196
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 13630 19156 13636 19168
rect 13403 19128 13636 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18601 19159 18659 19165
rect 18601 19156 18613 19159
rect 18196 19128 18613 19156
rect 18196 19116 18202 19128
rect 18601 19125 18613 19128
rect 18647 19125 18659 19159
rect 18601 19119 18659 19125
rect 20073 19159 20131 19165
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 20530 19156 20536 19168
rect 20119 19128 20536 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 20901 19159 20959 19165
rect 20901 19156 20913 19159
rect 20864 19128 20913 19156
rect 20864 19116 20870 19128
rect 20901 19125 20913 19128
rect 20947 19125 20959 19159
rect 21008 19156 21036 19196
rect 22756 19196 23520 19224
rect 23584 19196 24624 19224
rect 22756 19156 22784 19196
rect 21008 19128 22784 19156
rect 22833 19159 22891 19165
rect 20901 19119 20959 19125
rect 22833 19125 22845 19159
rect 22879 19156 22891 19159
rect 23198 19156 23204 19168
rect 22879 19128 23204 19156
rect 22879 19125 22891 19128
rect 22833 19119 22891 19125
rect 23198 19116 23204 19128
rect 23256 19116 23262 19168
rect 23290 19116 23296 19168
rect 23348 19116 23354 19168
rect 23492 19156 23520 19196
rect 23566 19156 23572 19168
rect 23492 19128 23572 19156
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 23934 19116 23940 19168
rect 23992 19116 23998 19168
rect 27522 19116 27528 19168
rect 27580 19116 27586 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 10870 18952 10876 18964
rect 10520 18924 10876 18952
rect 10520 18825 10548 18924
rect 10870 18912 10876 18924
rect 10928 18912 10934 18964
rect 13170 18952 13176 18964
rect 12406 18924 13176 18952
rect 10505 18819 10563 18825
rect 10505 18785 10517 18819
rect 10551 18785 10563 18819
rect 10505 18779 10563 18785
rect 12158 18776 12164 18828
rect 12216 18776 12222 18828
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 10796 18680 10824 18711
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 12253 18751 12311 18757
rect 12253 18748 12265 18751
rect 11664 18720 12265 18748
rect 11664 18708 11670 18720
rect 12253 18717 12265 18720
rect 12299 18748 12311 18751
rect 12406 18748 12434 18924
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13262 18912 13268 18964
rect 13320 18952 13326 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13320 18924 13553 18952
rect 13320 18912 13326 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 13541 18915 13599 18921
rect 17954 18912 17960 18964
rect 18012 18912 18018 18964
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18506 18952 18512 18964
rect 18187 18924 18512 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 20622 18912 20628 18964
rect 20680 18952 20686 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 20680 18924 21465 18952
rect 20680 18912 20686 18924
rect 21453 18921 21465 18924
rect 21499 18952 21511 18955
rect 22462 18952 22468 18964
rect 21499 18924 22468 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 22830 18912 22836 18964
rect 22888 18952 22894 18964
rect 22925 18955 22983 18961
rect 22925 18952 22937 18955
rect 22888 18924 22937 18952
rect 22888 18912 22894 18924
rect 22925 18921 22937 18924
rect 22971 18921 22983 18955
rect 22925 18915 22983 18921
rect 23753 18955 23811 18961
rect 23753 18921 23765 18955
rect 23799 18952 23811 18955
rect 23842 18952 23848 18964
rect 23799 18924 23848 18952
rect 23799 18921 23811 18924
rect 23753 18915 23811 18921
rect 12621 18887 12679 18893
rect 12621 18853 12633 18887
rect 12667 18884 12679 18887
rect 14550 18884 14556 18896
rect 12667 18856 14556 18884
rect 12667 18853 12679 18856
rect 12621 18847 12679 18853
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 19150 18884 19156 18896
rect 16960 18856 19156 18884
rect 12710 18776 12716 18828
rect 12768 18776 12774 18828
rect 13078 18776 13084 18828
rect 13136 18776 13142 18828
rect 13198 18819 13256 18825
rect 13198 18785 13210 18819
rect 13244 18816 13256 18819
rect 13354 18816 13360 18828
rect 13244 18788 13360 18816
rect 13244 18785 13256 18788
rect 13198 18779 13256 18785
rect 13354 18776 13360 18788
rect 13412 18816 13418 18828
rect 13412 18788 13676 18816
rect 13412 18776 13418 18788
rect 13538 18748 13544 18760
rect 12299 18720 12434 18748
rect 13004 18720 13544 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 13004 18692 13032 18720
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 13648 18757 13676 18788
rect 14734 18776 14740 18828
rect 14792 18776 14798 18828
rect 15197 18819 15255 18825
rect 15197 18785 15209 18819
rect 15243 18816 15255 18819
rect 15289 18819 15347 18825
rect 15289 18816 15301 18819
rect 15243 18788 15301 18816
rect 15243 18785 15255 18788
rect 15197 18779 15255 18785
rect 15289 18785 15301 18788
rect 15335 18816 15347 18819
rect 15470 18816 15476 18828
rect 15335 18788 15476 18816
rect 15335 18785 15347 18788
rect 15289 18779 15347 18785
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 16960 18825 16988 18856
rect 19150 18844 19156 18856
rect 19208 18844 19214 18896
rect 16945 18819 17003 18825
rect 16945 18785 16957 18819
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 18693 18819 18751 18825
rect 18693 18785 18705 18819
rect 18739 18816 18751 18819
rect 19702 18816 19708 18828
rect 18739 18788 19708 18816
rect 18739 18785 18751 18788
rect 18693 18779 18751 18785
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 14369 18751 14427 18757
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14458 18748 14464 18760
rect 14415 18720 14464 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 14458 18708 14464 18720
rect 14516 18708 14522 18760
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18748 14703 18751
rect 14752 18748 14780 18776
rect 14691 18720 14780 18748
rect 14921 18751 14979 18757
rect 14691 18717 14703 18720
rect 14645 18711 14703 18717
rect 14921 18717 14933 18751
rect 14967 18748 14979 18751
rect 15102 18748 15108 18760
rect 14967 18720 15108 18748
rect 14967 18717 14979 18720
rect 14921 18711 14979 18717
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15436 18720 15945 18748
rect 15436 18708 15442 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 16114 18708 16120 18760
rect 16172 18708 16178 18760
rect 16298 18708 16304 18760
rect 16356 18708 16362 18760
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16816 18720 16865 18748
rect 16816 18708 16822 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 16853 18711 16911 18717
rect 17144 18720 17325 18748
rect 9876 18652 10824 18680
rect 9876 18624 9904 18652
rect 12986 18640 12992 18692
rect 13044 18640 13050 18692
rect 16132 18680 16160 18708
rect 17144 18680 17172 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17586 18708 17592 18760
rect 17644 18708 17650 18760
rect 17770 18708 17776 18760
rect 17828 18708 17834 18760
rect 18138 18708 18144 18760
rect 18196 18708 18202 18760
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 18248 18720 18337 18748
rect 17451 18683 17509 18689
rect 17451 18680 17463 18683
rect 13372 18652 14964 18680
rect 16132 18652 17172 18680
rect 17236 18652 17463 18680
rect 9858 18572 9864 18624
rect 9916 18572 9922 18624
rect 13372 18621 13400 18652
rect 14936 18624 14964 18652
rect 13357 18615 13415 18621
rect 13357 18581 13369 18615
rect 13403 18581 13415 18615
rect 13357 18575 13415 18581
rect 14642 18572 14648 18624
rect 14700 18572 14706 18624
rect 14918 18572 14924 18624
rect 14976 18572 14982 18624
rect 17236 18621 17264 18652
rect 17451 18649 17463 18652
rect 17497 18649 17509 18683
rect 17451 18643 17509 18649
rect 17681 18683 17739 18689
rect 17681 18649 17693 18683
rect 17727 18680 17739 18683
rect 18156 18680 18184 18708
rect 17727 18652 18184 18680
rect 17727 18649 17739 18652
rect 17681 18643 17739 18649
rect 17221 18615 17279 18621
rect 17221 18581 17233 18615
rect 17267 18581 17279 18615
rect 17221 18575 17279 18581
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 18248 18612 18276 18720
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18432 18680 18460 18711
rect 18340 18652 18460 18680
rect 18340 18624 18368 18652
rect 18616 18624 18644 18779
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 20714 18776 20720 18828
rect 20772 18816 20778 18828
rect 20993 18819 21051 18825
rect 20993 18816 21005 18819
rect 20772 18788 21005 18816
rect 20772 18776 20778 18788
rect 20993 18785 21005 18788
rect 21039 18785 21051 18819
rect 20993 18779 21051 18785
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 21876 18788 21925 18816
rect 21876 18776 21882 18788
rect 21913 18785 21925 18788
rect 21959 18785 21971 18819
rect 22940 18816 22968 18915
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 24026 18912 24032 18964
rect 24084 18912 24090 18964
rect 24949 18955 25007 18961
rect 24949 18921 24961 18955
rect 24995 18952 25007 18955
rect 25406 18952 25412 18964
rect 24995 18924 25412 18952
rect 24995 18921 25007 18924
rect 24949 18915 25007 18921
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 28718 18952 28724 18964
rect 28679 18924 28724 18952
rect 28718 18912 28724 18924
rect 28776 18952 28782 18964
rect 30006 18952 30012 18964
rect 28776 18924 30012 18952
rect 28776 18912 28782 18924
rect 30006 18912 30012 18924
rect 30064 18912 30070 18964
rect 30285 18955 30343 18961
rect 30285 18921 30297 18955
rect 30331 18952 30343 18955
rect 30558 18952 30564 18964
rect 30331 18924 30564 18952
rect 30331 18921 30343 18924
rect 30285 18915 30343 18921
rect 30558 18912 30564 18924
rect 30616 18912 30622 18964
rect 23937 18887 23995 18893
rect 23937 18884 23949 18887
rect 23492 18856 23949 18884
rect 23492 18825 23520 18856
rect 23937 18853 23949 18856
rect 23983 18853 23995 18887
rect 23937 18847 23995 18853
rect 24044 18884 24072 18912
rect 24854 18884 24860 18896
rect 24044 18856 24860 18884
rect 23477 18819 23535 18825
rect 22940 18788 23428 18816
rect 21913 18779 21971 18785
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18840 18720 18889 18748
rect 18840 18708 18846 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 18877 18711 18935 18717
rect 21100 18720 21649 18748
rect 18969 18683 19027 18689
rect 18969 18649 18981 18683
rect 19015 18680 19027 18683
rect 19015 18652 19550 18680
rect 19015 18649 19027 18652
rect 18969 18643 19027 18649
rect 20438 18640 20444 18692
rect 20496 18680 20502 18692
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 20496 18652 20729 18680
rect 20496 18640 20502 18652
rect 20717 18649 20729 18652
rect 20763 18649 20775 18683
rect 21100 18680 21128 18720
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18748 22247 18751
rect 23198 18748 23204 18760
rect 22235 18720 23204 18748
rect 22235 18717 22247 18720
rect 22189 18711 22247 18717
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 23400 18757 23428 18788
rect 23477 18785 23489 18819
rect 23523 18785 23535 18819
rect 24044 18816 24072 18856
rect 24854 18844 24860 18856
rect 24912 18884 24918 18896
rect 25041 18887 25099 18893
rect 25041 18884 25053 18887
rect 24912 18856 25053 18884
rect 24912 18844 24918 18856
rect 25041 18853 25053 18856
rect 25087 18853 25099 18887
rect 25041 18847 25099 18853
rect 26050 18844 26056 18896
rect 26108 18884 26114 18896
rect 35434 18884 35440 18896
rect 26108 18856 27660 18884
rect 26108 18844 26114 18856
rect 23477 18779 23535 18785
rect 23860 18788 24072 18816
rect 23860 18757 23888 18788
rect 24118 18776 24124 18828
rect 24176 18776 24182 18828
rect 27522 18776 27528 18828
rect 27580 18776 27586 18828
rect 23385 18751 23443 18757
rect 23385 18717 23397 18751
rect 23431 18717 23443 18751
rect 23385 18711 23443 18717
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 24136 18748 24164 18776
rect 26970 18748 26976 18760
rect 24075 18720 24164 18748
rect 25332 18720 26976 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 20717 18643 20775 18649
rect 20916 18652 21128 18680
rect 20916 18624 20944 18652
rect 21174 18640 21180 18692
rect 21232 18680 21238 18692
rect 21542 18680 21548 18692
rect 21232 18652 21548 18680
rect 21232 18640 21238 18652
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 25332 18680 25360 18720
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 27062 18708 27068 18760
rect 27120 18748 27126 18760
rect 27249 18751 27307 18757
rect 27249 18748 27261 18751
rect 27120 18720 27261 18748
rect 27120 18708 27126 18720
rect 27249 18717 27261 18720
rect 27295 18717 27307 18751
rect 27249 18711 27307 18717
rect 27341 18751 27399 18757
rect 27341 18717 27353 18751
rect 27387 18748 27399 18751
rect 27540 18748 27568 18776
rect 27387 18720 27568 18748
rect 27632 18748 27660 18856
rect 31726 18856 35440 18884
rect 30374 18816 30380 18828
rect 30208 18788 30380 18816
rect 28629 18751 28687 18757
rect 28629 18748 28641 18751
rect 27632 18720 28641 18748
rect 27387 18717 27399 18720
rect 27341 18711 27399 18717
rect 28629 18717 28641 18720
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 29178 18708 29184 18760
rect 29236 18748 29242 18760
rect 30208 18757 30236 18788
rect 30374 18776 30380 18788
rect 30432 18776 30438 18828
rect 30193 18751 30251 18757
rect 30193 18748 30205 18751
rect 29236 18720 30205 18748
rect 29236 18708 29242 18720
rect 30193 18717 30205 18720
rect 30239 18748 30251 18751
rect 30745 18751 30803 18757
rect 30745 18748 30757 18751
rect 30239 18720 30757 18748
rect 30239 18717 30251 18720
rect 30193 18711 30251 18717
rect 30745 18717 30757 18720
rect 30791 18717 30803 18751
rect 30745 18711 30803 18717
rect 21652 18652 22094 18680
rect 18196 18584 18276 18612
rect 18196 18572 18202 18584
rect 18322 18572 18328 18624
rect 18380 18572 18386 18624
rect 18598 18572 18604 18624
rect 18656 18612 18662 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 18656 18584 19257 18612
rect 18656 18572 18662 18584
rect 19245 18581 19257 18584
rect 19291 18612 19303 18615
rect 19426 18612 19432 18624
rect 19291 18584 19432 18612
rect 19291 18581 19303 18584
rect 19245 18575 19303 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 20898 18572 20904 18624
rect 20956 18572 20962 18624
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21652 18612 21680 18652
rect 21140 18584 21680 18612
rect 21140 18572 21146 18584
rect 21726 18572 21732 18624
rect 21784 18572 21790 18624
rect 22066 18612 22094 18652
rect 23124 18652 25360 18680
rect 23124 18612 23152 18652
rect 25406 18640 25412 18692
rect 25464 18640 25470 18692
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 27157 18683 27215 18689
rect 27157 18680 27169 18683
rect 26200 18652 27169 18680
rect 26200 18640 26206 18652
rect 27157 18649 27169 18652
rect 27203 18649 27215 18683
rect 31726 18680 31754 18856
rect 35434 18844 35440 18856
rect 35492 18844 35498 18896
rect 27157 18643 27215 18649
rect 27264 18652 31754 18680
rect 22066 18584 23152 18612
rect 23198 18572 23204 18624
rect 23256 18612 23262 18624
rect 27264 18612 27292 18652
rect 23256 18584 27292 18612
rect 23256 18572 23262 18584
rect 27522 18572 27528 18624
rect 27580 18572 27586 18624
rect 30834 18572 30840 18624
rect 30892 18572 30898 18624
rect 1104 18522 38824 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 38824 18522
rect 1104 18448 38824 18470
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 12158 18408 12164 18420
rect 11572 18380 12164 18408
rect 11572 18368 11578 18380
rect 12158 18368 12164 18380
rect 12216 18408 12222 18420
rect 14366 18408 14372 18420
rect 12216 18380 14372 18408
rect 12216 18368 12222 18380
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14516 18380 15209 18408
rect 14516 18368 14522 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 16298 18368 16304 18420
rect 16356 18408 16362 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 16356 18380 16681 18408
rect 16356 18368 16362 18380
rect 16669 18377 16681 18380
rect 16715 18408 16727 18411
rect 16715 18380 17448 18408
rect 16715 18377 16727 18380
rect 16669 18371 16727 18377
rect 9766 18300 9772 18352
rect 9824 18300 9830 18352
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 17313 18343 17371 18349
rect 17313 18340 17325 18343
rect 16816 18312 17325 18340
rect 16816 18300 16822 18312
rect 17313 18309 17325 18312
rect 17359 18309 17371 18343
rect 17313 18303 17371 18309
rect 12992 18284 13044 18290
rect 15378 18232 15384 18284
rect 15436 18232 15442 18284
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16776 18272 16804 18300
rect 15979 18244 16804 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 12992 18226 13044 18232
rect 4062 18164 4068 18216
rect 4120 18164 4126 18216
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8352 18176 8493 18204
rect 8352 18164 8358 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 12526 18164 12532 18216
rect 12584 18164 12590 18216
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 14274 18204 14280 18216
rect 13403 18176 14280 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 14274 18164 14280 18176
rect 14332 18164 14338 18216
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 15841 18207 15899 18213
rect 15841 18204 15853 18207
rect 15703 18176 15853 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 15841 18173 15853 18176
rect 15887 18173 15899 18207
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 15841 18167 15899 18173
rect 16684 18176 17141 18204
rect 4080 18068 4108 18164
rect 15565 18139 15623 18145
rect 15565 18105 15577 18139
rect 15611 18136 15623 18139
rect 16684 18136 16712 18176
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17420 18204 17448 18380
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 17865 18411 17923 18417
rect 17865 18408 17877 18411
rect 17828 18380 17877 18408
rect 17828 18368 17834 18380
rect 17865 18377 17877 18380
rect 17911 18377 17923 18411
rect 17865 18371 17923 18377
rect 19061 18411 19119 18417
rect 19061 18377 19073 18411
rect 19107 18408 19119 18411
rect 19702 18408 19708 18420
rect 19107 18380 19708 18408
rect 19107 18377 19119 18380
rect 19061 18371 19119 18377
rect 18322 18340 18328 18352
rect 17788 18312 18328 18340
rect 17788 18213 17816 18312
rect 18322 18300 18328 18312
rect 18380 18300 18386 18352
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18272 18107 18275
rect 19076 18272 19104 18371
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 20530 18368 20536 18420
rect 20588 18368 20594 18420
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 23845 18411 23903 18417
rect 23845 18408 23857 18411
rect 23716 18380 23857 18408
rect 23716 18368 23722 18380
rect 23845 18377 23857 18380
rect 23891 18377 23903 18411
rect 23845 18371 23903 18377
rect 23934 18368 23940 18420
rect 23992 18368 23998 18420
rect 25314 18368 25320 18420
rect 25372 18408 25378 18420
rect 25409 18411 25467 18417
rect 25409 18408 25421 18411
rect 25372 18380 25421 18408
rect 25372 18368 25378 18380
rect 25409 18377 25421 18380
rect 25455 18377 25467 18411
rect 25409 18371 25467 18377
rect 26142 18368 26148 18420
rect 26200 18368 26206 18420
rect 27065 18411 27123 18417
rect 27065 18377 27077 18411
rect 27111 18377 27123 18411
rect 27065 18371 27123 18377
rect 27433 18411 27491 18417
rect 27433 18377 27445 18411
rect 27479 18408 27491 18411
rect 27522 18408 27528 18420
rect 27479 18380 27528 18408
rect 27479 18377 27491 18380
rect 27433 18371 27491 18377
rect 20073 18343 20131 18349
rect 20073 18309 20085 18343
rect 20119 18340 20131 18343
rect 20441 18343 20499 18349
rect 20441 18340 20453 18343
rect 20119 18312 20453 18340
rect 20119 18309 20131 18312
rect 20073 18303 20131 18309
rect 20441 18309 20453 18312
rect 20487 18309 20499 18343
rect 20441 18303 20499 18309
rect 18095 18244 19104 18272
rect 18095 18241 18107 18244
rect 18049 18235 18107 18241
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19208 18244 20177 18272
rect 19208 18232 19214 18244
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20548 18281 20576 18368
rect 20898 18300 20904 18352
rect 20956 18300 20962 18352
rect 23308 18281 23336 18368
rect 20349 18275 20407 18281
rect 20349 18272 20361 18275
rect 20312 18244 20361 18272
rect 20312 18232 20318 18244
rect 20349 18241 20361 18244
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 17773 18207 17831 18213
rect 17420 18176 17724 18204
rect 17129 18167 17187 18173
rect 15611 18108 16712 18136
rect 15611 18105 15623 18108
rect 15565 18099 15623 18105
rect 16758 18096 16764 18148
rect 16816 18096 16822 18148
rect 17144 18136 17172 18167
rect 17402 18136 17408 18148
rect 17144 18108 17408 18136
rect 17402 18096 17408 18108
rect 17460 18136 17466 18148
rect 17589 18139 17647 18145
rect 17589 18136 17601 18139
rect 17460 18108 17601 18136
rect 17460 18096 17466 18108
rect 17589 18105 17601 18108
rect 17635 18105 17647 18139
rect 17696 18136 17724 18176
rect 17773 18173 17785 18207
rect 17819 18173 17831 18207
rect 17773 18167 17831 18173
rect 18138 18164 18144 18216
rect 18196 18164 18202 18216
rect 19518 18164 19524 18216
rect 19576 18164 19582 18216
rect 19978 18164 19984 18216
rect 20036 18204 20042 18216
rect 20036 18176 21226 18204
rect 20036 18164 20042 18176
rect 18156 18136 18184 18164
rect 21082 18136 21088 18148
rect 17696 18108 18184 18136
rect 18248 18108 21088 18136
rect 17589 18099 17647 18105
rect 9858 18068 9864 18080
rect 4080 18040 9864 18068
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18248 18068 18276 18108
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 21198 18136 21226 18176
rect 21726 18164 21732 18216
rect 21784 18204 21790 18216
rect 23569 18207 23627 18213
rect 23569 18204 23581 18207
rect 21784 18176 23581 18204
rect 21784 18164 21790 18176
rect 23569 18173 23581 18176
rect 23615 18173 23627 18207
rect 23569 18167 23627 18173
rect 23474 18136 23480 18148
rect 21198 18108 23480 18136
rect 23474 18096 23480 18108
rect 23532 18096 23538 18148
rect 23952 18136 23980 18368
rect 24854 18300 24860 18352
rect 24912 18340 24918 18352
rect 24949 18343 25007 18349
rect 24949 18340 24961 18343
rect 24912 18312 24961 18340
rect 24912 18300 24918 18312
rect 24949 18309 24961 18312
rect 24995 18340 25007 18343
rect 24995 18312 25820 18340
rect 24995 18309 25007 18312
rect 24949 18303 25007 18309
rect 25792 18281 25820 18312
rect 25777 18275 25835 18281
rect 25777 18241 25789 18275
rect 25823 18241 25835 18275
rect 25777 18235 25835 18241
rect 26789 18275 26847 18281
rect 26789 18241 26801 18275
rect 26835 18272 26847 18275
rect 27080 18272 27108 18371
rect 27522 18368 27528 18380
rect 27580 18368 27586 18420
rect 29733 18411 29791 18417
rect 29733 18377 29745 18411
rect 29779 18377 29791 18411
rect 29733 18371 29791 18377
rect 29748 18340 29776 18371
rect 30101 18343 30159 18349
rect 30101 18340 30113 18343
rect 29748 18312 30113 18340
rect 30101 18309 30113 18312
rect 30147 18309 30159 18343
rect 30101 18303 30159 18309
rect 30834 18300 30840 18352
rect 30892 18300 30898 18352
rect 26835 18244 27108 18272
rect 26835 18241 26847 18244
rect 26789 18235 26847 18241
rect 29546 18232 29552 18284
rect 29604 18232 29610 18284
rect 32490 18272 32496 18284
rect 31588 18244 32496 18272
rect 25866 18164 25872 18216
rect 25924 18164 25930 18216
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 27356 18176 27537 18204
rect 23676 18108 23980 18136
rect 16172 18040 18276 18068
rect 18325 18071 18383 18077
rect 16172 18028 16178 18040
rect 18325 18037 18337 18071
rect 18371 18068 18383 18071
rect 18598 18068 18604 18080
rect 18371 18040 18604 18068
rect 18371 18037 18383 18040
rect 18325 18031 18383 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 23676 18077 23704 18108
rect 25314 18096 25320 18148
rect 25372 18136 25378 18148
rect 27356 18136 27384 18176
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27525 18167 27583 18173
rect 27614 18164 27620 18216
rect 27672 18164 27678 18216
rect 29454 18164 29460 18216
rect 29512 18204 29518 18216
rect 29825 18207 29883 18213
rect 29825 18204 29837 18207
rect 29512 18176 29837 18204
rect 29512 18164 29518 18176
rect 29825 18173 29837 18176
rect 29871 18173 29883 18207
rect 29825 18167 29883 18173
rect 25372 18108 27384 18136
rect 25372 18096 25378 18108
rect 27356 18080 27384 18108
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20496 18040 20729 18068
rect 20496 18028 20502 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 23661 18071 23719 18077
rect 23661 18037 23673 18071
rect 23707 18037 23719 18071
rect 23661 18031 23719 18037
rect 26602 18028 26608 18080
rect 26660 18028 26666 18080
rect 27338 18028 27344 18080
rect 27396 18028 27402 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 31588 18077 31616 18244
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 33597 18275 33655 18281
rect 33597 18272 33609 18275
rect 33244 18244 33609 18272
rect 32217 18207 32275 18213
rect 32217 18173 32229 18207
rect 32263 18173 32275 18207
rect 32217 18167 32275 18173
rect 32232 18136 32260 18167
rect 33244 18145 33272 18244
rect 33597 18241 33609 18244
rect 33643 18272 33655 18275
rect 35342 18272 35348 18284
rect 33643 18244 35348 18272
rect 33643 18241 33655 18244
rect 33597 18235 33655 18241
rect 35342 18232 35348 18244
rect 35400 18232 35406 18284
rect 33318 18164 33324 18216
rect 33376 18164 33382 18216
rect 33229 18139 33287 18145
rect 32232 18108 32352 18136
rect 32324 18080 32352 18108
rect 33229 18105 33241 18139
rect 33275 18105 33287 18139
rect 33229 18099 33287 18105
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 30800 18040 31585 18068
rect 30800 18028 30806 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 31573 18031 31631 18037
rect 32306 18028 32312 18080
rect 32364 18068 32370 18080
rect 32674 18068 32680 18080
rect 32364 18040 32680 18068
rect 32364 18028 32370 18040
rect 32674 18028 32680 18040
rect 32732 18028 32738 18080
rect 34330 18028 34336 18080
rect 34388 18028 34394 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 8754 17824 8760 17876
rect 8812 17864 8818 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 8812 17836 9045 17864
rect 8812 17824 8818 17836
rect 9033 17833 9045 17836
rect 9079 17833 9091 17867
rect 9033 17827 9091 17833
rect 9493 17867 9551 17873
rect 9493 17833 9505 17867
rect 9539 17864 9551 17867
rect 9766 17864 9772 17876
rect 9539 17836 9772 17864
rect 9539 17833 9551 17836
rect 9493 17827 9551 17833
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 9858 17824 9864 17876
rect 9916 17824 9922 17876
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 14826 17864 14832 17876
rect 12952 17836 14832 17864
rect 12952 17824 12958 17836
rect 14826 17824 14832 17836
rect 14884 17864 14890 17876
rect 20809 17867 20867 17873
rect 20809 17864 20821 17867
rect 14884 17836 20821 17864
rect 14884 17824 14890 17836
rect 20809 17833 20821 17836
rect 20855 17864 20867 17867
rect 21358 17864 21364 17876
rect 20855 17836 21364 17864
rect 20855 17833 20867 17836
rect 20809 17827 20867 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22278 17824 22284 17876
rect 22336 17864 22342 17876
rect 25222 17864 25228 17876
rect 22336 17836 23704 17864
rect 22336 17824 22342 17836
rect 14274 17756 14280 17808
rect 14332 17796 14338 17808
rect 20073 17799 20131 17805
rect 14332 17768 15056 17796
rect 14332 17756 14338 17768
rect 10870 17688 10876 17740
rect 10928 17688 10934 17740
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17728 11575 17731
rect 11606 17728 11612 17740
rect 11563 17700 11612 17728
rect 11563 17697 11575 17700
rect 11517 17691 11575 17697
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 15028 17737 15056 17768
rect 20073 17765 20085 17799
rect 20119 17796 20131 17799
rect 20254 17796 20260 17808
rect 20119 17768 20260 17796
rect 20119 17765 20131 17768
rect 20073 17759 20131 17765
rect 20254 17756 20260 17768
rect 20312 17756 20318 17808
rect 21634 17756 21640 17808
rect 21692 17796 21698 17808
rect 21818 17796 21824 17808
rect 21692 17768 21824 17796
rect 21692 17756 21698 17768
rect 21818 17756 21824 17768
rect 21876 17796 21882 17808
rect 21876 17768 21956 17796
rect 21876 17756 21882 17768
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 14292 17700 14749 17728
rect 9214 17620 9220 17672
rect 9272 17620 9278 17672
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 9674 17660 9680 17672
rect 9447 17632 9680 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9416 17592 9444 17623
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10284 17632 10609 17660
rect 10284 17620 10290 17632
rect 10597 17629 10609 17632
rect 10643 17660 10655 17663
rect 12345 17663 12403 17669
rect 10643 17632 11454 17660
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12526 17660 12532 17672
rect 12391 17632 12532 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12526 17620 12532 17632
rect 12584 17660 12590 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 12584 17632 12633 17660
rect 12584 17620 12590 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12805 17663 12863 17669
rect 12805 17629 12817 17663
rect 12851 17660 12863 17663
rect 12986 17660 12992 17672
rect 12851 17632 12992 17660
rect 12851 17629 12863 17632
rect 12805 17623 12863 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 14292 17669 14320 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 14737 17691 14795 17697
rect 15013 17731 15071 17737
rect 15013 17697 15025 17731
rect 15059 17697 15071 17731
rect 19978 17728 19984 17740
rect 15013 17691 15071 17697
rect 16132 17700 19984 17728
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14550 17660 14556 17672
rect 14507 17632 14556 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 14645 17663 14703 17669
rect 14645 17629 14657 17663
rect 14691 17660 14703 17663
rect 14826 17660 14832 17672
rect 14691 17632 14832 17660
rect 14691 17629 14703 17632
rect 14645 17623 14703 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 15102 17620 15108 17672
rect 15160 17620 15166 17672
rect 9140 17564 9444 17592
rect 14369 17595 14427 17601
rect 9140 17536 9168 17564
rect 14369 17561 14381 17595
rect 14415 17592 14427 17595
rect 14734 17592 14740 17604
rect 14415 17564 14740 17592
rect 14415 17561 14427 17564
rect 14369 17555 14427 17561
rect 14734 17552 14740 17564
rect 14792 17592 14798 17604
rect 16132 17592 16160 17700
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 21928 17728 21956 17768
rect 22005 17731 22063 17737
rect 22005 17728 22017 17731
rect 21928 17700 22017 17728
rect 22005 17697 22017 17700
rect 22051 17697 22063 17731
rect 23676 17728 23704 17836
rect 24596 17836 25228 17864
rect 23750 17728 23756 17740
rect 23676 17700 23756 17728
rect 22005 17691 22063 17697
rect 23750 17688 23756 17700
rect 23808 17688 23814 17740
rect 24596 17737 24624 17836
rect 25222 17824 25228 17836
rect 25280 17864 25286 17876
rect 25774 17864 25780 17876
rect 25280 17836 25780 17864
rect 25280 17824 25286 17836
rect 25774 17824 25780 17836
rect 25832 17824 25838 17876
rect 27338 17824 27344 17876
rect 27396 17864 27402 17876
rect 28077 17867 28135 17873
rect 28077 17864 28089 17867
rect 27396 17836 28089 17864
rect 27396 17824 27402 17836
rect 28077 17833 28089 17836
rect 28123 17833 28135 17867
rect 28077 17827 28135 17833
rect 29546 17824 29552 17876
rect 29604 17864 29610 17876
rect 30285 17867 30343 17873
rect 30285 17864 30297 17867
rect 29604 17836 30297 17864
rect 29604 17824 29610 17836
rect 30285 17833 30297 17836
rect 30331 17833 30343 17867
rect 30285 17827 30343 17833
rect 32490 17824 32496 17876
rect 32548 17864 32554 17876
rect 32769 17867 32827 17873
rect 32769 17864 32781 17867
rect 32548 17836 32781 17864
rect 32548 17824 32554 17836
rect 32769 17833 32781 17836
rect 32815 17833 32827 17867
rect 32769 17827 32827 17833
rect 32950 17824 32956 17876
rect 33008 17864 33014 17876
rect 33137 17867 33195 17873
rect 33137 17864 33149 17867
rect 33008 17836 33149 17864
rect 33008 17824 33014 17836
rect 33137 17833 33149 17836
rect 33183 17833 33195 17867
rect 33137 17827 33195 17833
rect 33502 17824 33508 17876
rect 33560 17864 33566 17876
rect 34330 17864 34336 17876
rect 33560 17836 34336 17864
rect 33560 17824 33566 17836
rect 34330 17824 34336 17836
rect 34388 17824 34394 17876
rect 25593 17799 25651 17805
rect 25593 17765 25605 17799
rect 25639 17765 25651 17799
rect 34054 17796 34060 17808
rect 25593 17759 25651 17765
rect 27632 17768 34060 17796
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17697 24639 17731
rect 25608 17728 25636 17759
rect 25682 17728 25688 17740
rect 25608 17700 25688 17728
rect 24581 17691 24639 17697
rect 25682 17688 25688 17700
rect 25740 17728 25746 17740
rect 27632 17728 27660 17768
rect 34054 17756 34060 17768
rect 34112 17756 34118 17808
rect 29178 17728 29184 17740
rect 25740 17700 27660 17728
rect 28644 17700 29184 17728
rect 25740 17688 25746 17700
rect 17678 17660 17684 17672
rect 16684 17632 17684 17660
rect 16684 17601 16712 17632
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17629 18659 17663
rect 18601 17623 18659 17629
rect 14792 17564 16160 17592
rect 16669 17595 16727 17601
rect 14792 17552 14798 17564
rect 16669 17561 16681 17595
rect 16715 17561 16727 17595
rect 16669 17555 16727 17561
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 12710 17484 12716 17536
rect 12768 17484 12774 17536
rect 14090 17484 14096 17536
rect 14148 17484 14154 17536
rect 16393 17527 16451 17533
rect 16393 17493 16405 17527
rect 16439 17524 16451 17527
rect 17034 17524 17040 17536
rect 16439 17496 17040 17524
rect 16439 17493 16451 17496
rect 16393 17487 16451 17493
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 18616 17524 18644 17623
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 18840 17632 18889 17660
rect 18840 17620 18846 17632
rect 18877 17629 18889 17632
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 19518 17620 19524 17672
rect 19576 17660 19582 17672
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 19576 17632 20269 17660
rect 19576 17620 19582 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17660 20407 17663
rect 21726 17660 21732 17672
rect 20395 17632 21732 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 22281 17663 22339 17669
rect 22281 17660 22293 17663
rect 22066 17632 22293 17660
rect 22066 17604 22094 17632
rect 22281 17629 22293 17632
rect 22327 17660 22339 17663
rect 23293 17663 23351 17669
rect 22327 17632 22784 17660
rect 22327 17629 22339 17632
rect 22281 17623 22339 17629
rect 20073 17595 20131 17601
rect 20073 17561 20085 17595
rect 20119 17592 20131 17595
rect 20622 17592 20628 17604
rect 20119 17564 20628 17592
rect 20119 17561 20131 17564
rect 20073 17555 20131 17561
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 20898 17552 20904 17604
rect 20956 17592 20962 17604
rect 21085 17595 21143 17601
rect 21085 17592 21097 17595
rect 20956 17564 21097 17592
rect 20956 17552 20962 17564
rect 21085 17561 21097 17564
rect 21131 17561 21143 17595
rect 21085 17555 21143 17561
rect 21542 17552 21548 17604
rect 21600 17552 21606 17604
rect 22002 17552 22008 17604
rect 22060 17564 22094 17604
rect 22060 17552 22066 17564
rect 22756 17536 22784 17632
rect 23293 17629 23305 17663
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23308 17536 23336 17623
rect 24026 17620 24032 17672
rect 24084 17620 24090 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17660 24915 17663
rect 25314 17660 25320 17672
rect 24903 17632 25320 17660
rect 24903 17629 24915 17632
rect 24857 17623 24915 17629
rect 25314 17620 25320 17632
rect 25372 17620 25378 17672
rect 28644 17669 28672 17700
rect 29178 17688 29184 17700
rect 29236 17688 29242 17740
rect 29546 17688 29552 17740
rect 29604 17728 29610 17740
rect 29641 17731 29699 17737
rect 29641 17728 29653 17731
rect 29604 17700 29653 17728
rect 29604 17688 29610 17700
rect 29641 17697 29653 17700
rect 29687 17697 29699 17731
rect 29641 17691 29699 17697
rect 30190 17688 30196 17740
rect 30248 17728 30254 17740
rect 30837 17731 30895 17737
rect 30837 17728 30849 17731
rect 30248 17700 30849 17728
rect 30248 17688 30254 17700
rect 30837 17697 30849 17700
rect 30883 17697 30895 17731
rect 30837 17691 30895 17697
rect 32490 17688 32496 17740
rect 32548 17728 32554 17740
rect 32548 17700 33272 17728
rect 32548 17688 32554 17700
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 28353 17663 28411 17669
rect 28353 17629 28365 17663
rect 28399 17660 28411 17663
rect 28629 17663 28687 17669
rect 28629 17660 28641 17663
rect 28399 17632 28641 17660
rect 28399 17629 28411 17632
rect 28353 17623 28411 17629
rect 28629 17629 28641 17632
rect 28675 17629 28687 17663
rect 28629 17623 28687 17629
rect 21726 17524 21732 17536
rect 18616 17496 21732 17524
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 21821 17527 21879 17533
rect 21821 17493 21833 17527
rect 21867 17524 21879 17527
rect 22186 17524 22192 17536
rect 21867 17496 22192 17524
rect 21867 17493 21879 17496
rect 21821 17487 21879 17493
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 23014 17484 23020 17536
rect 23072 17484 23078 17536
rect 23198 17484 23204 17536
rect 23256 17484 23262 17536
rect 23290 17484 23296 17536
rect 23348 17484 23354 17536
rect 26344 17524 26372 17623
rect 26602 17552 26608 17604
rect 26660 17552 26666 17604
rect 28261 17595 28319 17601
rect 28261 17592 28273 17595
rect 27830 17564 28273 17592
rect 28261 17561 28273 17564
rect 28307 17561 28319 17595
rect 28261 17555 28319 17561
rect 28368 17536 28396 17623
rect 29362 17620 29368 17672
rect 29420 17660 29426 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29420 17632 29745 17660
rect 29420 17620 29426 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 29748 17592 29776 17623
rect 30558 17620 30564 17672
rect 30616 17660 30622 17672
rect 31294 17660 31300 17672
rect 30616 17632 31300 17660
rect 30616 17620 30622 17632
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 33244 17669 33272 17700
rect 32677 17663 32735 17669
rect 32677 17629 32689 17663
rect 32723 17629 32735 17663
rect 32677 17623 32735 17629
rect 33229 17663 33287 17669
rect 33229 17629 33241 17663
rect 33275 17629 33287 17663
rect 33229 17623 33287 17629
rect 32398 17592 32404 17604
rect 29748 17564 32404 17592
rect 32398 17552 32404 17564
rect 32456 17552 32462 17604
rect 32692 17592 32720 17623
rect 33502 17620 33508 17672
rect 33560 17620 33566 17672
rect 32858 17592 32864 17604
rect 32692 17564 32864 17592
rect 32858 17552 32864 17564
rect 32916 17592 32922 17604
rect 33520 17592 33548 17620
rect 32916 17564 33548 17592
rect 32916 17552 32922 17564
rect 27522 17524 27528 17536
rect 26344 17496 27528 17524
rect 27522 17484 27528 17496
rect 27580 17484 27586 17536
rect 28350 17484 28356 17536
rect 28408 17484 28414 17536
rect 28626 17484 28632 17536
rect 28684 17524 28690 17536
rect 28721 17527 28779 17533
rect 28721 17524 28733 17527
rect 28684 17496 28733 17524
rect 28684 17484 28690 17496
rect 28721 17493 28733 17496
rect 28767 17493 28779 17527
rect 28721 17487 28779 17493
rect 30098 17484 30104 17536
rect 30156 17484 30162 17536
rect 30650 17484 30656 17536
rect 30708 17484 30714 17536
rect 30742 17484 30748 17536
rect 30800 17484 30806 17536
rect 32214 17484 32220 17536
rect 32272 17524 32278 17536
rect 33042 17524 33048 17536
rect 32272 17496 33048 17524
rect 32272 17484 32278 17496
rect 33042 17484 33048 17496
rect 33100 17484 33106 17536
rect 33686 17484 33692 17536
rect 33744 17484 33750 17536
rect 1104 17434 38824 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 38824 17434
rect 1104 17360 38824 17382
rect 11606 17280 11612 17332
rect 11664 17280 11670 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 12768 17292 13829 17320
rect 12768 17280 12774 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 14645 17323 14703 17329
rect 14645 17289 14657 17323
rect 14691 17320 14703 17323
rect 15102 17320 15108 17332
rect 14691 17292 15108 17320
rect 14691 17289 14703 17292
rect 14645 17283 14703 17289
rect 10413 17255 10471 17261
rect 10413 17221 10425 17255
rect 10459 17252 10471 17255
rect 11330 17252 11336 17264
rect 10459 17224 11336 17252
rect 10459 17221 10471 17224
rect 10413 17215 10471 17221
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17184 11575 17187
rect 11624 17184 11652 17280
rect 14660 17252 14688 17283
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 18874 17320 18880 17332
rect 17328 17292 18880 17320
rect 14200 17224 14688 17252
rect 14200 17193 14228 17224
rect 11563 17156 11652 17184
rect 14185 17187 14243 17193
rect 11563 17153 11575 17156
rect 11517 17147 11575 17153
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 14274 17144 14280 17196
rect 14332 17144 14338 17196
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17184 14611 17187
rect 14642 17184 14648 17196
rect 14599 17156 14648 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 14737 17187 14795 17193
rect 14737 17153 14749 17187
rect 14783 17184 14795 17187
rect 14918 17184 14924 17196
rect 14783 17156 14924 17184
rect 14783 17153 14795 17156
rect 14737 17147 14795 17153
rect 14918 17144 14924 17156
rect 14976 17144 14982 17196
rect 17328 17193 17356 17292
rect 18874 17280 18880 17292
rect 18932 17320 18938 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 18932 17292 19625 17320
rect 18932 17280 18938 17292
rect 19613 17289 19625 17292
rect 19659 17289 19671 17323
rect 19613 17283 19671 17289
rect 21637 17323 21695 17329
rect 21637 17289 21649 17323
rect 21683 17289 21695 17323
rect 21637 17283 21695 17289
rect 17402 17212 17408 17264
rect 17460 17212 17466 17264
rect 21652 17252 21680 17283
rect 22738 17280 22744 17332
rect 22796 17320 22802 17332
rect 23569 17323 23627 17329
rect 23569 17320 23581 17323
rect 22796 17292 23581 17320
rect 22796 17280 22802 17292
rect 23569 17289 23581 17292
rect 23615 17289 23627 17323
rect 23569 17283 23627 17289
rect 23750 17280 23756 17332
rect 23808 17280 23814 17332
rect 24026 17280 24032 17332
rect 24084 17320 24090 17332
rect 24084 17292 30604 17320
rect 24084 17280 24090 17292
rect 22097 17255 22155 17261
rect 22097 17252 22109 17255
rect 17788 17224 19748 17252
rect 21652 17224 22109 17252
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17420 17184 17448 17212
rect 17788 17193 17816 17224
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17420 17156 17785 17184
rect 17313 17147 17371 17153
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 18414 17144 18420 17196
rect 18472 17184 18478 17196
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 18472 17156 18613 17184
rect 18472 17144 18478 17156
rect 18601 17153 18613 17156
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 18874 17144 18880 17196
rect 18932 17144 18938 17196
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 17405 17119 17463 17125
rect 11020 17088 17080 17116
rect 11020 17076 11026 17088
rect 17052 17060 17080 17088
rect 17405 17085 17417 17119
rect 17451 17116 17463 17119
rect 17862 17116 17868 17128
rect 17451 17088 17868 17116
rect 17451 17085 17463 17088
rect 17405 17079 17463 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 16942 17008 16948 17060
rect 17000 17008 17006 17060
rect 17034 17008 17040 17060
rect 17092 17008 17098 17060
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8941 16983 8999 16989
rect 8941 16980 8953 16983
rect 8352 16952 8953 16980
rect 8352 16940 8358 16952
rect 8941 16949 8953 16952
rect 8987 16949 8999 16983
rect 8941 16943 8999 16949
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11974 16980 11980 16992
rect 11655 16952 11980 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 14458 16940 14464 16992
rect 14516 16940 14522 16992
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 18966 16980 18972 16992
rect 17828 16952 18972 16980
rect 17828 16940 17834 16952
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19720 16980 19748 17224
rect 22097 17221 22109 17224
rect 22143 17221 22155 17255
rect 22097 17215 22155 17221
rect 21450 17144 21456 17196
rect 21508 17144 21514 17196
rect 23198 17144 23204 17196
rect 23256 17144 23262 17196
rect 23768 17184 23796 17280
rect 28626 17212 28632 17264
rect 28684 17212 28690 17264
rect 30576 17252 30604 17292
rect 30650 17280 30656 17332
rect 30708 17320 30714 17332
rect 30837 17323 30895 17329
rect 30837 17320 30849 17323
rect 30708 17292 30849 17320
rect 30708 17280 30714 17292
rect 30837 17289 30849 17292
rect 30883 17289 30895 17323
rect 32214 17320 32220 17332
rect 30837 17283 30895 17289
rect 30944 17292 32220 17320
rect 30944 17252 30972 17292
rect 32214 17280 32220 17292
rect 32272 17280 32278 17332
rect 32877 17323 32935 17329
rect 32877 17320 32889 17323
rect 32324 17292 32889 17320
rect 32324 17252 32352 17292
rect 32877 17289 32889 17292
rect 32923 17289 32935 17323
rect 32877 17283 32935 17289
rect 33042 17280 33048 17332
rect 33100 17320 33106 17332
rect 38289 17323 38347 17329
rect 38289 17320 38301 17323
rect 33100 17292 38301 17320
rect 33100 17280 33106 17292
rect 38289 17289 38301 17292
rect 38335 17289 38347 17323
rect 38289 17283 38347 17289
rect 29564 17224 30512 17252
rect 30576 17224 30972 17252
rect 31036 17224 32352 17252
rect 29564 17196 29592 17224
rect 24305 17187 24363 17193
rect 24305 17184 24317 17187
rect 23768 17156 24317 17184
rect 24305 17153 24317 17156
rect 24351 17184 24363 17187
rect 24397 17187 24455 17193
rect 24397 17184 24409 17187
rect 24351 17156 24409 17184
rect 24351 17153 24363 17156
rect 24305 17147 24363 17153
rect 24397 17153 24409 17156
rect 24443 17153 24455 17187
rect 25682 17184 25688 17196
rect 25645 17156 25688 17184
rect 24397 17147 24455 17153
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 25774 17144 25780 17196
rect 25832 17184 25838 17196
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25832 17156 25973 17184
rect 25832 17144 25838 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 29546 17144 29552 17196
rect 29604 17144 29610 17196
rect 29822 17144 29828 17196
rect 29880 17144 29886 17196
rect 30484 17184 30512 17224
rect 31036 17184 31064 17224
rect 32324 17193 32352 17224
rect 32398 17212 32404 17264
rect 32456 17212 32462 17264
rect 32582 17212 32588 17264
rect 32640 17212 32646 17264
rect 32677 17255 32735 17261
rect 32677 17221 32689 17255
rect 32723 17221 32735 17255
rect 32677 17215 32735 17221
rect 30484 17156 31064 17184
rect 31113 17188 31171 17193
rect 31113 17187 31248 17188
rect 31113 17153 31125 17187
rect 31159 17184 31248 17187
rect 32309 17187 32367 17193
rect 31159 17160 31708 17184
rect 31159 17153 31171 17160
rect 31220 17156 31708 17160
rect 31113 17147 31171 17153
rect 31680 17128 31708 17156
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32416 17184 32444 17212
rect 32692 17184 32720 17215
rect 32766 17212 32772 17264
rect 32824 17252 32830 17264
rect 33137 17255 33195 17261
rect 33137 17252 33149 17255
rect 32824 17224 33149 17252
rect 32824 17212 32830 17224
rect 33137 17221 33149 17224
rect 33183 17221 33195 17255
rect 33137 17215 33195 17221
rect 33226 17184 33232 17196
rect 32416 17156 33232 17184
rect 32309 17147 32367 17153
rect 33226 17144 33232 17156
rect 33284 17144 33290 17196
rect 33413 17187 33471 17193
rect 33413 17153 33425 17187
rect 33459 17153 33471 17187
rect 33413 17147 33471 17153
rect 38473 17187 38531 17193
rect 38473 17153 38485 17187
rect 38519 17184 38531 17187
rect 38519 17156 38884 17184
rect 38519 17153 38531 17156
rect 38473 17147 38531 17153
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21818 17116 21824 17128
rect 20772 17088 21824 17116
rect 20772 17076 20778 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 23290 17116 23296 17128
rect 23216 17088 23296 17116
rect 23216 16992 23244 17088
rect 23290 17076 23296 17088
rect 23348 17116 23354 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23348 17088 24041 17116
rect 23348 17076 23354 17088
rect 24029 17085 24041 17088
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 24673 17119 24731 17125
rect 24673 17085 24685 17119
rect 24719 17116 24731 17119
rect 24719 17088 25360 17116
rect 24719 17085 24731 17088
rect 24673 17079 24731 17085
rect 24854 17008 24860 17060
rect 24912 17048 24918 17060
rect 24949 17051 25007 17057
rect 24949 17048 24961 17051
rect 24912 17020 24961 17048
rect 24912 17008 24918 17020
rect 24949 17017 24961 17020
rect 24995 17017 25007 17051
rect 24949 17011 25007 17017
rect 23198 16980 23204 16992
rect 19720 16952 23204 16980
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 25332 16980 25360 17088
rect 27522 17076 27528 17128
rect 27580 17116 27586 17128
rect 27617 17119 27675 17125
rect 27617 17116 27629 17119
rect 27580 17088 27629 17116
rect 27580 17076 27586 17088
rect 27617 17085 27629 17088
rect 27663 17085 27675 17119
rect 27617 17079 27675 17085
rect 27890 17076 27896 17128
rect 27948 17076 27954 17128
rect 29365 17119 29423 17125
rect 29365 17085 29377 17119
rect 29411 17116 29423 17119
rect 29914 17116 29920 17128
rect 29411 17088 29920 17116
rect 29411 17085 29423 17088
rect 29365 17079 29423 17085
rect 29914 17076 29920 17088
rect 29972 17076 29978 17128
rect 30101 17119 30159 17125
rect 30101 17085 30113 17119
rect 30147 17116 30159 17119
rect 30190 17116 30196 17128
rect 30147 17088 30196 17116
rect 30147 17085 30159 17088
rect 30101 17079 30159 17085
rect 30190 17076 30196 17088
rect 30248 17076 30254 17128
rect 30837 17119 30895 17125
rect 30837 17085 30849 17119
rect 30883 17085 30895 17119
rect 30837 17079 30895 17085
rect 29270 17008 29276 17060
rect 29328 17048 29334 17060
rect 29457 17051 29515 17057
rect 29457 17048 29469 17051
rect 29328 17020 29469 17048
rect 29328 17008 29334 17020
rect 29457 17017 29469 17020
rect 29503 17017 29515 17051
rect 30852 17048 30880 17079
rect 31662 17076 31668 17128
rect 31720 17076 31726 17128
rect 33137 17119 33195 17125
rect 33137 17116 33149 17119
rect 32508 17108 32812 17116
rect 32968 17108 33149 17116
rect 32508 17088 33149 17108
rect 32398 17048 32404 17060
rect 30852 17020 32404 17048
rect 29457 17011 29515 17017
rect 32398 17008 32404 17020
rect 32456 17008 32462 17060
rect 28350 16980 28356 16992
rect 25332 16952 28356 16980
rect 28350 16940 28356 16952
rect 28408 16940 28414 16992
rect 31018 16940 31024 16992
rect 31076 16940 31082 16992
rect 31294 16940 31300 16992
rect 31352 16980 31358 16992
rect 32508 16980 32536 17088
rect 32784 17080 32996 17088
rect 33137 17085 33149 17088
rect 33183 17085 33195 17119
rect 33137 17079 33195 17085
rect 32585 17051 32643 17057
rect 32585 17017 32597 17051
rect 32631 17048 32643 17051
rect 33321 17051 33379 17057
rect 33321 17048 33333 17051
rect 32631 17020 33333 17048
rect 32631 17017 32643 17020
rect 32585 17011 32643 17017
rect 33321 17017 33333 17020
rect 33367 17017 33379 17051
rect 33321 17011 33379 17017
rect 31352 16952 32536 16980
rect 31352 16940 31358 16952
rect 32858 16940 32864 16992
rect 32916 16940 32922 16992
rect 33042 16940 33048 16992
rect 33100 16980 33106 16992
rect 33428 16980 33456 17147
rect 38856 17128 38884 17156
rect 38838 17076 38844 17128
rect 38896 17076 38902 17128
rect 33100 16952 33456 16980
rect 33100 16940 33106 16952
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 9585 16779 9643 16785
rect 9585 16776 9597 16779
rect 9272 16748 9597 16776
rect 9272 16736 9278 16748
rect 9585 16745 9597 16748
rect 9631 16745 9643 16779
rect 9585 16739 9643 16745
rect 10226 16736 10232 16788
rect 10284 16776 10290 16788
rect 11885 16779 11943 16785
rect 11885 16776 11897 16779
rect 10284 16748 11897 16776
rect 10284 16736 10290 16748
rect 11885 16745 11897 16748
rect 11931 16776 11943 16779
rect 12437 16779 12495 16785
rect 12437 16776 12449 16779
rect 11931 16748 12449 16776
rect 11931 16745 11943 16748
rect 11885 16739 11943 16745
rect 12437 16745 12449 16748
rect 12483 16745 12495 16779
rect 12437 16739 12495 16745
rect 12710 16736 12716 16788
rect 12768 16736 12774 16788
rect 13541 16779 13599 16785
rect 13541 16745 13553 16779
rect 13587 16776 13599 16779
rect 13814 16776 13820 16788
rect 13587 16748 13820 16776
rect 13587 16745 13599 16748
rect 13541 16739 13599 16745
rect 13814 16736 13820 16748
rect 13872 16736 13878 16788
rect 14274 16736 14280 16788
rect 14332 16736 14338 16788
rect 14458 16736 14464 16788
rect 14516 16736 14522 16788
rect 20714 16776 20720 16788
rect 15764 16748 20720 16776
rect 10244 16708 10272 16736
rect 10060 16680 10272 16708
rect 10060 16649 10088 16680
rect 9217 16643 9275 16649
rect 9217 16609 9229 16643
rect 9263 16640 9275 16643
rect 10045 16643 10103 16649
rect 9263 16612 9996 16640
rect 9263 16609 9275 16612
rect 9217 16603 9275 16609
rect 9968 16584 9996 16612
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16640 10287 16643
rect 10318 16640 10324 16652
rect 10275 16612 10324 16640
rect 10275 16609 10287 16612
rect 10229 16603 10287 16609
rect 10318 16600 10324 16612
rect 10376 16640 10382 16652
rect 10962 16640 10968 16652
rect 10376 16612 10968 16640
rect 10376 16600 10382 16612
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 11204 16612 11345 16640
rect 11204 16600 11210 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 11839 16612 12633 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 9950 16532 9956 16584
rect 10008 16532 10014 16584
rect 10686 16532 10692 16584
rect 10744 16572 10750 16584
rect 11900 16581 11928 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12728 16640 12756 16736
rect 13633 16711 13691 16717
rect 13633 16677 13645 16711
rect 13679 16708 13691 16711
rect 13722 16708 13728 16720
rect 13679 16680 13728 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 13722 16668 13728 16680
rect 13780 16668 13786 16720
rect 13357 16643 13415 16649
rect 13357 16640 13369 16643
rect 12728 16612 13369 16640
rect 12621 16603 12679 16609
rect 13357 16609 13369 16612
rect 13403 16609 13415 16643
rect 14292 16640 14320 16736
rect 13357 16603 13415 16609
rect 13924 16612 14320 16640
rect 14369 16643 14427 16649
rect 10873 16575 10931 16581
rect 10873 16572 10885 16575
rect 10744 16544 10885 16572
rect 10744 16532 10750 16544
rect 10873 16541 10885 16544
rect 10919 16572 10931 16575
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10919 16544 11437 16572
rect 10919 16541 10931 16544
rect 10873 16535 10931 16541
rect 11425 16541 11437 16544
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16541 11943 16575
rect 11885 16535 11943 16541
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12032 16544 12357 16572
rect 12032 16532 12038 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 13265 16575 13323 16581
rect 13265 16572 13277 16575
rect 12345 16535 12403 16541
rect 12636 16544 13277 16572
rect 9398 16464 9404 16516
rect 9456 16464 9462 16516
rect 12158 16504 12164 16516
rect 9968 16476 12164 16504
rect 9968 16445 9996 16476
rect 12158 16464 12164 16476
rect 12216 16464 12222 16516
rect 12636 16513 12664 16544
rect 13265 16541 13277 16544
rect 13311 16572 13323 16575
rect 13538 16572 13544 16584
rect 13311 16544 13544 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13538 16532 13544 16544
rect 13596 16572 13602 16584
rect 13924 16581 13952 16612
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 14476 16640 14504 16736
rect 15764 16649 15792 16748
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 21450 16736 21456 16788
rect 21508 16776 21514 16788
rect 21637 16779 21695 16785
rect 21637 16776 21649 16779
rect 21508 16748 21649 16776
rect 21508 16736 21514 16748
rect 21637 16745 21649 16748
rect 21683 16745 21695 16779
rect 21637 16739 21695 16745
rect 21726 16736 21732 16788
rect 21784 16776 21790 16788
rect 21784 16748 23704 16776
rect 21784 16736 21790 16748
rect 18785 16711 18843 16717
rect 18785 16677 18797 16711
rect 18831 16708 18843 16711
rect 18874 16708 18880 16720
rect 18831 16680 18880 16708
rect 18831 16677 18843 16680
rect 18785 16671 18843 16677
rect 18874 16668 18880 16680
rect 18932 16708 18938 16720
rect 18932 16680 19288 16708
rect 18932 16668 18938 16680
rect 19260 16652 19288 16680
rect 14415 16612 14504 16640
rect 15749 16643 15807 16649
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 15749 16609 15761 16643
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 17770 16600 17776 16652
rect 17828 16600 17834 16652
rect 19242 16600 19248 16652
rect 19300 16600 19306 16652
rect 20165 16643 20223 16649
rect 19536 16612 19840 16640
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 13596 16544 13645 16572
rect 13596 16532 13602 16544
rect 13633 16541 13645 16544
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 13909 16575 13967 16581
rect 13909 16541 13921 16575
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 17678 16572 17684 16584
rect 17158 16544 17684 16572
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17880 16544 18061 16572
rect 12621 16507 12679 16513
rect 12621 16473 12633 16507
rect 12667 16473 12679 16507
rect 13354 16504 13360 16516
rect 12621 16467 12679 16473
rect 12912 16476 13360 16504
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16405 10011 16439
rect 9953 16399 10011 16405
rect 10410 16396 10416 16448
rect 10468 16396 10474 16448
rect 10778 16396 10784 16448
rect 10836 16396 10842 16448
rect 12912 16445 12940 16476
rect 13354 16464 13360 16476
rect 13412 16504 13418 16516
rect 13725 16507 13783 16513
rect 13725 16504 13737 16507
rect 13412 16476 13737 16504
rect 13412 16464 13418 16476
rect 13725 16473 13737 16476
rect 13771 16473 13783 16507
rect 13725 16467 13783 16473
rect 16022 16464 16028 16516
rect 16080 16464 16086 16516
rect 17880 16448 17908 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 18049 16535 18107 16541
rect 18984 16544 19441 16572
rect 18984 16448 19012 16544
rect 19429 16541 19441 16544
rect 19475 16572 19487 16575
rect 19536 16572 19564 16612
rect 19475 16544 19564 16572
rect 19613 16575 19671 16581
rect 19475 16541 19487 16544
rect 19429 16535 19487 16541
rect 19613 16541 19625 16575
rect 19659 16572 19671 16575
rect 19659 16544 19748 16572
rect 19659 16541 19671 16544
rect 19613 16535 19671 16541
rect 12253 16439 12311 16445
rect 12253 16405 12265 16439
rect 12299 16436 12311 16439
rect 12897 16439 12955 16445
rect 12897 16436 12909 16439
rect 12299 16408 12909 16436
rect 12299 16405 12311 16408
rect 12253 16399 12311 16405
rect 12897 16405 12909 16408
rect 12943 16405 12955 16439
rect 12897 16399 12955 16405
rect 14642 16396 14648 16448
rect 14700 16396 14706 16448
rect 17497 16439 17555 16445
rect 17497 16405 17509 16439
rect 17543 16436 17555 16439
rect 17862 16436 17868 16448
rect 17543 16408 17868 16436
rect 17543 16405 17555 16408
rect 17497 16399 17555 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 18966 16396 18972 16448
rect 19024 16396 19030 16448
rect 19610 16396 19616 16448
rect 19668 16396 19674 16448
rect 19720 16445 19748 16544
rect 19812 16504 19840 16612
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 22002 16640 22008 16652
rect 20211 16612 22008 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 22002 16600 22008 16612
rect 22060 16640 22066 16652
rect 22097 16643 22155 16649
rect 22097 16640 22109 16643
rect 22060 16612 22109 16640
rect 22060 16600 22066 16612
rect 22097 16609 22109 16612
rect 22143 16609 22155 16643
rect 22097 16603 22155 16609
rect 22186 16600 22192 16652
rect 22244 16600 22250 16652
rect 23676 16649 23704 16748
rect 27890 16736 27896 16788
rect 27948 16776 27954 16788
rect 28169 16779 28227 16785
rect 28169 16776 28181 16779
rect 27948 16748 28181 16776
rect 27948 16736 27954 16748
rect 28169 16745 28181 16748
rect 28215 16745 28227 16779
rect 28169 16739 28227 16745
rect 29641 16779 29699 16785
rect 29641 16745 29653 16779
rect 29687 16776 29699 16779
rect 29822 16776 29828 16788
rect 29687 16748 29828 16776
rect 29687 16745 29699 16748
rect 29641 16739 29699 16745
rect 29822 16736 29828 16748
rect 29880 16736 29886 16788
rect 30745 16779 30803 16785
rect 30745 16745 30757 16779
rect 30791 16776 30803 16779
rect 31018 16776 31024 16788
rect 30791 16748 31024 16776
rect 30791 16745 30803 16748
rect 30745 16739 30803 16745
rect 31018 16736 31024 16748
rect 31076 16736 31082 16788
rect 31128 16748 31616 16776
rect 31128 16708 31156 16748
rect 30944 16680 31156 16708
rect 31588 16708 31616 16748
rect 31662 16736 31668 16788
rect 31720 16736 31726 16788
rect 32950 16736 32956 16788
rect 33008 16776 33014 16788
rect 33689 16779 33747 16785
rect 33689 16776 33701 16779
rect 33008 16748 33701 16776
rect 33008 16736 33014 16748
rect 33689 16745 33701 16748
rect 33735 16745 33747 16779
rect 33689 16739 33747 16745
rect 31588 16680 31708 16708
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 29270 16600 29276 16652
rect 29328 16600 29334 16652
rect 30944 16640 30972 16680
rect 29932 16612 30972 16640
rect 19886 16532 19892 16584
rect 19944 16572 19950 16584
rect 20073 16575 20131 16581
rect 20073 16572 20085 16575
rect 19944 16544 20085 16572
rect 19944 16532 19950 16544
rect 20073 16541 20085 16544
rect 20119 16541 20131 16575
rect 20073 16535 20131 16541
rect 20349 16507 20407 16513
rect 20349 16504 20361 16507
rect 19812 16476 20361 16504
rect 20349 16473 20361 16476
rect 20395 16473 20407 16507
rect 20349 16467 20407 16473
rect 20533 16507 20591 16513
rect 20533 16473 20545 16507
rect 20579 16473 20591 16507
rect 22204 16504 22232 16600
rect 22554 16532 22560 16584
rect 22612 16532 22618 16584
rect 23014 16532 23020 16584
rect 23072 16572 23078 16584
rect 23385 16575 23443 16581
rect 23385 16572 23397 16575
rect 23072 16544 23397 16572
rect 23072 16532 23078 16544
rect 23385 16541 23397 16544
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23290 16504 23296 16516
rect 22204 16476 23296 16504
rect 20533 16467 20591 16473
rect 19705 16439 19763 16445
rect 19705 16405 19717 16439
rect 19751 16436 19763 16439
rect 20548 16436 20576 16467
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 23400 16504 23428 16535
rect 24670 16532 24676 16584
rect 24728 16532 24734 16584
rect 28353 16575 28411 16581
rect 24780 16544 26188 16572
rect 24780 16504 24808 16544
rect 23400 16476 24808 16504
rect 26050 16464 26056 16516
rect 26108 16464 26114 16516
rect 26160 16504 26188 16544
rect 28353 16541 28365 16575
rect 28399 16572 28411 16575
rect 29288 16572 29316 16600
rect 29932 16581 29960 16612
rect 28399 16544 29316 16572
rect 29825 16575 29883 16581
rect 28399 16541 28411 16544
rect 28353 16535 28411 16541
rect 29825 16541 29837 16575
rect 29871 16541 29883 16575
rect 29825 16535 29883 16541
rect 29917 16575 29975 16581
rect 29917 16541 29929 16575
rect 29963 16541 29975 16575
rect 29917 16535 29975 16541
rect 29270 16504 29276 16516
rect 26160 16476 29276 16504
rect 29270 16464 29276 16476
rect 29328 16464 29334 16516
rect 19751 16408 20576 16436
rect 19751 16405 19763 16408
rect 19705 16399 19763 16405
rect 20714 16396 20720 16448
rect 20772 16396 20778 16448
rect 22005 16439 22063 16445
rect 22005 16405 22017 16439
rect 22051 16436 22063 16439
rect 22462 16436 22468 16448
rect 22051 16408 22468 16436
rect 22051 16405 22063 16408
rect 22005 16399 22063 16405
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 24489 16439 24547 16445
rect 24489 16405 24501 16439
rect 24535 16436 24547 16439
rect 25406 16436 25412 16448
rect 24535 16408 25412 16436
rect 24535 16405 24547 16408
rect 24489 16399 24547 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 26142 16396 26148 16448
rect 26200 16436 26206 16448
rect 27062 16436 27068 16448
rect 26200 16408 27068 16436
rect 26200 16396 26206 16408
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 29840 16436 29868 16535
rect 30098 16532 30104 16584
rect 30156 16581 30162 16584
rect 30156 16575 30185 16581
rect 30173 16541 30185 16575
rect 30156 16535 30185 16541
rect 30285 16575 30343 16581
rect 30285 16541 30297 16575
rect 30331 16572 30343 16575
rect 30558 16572 30564 16584
rect 30331 16544 30564 16572
rect 30331 16541 30343 16544
rect 30285 16535 30343 16541
rect 30156 16532 30162 16535
rect 30558 16532 30564 16544
rect 30616 16532 30622 16584
rect 30944 16581 30972 16612
rect 31018 16600 31024 16652
rect 31076 16640 31082 16652
rect 31570 16640 31576 16652
rect 31076 16612 31121 16640
rect 31076 16600 31082 16612
rect 31205 16609 31263 16615
rect 30929 16575 30987 16581
rect 30929 16541 30941 16575
rect 30975 16541 30987 16575
rect 30929 16535 30987 16541
rect 31113 16575 31171 16581
rect 31113 16541 31125 16575
rect 31159 16541 31171 16575
rect 31205 16575 31217 16609
rect 31251 16606 31263 16609
rect 31312 16612 31576 16640
rect 31312 16606 31340 16612
rect 31251 16578 31340 16606
rect 31570 16600 31576 16612
rect 31628 16600 31634 16652
rect 31251 16575 31263 16578
rect 31205 16569 31263 16575
rect 31389 16575 31447 16581
rect 31113 16535 31171 16541
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31680 16572 31708 16680
rect 32968 16640 32996 16736
rect 33226 16668 33232 16720
rect 33284 16668 33290 16720
rect 32784 16612 32996 16640
rect 32784 16581 32812 16612
rect 31435 16544 31708 16572
rect 32585 16575 32643 16581
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 32585 16541 32597 16575
rect 32631 16541 32643 16575
rect 32585 16535 32643 16541
rect 32769 16575 32827 16581
rect 32769 16541 32781 16575
rect 32815 16541 32827 16575
rect 32769 16535 32827 16541
rect 32861 16575 32919 16581
rect 32861 16541 32873 16575
rect 32907 16572 32919 16575
rect 33686 16572 33692 16584
rect 32907 16544 33692 16572
rect 32907 16541 32919 16544
rect 32861 16535 32919 16541
rect 30006 16464 30012 16516
rect 30064 16464 30070 16516
rect 30466 16464 30472 16516
rect 30524 16504 30530 16516
rect 30944 16504 30972 16535
rect 30524 16476 30972 16504
rect 31128 16504 31156 16535
rect 31665 16507 31723 16513
rect 31665 16504 31677 16507
rect 31128 16476 31677 16504
rect 30524 16464 30530 16476
rect 31665 16473 31677 16476
rect 31711 16504 31723 16507
rect 32122 16504 32128 16516
rect 31711 16476 32128 16504
rect 31711 16473 31723 16476
rect 31665 16467 31723 16473
rect 32122 16464 32128 16476
rect 32180 16464 32186 16516
rect 32600 16504 32628 16535
rect 33686 16532 33692 16544
rect 33744 16532 33750 16584
rect 32600 16476 32904 16504
rect 31018 16436 31024 16448
rect 29840 16408 31024 16436
rect 31018 16396 31024 16408
rect 31076 16396 31082 16448
rect 31110 16396 31116 16448
rect 31168 16436 31174 16448
rect 31386 16436 31392 16448
rect 31168 16408 31392 16436
rect 31168 16396 31174 16408
rect 31386 16396 31392 16408
rect 31444 16436 31450 16448
rect 31481 16439 31539 16445
rect 31481 16436 31493 16439
rect 31444 16408 31493 16436
rect 31444 16396 31450 16408
rect 31481 16405 31493 16408
rect 31527 16405 31539 16439
rect 31481 16399 31539 16405
rect 32398 16396 32404 16448
rect 32456 16396 32462 16448
rect 32876 16436 32904 16476
rect 32950 16464 32956 16516
rect 33008 16464 33014 16516
rect 33873 16507 33931 16513
rect 33873 16504 33885 16507
rect 33428 16476 33885 16504
rect 33428 16445 33456 16476
rect 33873 16473 33885 16476
rect 33919 16473 33931 16507
rect 33873 16467 33931 16473
rect 33413 16439 33471 16445
rect 33413 16436 33425 16439
rect 32876 16408 33425 16436
rect 33413 16405 33425 16408
rect 33459 16405 33471 16439
rect 33413 16399 33471 16405
rect 33502 16396 33508 16448
rect 33560 16396 33566 16448
rect 33686 16445 33692 16448
rect 33673 16439 33692 16445
rect 33673 16405 33685 16439
rect 33673 16399 33692 16405
rect 33686 16396 33692 16399
rect 33744 16396 33750 16448
rect 1104 16346 38824 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 38824 16346
rect 1104 16272 38824 16294
rect 10778 16192 10784 16244
rect 10836 16232 10842 16244
rect 13541 16235 13599 16241
rect 10836 16204 13400 16232
rect 10836 16192 10842 16204
rect 8294 16164 8300 16176
rect 7760 16136 8300 16164
rect 7760 16040 7788 16136
rect 8294 16124 8300 16136
rect 8352 16124 8358 16176
rect 9677 16167 9735 16173
rect 9677 16164 9689 16167
rect 9246 16136 9689 16164
rect 9677 16133 9689 16136
rect 9723 16133 9735 16167
rect 9677 16127 9735 16133
rect 11057 16167 11115 16173
rect 11057 16133 11069 16167
rect 11103 16164 11115 16167
rect 11146 16164 11152 16176
rect 11103 16136 11152 16164
rect 11103 16133 11115 16136
rect 11057 16127 11115 16133
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 7742 15988 7748 16040
rect 7800 15988 7806 16040
rect 8018 15988 8024 16040
rect 8076 15988 8082 16040
rect 9784 16028 9812 16059
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 10100 16068 10149 16096
rect 10100 16056 10106 16068
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10137 16059 10195 16065
rect 9140 16000 9812 16028
rect 9861 16031 9919 16037
rect 9140 15972 9168 16000
rect 9861 15997 9873 16031
rect 9907 15997 9919 16031
rect 11072 16028 11100 16127
rect 11146 16124 11152 16136
rect 11204 16164 11210 16176
rect 11204 16136 11836 16164
rect 11204 16124 11210 16136
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16096 11391 16099
rect 11514 16096 11520 16108
rect 11379 16068 11520 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 9861 15991 9919 15997
rect 10888 16000 11100 16028
rect 11256 16028 11284 16059
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 11606 16056 11612 16108
rect 11664 16056 11670 16108
rect 11808 16105 11836 16136
rect 12066 16124 12072 16176
rect 12124 16164 12130 16176
rect 12437 16167 12495 16173
rect 12437 16164 12449 16167
rect 12124 16136 12449 16164
rect 12124 16124 12130 16136
rect 12437 16133 12449 16136
rect 12483 16133 12495 16167
rect 13372 16164 13400 16204
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 14274 16232 14280 16244
rect 13587 16204 14280 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 14274 16192 14280 16204
rect 14332 16192 14338 16244
rect 14369 16235 14427 16241
rect 14369 16201 14381 16235
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 14384 16164 14412 16195
rect 14642 16192 14648 16244
rect 14700 16192 14706 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 16080 16204 16313 16232
rect 16080 16192 16086 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 16301 16195 16359 16201
rect 18966 16192 18972 16244
rect 19024 16192 19030 16244
rect 19610 16192 19616 16244
rect 19668 16192 19674 16244
rect 25424 16204 26740 16232
rect 14660 16164 14688 16192
rect 13372 16136 14412 16164
rect 14568 16136 14688 16164
rect 17313 16167 17371 16173
rect 12437 16127 12495 16133
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 11624 16028 11652 16056
rect 11256 16000 11652 16028
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 9876 15960 9904 15991
rect 10888 15969 10916 16000
rect 10873 15963 10931 15969
rect 9876 15932 9996 15960
rect 9968 15904 9996 15932
rect 10873 15929 10885 15963
rect 10919 15929 10931 15963
rect 10873 15923 10931 15929
rect 11057 15963 11115 15969
rect 11057 15929 11069 15963
rect 11103 15960 11115 15963
rect 12268 15960 12296 16059
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 14568 16105 14596 16136
rect 17313 16133 17325 16167
rect 17359 16164 17371 16167
rect 17862 16164 17868 16176
rect 17359 16136 17868 16164
rect 17359 16133 17371 16136
rect 17313 16127 17371 16133
rect 17862 16124 17868 16136
rect 17920 16164 17926 16176
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 17920 16136 18521 16164
rect 17920 16124 17926 16136
rect 18509 16133 18521 16136
rect 18555 16133 18567 16167
rect 18509 16127 18567 16133
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 14642 16056 14648 16108
rect 14700 16056 14706 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15102 16096 15108 16108
rect 14967 16068 15108 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 12621 16031 12679 16037
rect 12621 15997 12633 16031
rect 12667 16028 12679 16031
rect 14752 16028 14780 16059
rect 15102 16056 15108 16068
rect 15160 16096 15166 16108
rect 16114 16096 16120 16108
rect 15160 16068 16120 16096
rect 15160 16056 15166 16068
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 17221 16099 17279 16105
rect 16531 16068 16896 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 12667 16000 14780 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 16868 15969 16896 16068
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 18414 16096 18420 16108
rect 17267 16068 18420 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 19628 16096 19656 16192
rect 25424 16176 25452 16204
rect 20714 16124 20720 16176
rect 20772 16124 20778 16176
rect 20901 16167 20959 16173
rect 20901 16133 20913 16167
rect 20947 16164 20959 16167
rect 22002 16164 22008 16176
rect 20947 16136 22008 16164
rect 20947 16133 20959 16136
rect 20901 16127 20959 16133
rect 22002 16124 22008 16136
rect 22060 16124 22066 16176
rect 23658 16124 23664 16176
rect 23716 16124 23722 16176
rect 25406 16124 25412 16176
rect 25464 16124 25470 16176
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19628 16068 19993 16096
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16096 20223 16099
rect 20732 16096 20760 16124
rect 20211 16068 20760 16096
rect 20211 16065 20223 16068
rect 20165 16059 20223 16065
rect 23750 16056 23756 16108
rect 23808 16096 23814 16108
rect 24121 16099 24179 16105
rect 24121 16096 24133 16099
rect 23808 16068 24133 16096
rect 23808 16056 23814 16068
rect 24121 16065 24133 16068
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 26418 16056 26424 16108
rect 26476 16056 26482 16108
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 17092 16000 17417 16028
rect 17092 15988 17098 16000
rect 17405 15997 17417 16000
rect 17451 15997 17463 16031
rect 17405 15991 17463 15997
rect 23845 16031 23903 16037
rect 23845 15997 23857 16031
rect 23891 15997 23903 16031
rect 23845 15991 23903 15997
rect 25041 16031 25099 16037
rect 25041 15997 25053 16031
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 25317 16031 25375 16037
rect 25317 15997 25329 16031
rect 25363 16028 25375 16031
rect 25866 16028 25872 16040
rect 25363 16000 25872 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 11103 15932 12296 15960
rect 16853 15963 16911 15969
rect 11103 15929 11115 15932
rect 11057 15923 11115 15929
rect 16853 15929 16865 15963
rect 16899 15929 16911 15963
rect 16853 15923 16911 15929
rect 18782 15920 18788 15972
rect 18840 15960 18846 15972
rect 19794 15960 19800 15972
rect 18840 15932 19800 15960
rect 18840 15920 18846 15932
rect 19794 15920 19800 15932
rect 19852 15920 19858 15972
rect 19886 15920 19892 15972
rect 19944 15960 19950 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 19944 15932 21189 15960
rect 19944 15920 19950 15932
rect 21177 15929 21189 15932
rect 21223 15960 21235 15963
rect 22554 15960 22560 15972
rect 21223 15932 22560 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 22554 15920 22560 15932
rect 22612 15920 22618 15972
rect 23860 15960 23888 15991
rect 23860 15932 23980 15960
rect 23952 15904 23980 15932
rect 9493 15895 9551 15901
rect 9493 15861 9505 15895
rect 9539 15892 9551 15895
rect 9858 15892 9864 15904
rect 9539 15864 9864 15892
rect 9539 15861 9551 15864
rect 9493 15855 9551 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 9950 15852 9956 15904
rect 10008 15852 10014 15904
rect 11974 15852 11980 15904
rect 12032 15852 12038 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 14090 15892 14096 15904
rect 12216 15864 14096 15892
rect 12216 15852 12222 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 20070 15852 20076 15904
rect 20128 15852 20134 15904
rect 21361 15895 21419 15901
rect 21361 15861 21373 15895
rect 21407 15892 21419 15895
rect 21542 15892 21548 15904
rect 21407 15864 21548 15892
rect 21407 15861 21419 15864
rect 21361 15855 21419 15861
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 23569 15895 23627 15901
rect 23569 15861 23581 15895
rect 23615 15892 23627 15895
rect 23934 15892 23940 15904
rect 23615 15864 23940 15892
rect 23615 15861 23627 15864
rect 23569 15855 23627 15861
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 24854 15852 24860 15904
rect 24912 15852 24918 15904
rect 25056 15892 25084 15991
rect 25866 15988 25872 16000
rect 25924 15988 25930 16040
rect 26712 15960 26740 16204
rect 29914 16192 29920 16244
rect 29972 16192 29978 16244
rect 32122 16232 32128 16244
rect 30760 16204 32128 16232
rect 29932 16164 29960 16192
rect 30760 16173 30788 16204
rect 32122 16192 32128 16204
rect 32180 16192 32186 16244
rect 32950 16232 32956 16244
rect 32892 16204 32956 16232
rect 29012 16136 29960 16164
rect 30745 16167 30803 16173
rect 27246 16096 27252 16108
rect 26804 16068 27252 16096
rect 26804 16037 26832 16068
rect 27246 16056 27252 16068
rect 27304 16056 27310 16108
rect 28905 16099 28963 16105
rect 28905 16065 28917 16099
rect 28951 16096 28963 16099
rect 29012 16096 29040 16136
rect 30745 16133 30757 16167
rect 30791 16133 30803 16167
rect 30745 16127 30803 16133
rect 30834 16124 30840 16176
rect 30892 16164 30898 16176
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30892 16136 31033 16164
rect 30892 16124 30898 16136
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 31128 16136 31616 16164
rect 31128 16108 31156 16136
rect 28951 16068 29040 16096
rect 30561 16099 30619 16105
rect 28951 16065 28963 16068
rect 28905 16059 28963 16065
rect 30561 16065 30573 16099
rect 30607 16096 30619 16099
rect 30650 16096 30656 16108
rect 30607 16068 30656 16096
rect 30607 16065 30619 16068
rect 30561 16059 30619 16065
rect 30650 16056 30656 16068
rect 30708 16056 30714 16108
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16096 30987 16099
rect 31110 16096 31116 16108
rect 30975 16068 31116 16096
rect 30975 16065 30987 16068
rect 30929 16059 30987 16065
rect 31110 16056 31116 16068
rect 31168 16056 31174 16108
rect 31205 16099 31263 16105
rect 31205 16065 31217 16099
rect 31251 16096 31263 16099
rect 31294 16096 31300 16108
rect 31251 16068 31300 16096
rect 31251 16065 31263 16068
rect 31205 16059 31263 16065
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 31588 16105 31616 16136
rect 32892 16126 32920 16204
rect 32950 16192 32956 16204
rect 33008 16192 33014 16244
rect 33226 16192 33232 16244
rect 33284 16232 33290 16244
rect 33781 16235 33839 16241
rect 33781 16232 33793 16235
rect 33284 16204 33793 16232
rect 33284 16192 33290 16204
rect 33781 16201 33793 16204
rect 33827 16201 33839 16235
rect 33781 16195 33839 16201
rect 32953 16129 33011 16135
rect 32953 16126 32965 16129
rect 31573 16099 31631 16105
rect 31573 16065 31585 16099
rect 31619 16065 31631 16099
rect 31573 16059 31631 16065
rect 31757 16099 31815 16105
rect 31757 16065 31769 16099
rect 31803 16096 31815 16099
rect 32398 16096 32404 16108
rect 31803 16068 32404 16096
rect 31803 16065 31815 16068
rect 31757 16059 31815 16065
rect 32398 16056 32404 16068
rect 32456 16096 32462 16108
rect 32563 16099 32621 16105
rect 32563 16096 32575 16099
rect 32456 16068 32575 16096
rect 32456 16056 32462 16068
rect 32563 16065 32575 16068
rect 32609 16065 32621 16099
rect 32892 16098 32965 16126
rect 32953 16095 32965 16098
rect 32999 16095 33011 16129
rect 34517 16099 34575 16105
rect 34517 16096 34529 16099
rect 32953 16089 33011 16095
rect 32563 16059 32621 16065
rect 33704 16068 34529 16096
rect 26789 16031 26847 16037
rect 26789 15997 26801 16031
rect 26835 15997 26847 16031
rect 26789 15991 26847 15997
rect 26973 16031 27031 16037
rect 26973 15997 26985 16031
rect 27019 15997 27031 16031
rect 26973 15991 27031 15997
rect 28997 16031 29055 16037
rect 28997 15997 29009 16031
rect 29043 16028 29055 16031
rect 29362 16028 29368 16040
rect 29043 16000 29368 16028
rect 29043 15997 29055 16000
rect 28997 15991 29055 15997
rect 26988 15960 27016 15991
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 29914 15988 29920 16040
rect 29972 16028 29978 16040
rect 31386 16028 31392 16040
rect 29972 16000 31392 16028
rect 29972 15988 29978 16000
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 31478 15988 31484 16040
rect 31536 15988 31542 16040
rect 32306 15988 32312 16040
rect 32364 16028 32370 16040
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 32364 16000 32689 16028
rect 32364 15988 32370 16000
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 32677 15991 32735 15997
rect 26712 15932 27016 15960
rect 25498 15892 25504 15904
rect 25056 15864 25504 15892
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 26988 15892 27016 15932
rect 27982 15920 27988 15972
rect 28040 15960 28046 15972
rect 33704 15969 33732 16068
rect 34517 16065 34529 16068
rect 34563 16096 34575 16099
rect 37274 16096 37280 16108
rect 34563 16068 37280 16096
rect 34563 16065 34575 16068
rect 34517 16059 34575 16065
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 34793 16031 34851 16037
rect 34793 15997 34805 16031
rect 34839 15997 34851 16031
rect 34793 15991 34851 15997
rect 33689 15963 33747 15969
rect 28040 15932 29316 15960
rect 28040 15920 28046 15932
rect 29288 15904 29316 15932
rect 33689 15929 33701 15963
rect 33735 15929 33747 15963
rect 33689 15923 33747 15929
rect 28166 15892 28172 15904
rect 26988 15864 28172 15892
rect 28166 15852 28172 15864
rect 28224 15852 28230 15904
rect 29178 15852 29184 15904
rect 29236 15852 29242 15904
rect 29270 15852 29276 15904
rect 29328 15852 29334 15904
rect 31294 15852 31300 15904
rect 31352 15892 31358 15904
rect 32493 15895 32551 15901
rect 32493 15892 32505 15895
rect 31352 15864 32505 15892
rect 31352 15852 31358 15864
rect 32493 15861 32505 15864
rect 32539 15892 32551 15895
rect 33502 15892 33508 15904
rect 32539 15864 33508 15892
rect 32539 15861 32551 15864
rect 32493 15855 32551 15861
rect 33502 15852 33508 15864
rect 33560 15852 33566 15904
rect 33778 15852 33784 15904
rect 33836 15892 33842 15904
rect 34808 15892 34836 15991
rect 33836 15864 34836 15892
rect 33836 15852 33842 15864
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8018 15648 8024 15700
rect 8076 15688 8082 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 8076 15660 8401 15688
rect 8076 15648 8082 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 10410 15688 10416 15700
rect 8389 15651 8447 15657
rect 8588 15660 10416 15688
rect 8588 15493 8616 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 13722 15648 13728 15700
rect 13780 15648 13786 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 14918 15688 14924 15700
rect 14783 15660 14924 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 11057 15623 11115 15629
rect 11057 15589 11069 15623
rect 11103 15620 11115 15623
rect 11146 15620 11152 15632
rect 11103 15592 11152 15620
rect 11103 15589 11115 15592
rect 11057 15583 11115 15589
rect 11146 15580 11152 15592
rect 11204 15580 11210 15632
rect 14752 15620 14780 15651
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 27157 15691 27215 15697
rect 27157 15657 27169 15691
rect 27203 15688 27215 15691
rect 27203 15660 28580 15688
rect 27203 15657 27215 15660
rect 27157 15651 27215 15657
rect 28552 15632 28580 15660
rect 29178 15648 29184 15700
rect 29236 15648 29242 15700
rect 29270 15648 29276 15700
rect 29328 15688 29334 15700
rect 35434 15688 35440 15700
rect 29328 15660 35440 15688
rect 29328 15648 29334 15660
rect 35434 15648 35440 15660
rect 35492 15648 35498 15700
rect 13464 15592 14780 15620
rect 20257 15623 20315 15629
rect 10686 15512 10692 15564
rect 10744 15512 10750 15564
rect 11974 15512 11980 15564
rect 12032 15512 12038 15564
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 10008 15456 10149 15484
rect 10008 15444 10014 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 2774 15376 2780 15428
rect 2832 15376 2838 15428
rect 9876 15416 9904 15444
rect 10704 15416 10732 15512
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11572 15456 11897 15484
rect 11572 15444 11578 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 11992 15484 12020 15512
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 11992 15456 12081 15484
rect 11885 15447 11943 15453
rect 12069 15453 12081 15456
rect 12115 15484 12127 15487
rect 12158 15484 12164 15496
rect 12115 15456 12164 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 9876 15388 10732 15416
rect 11900 15416 11928 15447
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 13464 15493 13492 15592
rect 20257 15589 20269 15623
rect 20303 15620 20315 15623
rect 23293 15623 23351 15629
rect 23293 15620 23305 15623
rect 20303 15592 20668 15620
rect 20303 15589 20315 15592
rect 20257 15583 20315 15589
rect 20640 15564 20668 15592
rect 22066 15592 23305 15620
rect 22066 15564 22094 15592
rect 23293 15589 23305 15592
rect 23339 15589 23351 15623
rect 23293 15583 23351 15589
rect 28166 15580 28172 15632
rect 28224 15580 28230 15632
rect 28534 15580 28540 15632
rect 28592 15580 28598 15632
rect 13722 15512 13728 15564
rect 13780 15552 13786 15564
rect 13780 15524 14504 15552
rect 13780 15512 13786 15524
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13587 15487 13645 15493
rect 13587 15453 13599 15487
rect 13633 15484 13645 15487
rect 13633 15456 13768 15484
rect 13633 15453 13645 15456
rect 13587 15447 13645 15453
rect 11974 15416 11980 15428
rect 11900 15388 11980 15416
rect 11974 15376 11980 15388
rect 12032 15376 12038 15428
rect 13740 15416 13768 15456
rect 13814 15444 13820 15496
rect 13872 15484 13878 15496
rect 14476 15493 14504 15524
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15552 16911 15555
rect 17126 15552 17132 15564
rect 16899 15524 17132 15552
rect 16899 15521 16911 15524
rect 16853 15515 16911 15521
rect 17126 15512 17132 15524
rect 17184 15512 17190 15564
rect 20070 15512 20076 15564
rect 20128 15512 20134 15564
rect 20441 15555 20499 15561
rect 20441 15521 20453 15555
rect 20487 15521 20499 15555
rect 20441 15515 20499 15521
rect 13909 15487 13967 15493
rect 13909 15484 13921 15487
rect 13872 15456 13921 15484
rect 13872 15444 13878 15456
rect 13909 15453 13921 15456
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 14568 15416 14596 15512
rect 14734 15444 14740 15496
rect 14792 15444 14798 15496
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 16942 15484 16948 15496
rect 16807 15456 16948 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 16942 15444 16948 15456
rect 17000 15444 17006 15496
rect 20088 15484 20116 15512
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 20088 15456 20177 15484
rect 20165 15453 20177 15456
rect 20211 15453 20223 15487
rect 20456 15484 20484 15515
rect 20622 15512 20628 15564
rect 20680 15512 20686 15564
rect 22066 15552 22100 15564
rect 20916 15524 22100 15552
rect 20714 15484 20720 15496
rect 20456 15456 20720 15484
rect 20165 15447 20223 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 20916 15493 20944 15524
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 23750 15512 23756 15564
rect 23808 15512 23814 15564
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21039 15456 21588 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21266 15416 21272 15428
rect 13740 15388 14596 15416
rect 20456 15388 21272 15416
rect 2792 15348 2820 15376
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 2792 15320 9137 15348
rect 9125 15317 9137 15320
rect 9171 15348 9183 15351
rect 10042 15348 10048 15360
rect 9171 15320 10048 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 11146 15308 11152 15360
rect 11204 15308 11210 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 12124 15320 12265 15348
rect 12124 15308 12130 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 13906 15308 13912 15360
rect 13964 15308 13970 15360
rect 14918 15308 14924 15360
rect 14976 15308 14982 15360
rect 17129 15351 17187 15357
rect 17129 15317 17141 15351
rect 17175 15348 17187 15351
rect 17770 15348 17776 15360
rect 17175 15320 17776 15348
rect 17175 15317 17187 15320
rect 17129 15311 17187 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 20456 15357 20484 15388
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 21560 15360 21588 15456
rect 23566 15444 23572 15496
rect 23624 15444 23630 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 23842 15484 23848 15496
rect 23707 15456 23848 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 23842 15444 23848 15456
rect 23900 15484 23906 15496
rect 24394 15484 24400 15496
rect 23900 15456 24400 15484
rect 23900 15444 23906 15456
rect 24394 15444 24400 15456
rect 24452 15444 24458 15496
rect 27893 15487 27951 15493
rect 27893 15453 27905 15487
rect 27939 15484 27951 15487
rect 27982 15484 27988 15496
rect 27939 15456 27988 15484
rect 27939 15453 27951 15456
rect 27893 15447 27951 15453
rect 27982 15444 27988 15456
rect 28040 15444 28046 15496
rect 28184 15493 28212 15580
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 29196 15484 29224 15648
rect 30466 15580 30472 15632
rect 30524 15580 30530 15632
rect 31018 15580 31024 15632
rect 31076 15580 31082 15632
rect 32306 15580 32312 15632
rect 32364 15620 32370 15632
rect 33778 15620 33784 15632
rect 32364 15592 33784 15620
rect 32364 15580 32370 15592
rect 33778 15580 33784 15592
rect 33836 15580 33842 15632
rect 30944 15524 31340 15552
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29196 15456 29745 15484
rect 28169 15447 28227 15453
rect 29733 15453 29745 15456
rect 29779 15484 29791 15487
rect 30009 15487 30067 15493
rect 30009 15484 30021 15487
rect 29779 15456 30021 15484
rect 29779 15453 29791 15456
rect 29733 15447 29791 15453
rect 30009 15453 30021 15456
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 30193 15487 30251 15493
rect 30193 15453 30205 15487
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 23584 15416 23612 15444
rect 25225 15419 25283 15425
rect 25225 15416 25237 15419
rect 23584 15388 25237 15416
rect 25225 15385 25237 15388
rect 25271 15385 25283 15419
rect 25225 15379 25283 15385
rect 26973 15419 27031 15425
rect 26973 15385 26985 15419
rect 27019 15385 27031 15419
rect 26973 15379 27031 15385
rect 20441 15351 20499 15357
rect 20441 15317 20453 15351
rect 20487 15317 20499 15351
rect 20441 15311 20499 15317
rect 20530 15308 20536 15360
rect 20588 15308 20594 15360
rect 21542 15308 21548 15360
rect 21600 15308 21606 15360
rect 25590 15308 25596 15360
rect 25648 15348 25654 15360
rect 26988 15348 27016 15379
rect 27246 15376 27252 15428
rect 27304 15416 27310 15428
rect 28258 15416 28264 15428
rect 27304 15388 28264 15416
rect 27304 15376 27310 15388
rect 28258 15376 28264 15388
rect 28316 15376 28322 15428
rect 29454 15416 29460 15428
rect 28368 15388 29460 15416
rect 27522 15348 27528 15360
rect 25648 15320 27528 15348
rect 25648 15308 25654 15320
rect 27522 15308 27528 15320
rect 27580 15348 27586 15360
rect 28368 15348 28396 15388
rect 29454 15376 29460 15388
rect 29512 15376 29518 15428
rect 29549 15419 29607 15425
rect 29549 15385 29561 15419
rect 29595 15416 29607 15419
rect 30208 15416 30236 15447
rect 30650 15444 30656 15496
rect 30708 15444 30714 15496
rect 30944 15493 30972 15524
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15453 30987 15487
rect 30929 15447 30987 15453
rect 31021 15487 31079 15493
rect 31021 15453 31033 15487
rect 31067 15453 31079 15487
rect 31021 15447 31079 15453
rect 29595 15388 30236 15416
rect 30668 15416 30696 15444
rect 31036 15416 31064 15447
rect 31312 15425 31340 15524
rect 30668 15388 31064 15416
rect 31113 15419 31171 15425
rect 29595 15385 29607 15388
rect 29549 15379 29607 15385
rect 31113 15385 31125 15419
rect 31159 15385 31171 15419
rect 31113 15379 31171 15385
rect 31297 15419 31355 15425
rect 31297 15385 31309 15419
rect 31343 15416 31355 15419
rect 31570 15416 31576 15428
rect 31343 15388 31576 15416
rect 31343 15385 31355 15388
rect 31297 15379 31355 15385
rect 27580 15320 28396 15348
rect 28721 15351 28779 15357
rect 27580 15308 27586 15320
rect 28721 15317 28733 15351
rect 28767 15348 28779 15351
rect 28994 15348 29000 15360
rect 28767 15320 29000 15348
rect 28767 15317 28779 15320
rect 28721 15311 28779 15317
rect 28994 15308 29000 15320
rect 29052 15348 29058 15360
rect 29564 15348 29592 15379
rect 29052 15320 29592 15348
rect 29052 15308 29058 15320
rect 29914 15308 29920 15360
rect 29972 15308 29978 15360
rect 30098 15308 30104 15360
rect 30156 15308 30162 15360
rect 30837 15351 30895 15357
rect 30837 15317 30849 15351
rect 30883 15348 30895 15351
rect 31128 15348 31156 15379
rect 31570 15376 31576 15388
rect 31628 15376 31634 15428
rect 31478 15348 31484 15360
rect 30883 15320 31484 15348
rect 30883 15317 30895 15320
rect 30837 15311 30895 15317
rect 31478 15308 31484 15320
rect 31536 15308 31542 15360
rect 1104 15258 38824 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 38824 15258
rect 1104 15184 38824 15206
rect 14734 15104 14740 15156
rect 14792 15104 14798 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 18509 15147 18567 15153
rect 18509 15144 18521 15147
rect 18472 15116 18521 15144
rect 18472 15104 18478 15116
rect 18509 15113 18521 15116
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 22189 15147 22247 15153
rect 22189 15144 22201 15147
rect 21876 15116 22201 15144
rect 21876 15104 21882 15116
rect 22189 15113 22201 15116
rect 22235 15113 22247 15147
rect 22189 15107 22247 15113
rect 25866 15104 25872 15156
rect 25924 15104 25930 15156
rect 26418 15104 26424 15156
rect 26476 15104 26482 15156
rect 26973 15147 27031 15153
rect 26973 15113 26985 15147
rect 27019 15113 27031 15147
rect 26973 15107 27031 15113
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11701 15079 11759 15085
rect 11701 15076 11713 15079
rect 11204 15048 11713 15076
rect 11204 15036 11210 15048
rect 11701 15045 11713 15048
rect 11747 15045 11759 15079
rect 11701 15039 11759 15045
rect 17313 15079 17371 15085
rect 17313 15045 17325 15079
rect 17359 15076 17371 15079
rect 18598 15076 18604 15088
rect 17359 15048 18604 15076
rect 17359 15045 17371 15048
rect 17313 15039 17371 15045
rect 18598 15036 18604 15048
rect 18656 15076 18662 15088
rect 21177 15079 21235 15085
rect 21177 15076 21189 15079
rect 18656 15048 20208 15076
rect 18656 15036 18662 15048
rect 11514 14968 11520 15020
rect 11572 14968 11578 15020
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14139 14980 14381 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14001 14943 14059 14949
rect 14001 14940 14013 14943
rect 13964 14912 14013 14940
rect 13964 14900 13970 14912
rect 14001 14909 14013 14912
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 13722 14832 13728 14884
rect 13780 14832 13786 14884
rect 14108 14816 14136 14971
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14516 14980 14565 15008
rect 14516 14968 14522 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 16942 14968 16948 15020
rect 17000 15008 17006 15020
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 17000 14980 17049 15008
rect 17000 14968 17006 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 18233 15011 18291 15017
rect 18233 15008 18245 15011
rect 17037 14971 17095 14977
rect 17604 14980 18245 15008
rect 17604 14952 17632 14980
rect 18233 14977 18245 14980
rect 18279 14977 18291 15011
rect 18233 14971 18291 14977
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 20180 15017 20208 15048
rect 20456 15048 21189 15076
rect 20456 15017 20484 15048
rect 21177 15045 21189 15048
rect 21223 15045 21235 15079
rect 21177 15039 21235 15045
rect 21361 15079 21419 15085
rect 21361 15045 21373 15079
rect 21407 15076 21419 15079
rect 22094 15076 22100 15088
rect 21407 15048 22100 15076
rect 21407 15045 21419 15048
rect 21361 15039 21419 15045
rect 22094 15036 22100 15048
rect 22152 15036 22158 15088
rect 23566 15036 23572 15088
rect 23624 15076 23630 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 23624 15048 23673 15076
rect 23624 15036 23630 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 24794 15048 25697 15076
rect 23661 15039 23719 15045
rect 25685 15045 25697 15048
rect 25731 15045 25743 15079
rect 26988 15076 27016 15107
rect 27246 15104 27252 15156
rect 27304 15144 27310 15156
rect 27433 15147 27491 15153
rect 27433 15144 27445 15147
rect 27304 15116 27445 15144
rect 27304 15104 27310 15116
rect 27433 15113 27445 15116
rect 27479 15113 27491 15147
rect 27433 15107 27491 15113
rect 27540 15116 30052 15144
rect 25685 15039 25743 15045
rect 26068 15048 27016 15076
rect 20165 15011 20223 15017
rect 20165 14977 20177 15011
rect 20211 14977 20223 15011
rect 20165 14971 20223 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 15010 14900 15016 14952
rect 15068 14900 15074 14952
rect 16666 14900 16672 14952
rect 16724 14900 16730 14952
rect 17126 14900 17132 14952
rect 17184 14900 17190 14952
rect 17586 14900 17592 14952
rect 17644 14900 17650 14952
rect 17681 14943 17739 14949
rect 17681 14909 17693 14943
rect 17727 14909 17739 14943
rect 17681 14903 17739 14909
rect 15028 14872 15056 14900
rect 17696 14872 17724 14903
rect 17770 14900 17776 14952
rect 17828 14900 17834 14952
rect 17862 14900 17868 14952
rect 17920 14900 17926 14952
rect 17954 14900 17960 14952
rect 18012 14900 18018 14952
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14940 18567 14943
rect 19702 14940 19708 14952
rect 18555 14912 19708 14940
rect 18555 14909 18567 14912
rect 18509 14903 18567 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 15028 14844 17724 14872
rect 17788 14872 17816 14900
rect 19150 14872 19156 14884
rect 17788 14844 19156 14872
rect 19150 14832 19156 14844
rect 19208 14832 19214 14884
rect 11885 14807 11943 14813
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 12986 14804 12992 14816
rect 11931 14776 12992 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 14090 14764 14096 14816
rect 14148 14764 14154 14816
rect 18141 14807 18199 14813
rect 18141 14773 18153 14807
rect 18187 14804 18199 14807
rect 18325 14807 18383 14813
rect 18325 14804 18337 14807
rect 18187 14776 18337 14804
rect 18187 14773 18199 14776
rect 18141 14767 18199 14773
rect 18325 14773 18337 14776
rect 18371 14773 18383 14807
rect 18325 14767 18383 14773
rect 19610 14764 19616 14816
rect 19668 14804 19674 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19668 14776 19809 14804
rect 19668 14764 19674 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 20088 14804 20116 14968
rect 20272 14940 20300 14971
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20640 14980 20729 15008
rect 20548 14940 20576 14968
rect 20272 14912 20576 14940
rect 20640 14804 20668 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 21542 14968 21548 15020
rect 21600 14968 21606 15020
rect 25501 15011 25559 15017
rect 25501 14977 25513 15011
rect 25547 15008 25559 15011
rect 25590 15008 25596 15020
rect 25547 14980 25596 15008
rect 25547 14977 25559 14980
rect 25501 14971 25559 14977
rect 25590 14968 25596 14980
rect 25648 14968 25654 15020
rect 26068 15017 26096 15048
rect 25777 15011 25835 15017
rect 25777 14977 25789 15011
rect 25823 14977 25835 15011
rect 25777 14971 25835 14977
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 14977 26111 15011
rect 26053 14971 26111 14977
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 15008 26571 15011
rect 26559 14980 27292 15008
rect 26559 14977 26571 14980
rect 26513 14971 26571 14977
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 20732 14912 20821 14940
rect 20732 14816 20760 14912
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 20809 14903 20867 14909
rect 23566 14900 23572 14952
rect 23624 14940 23630 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 23624 14912 25237 14940
rect 23624 14900 23630 14912
rect 25225 14909 25237 14912
rect 25271 14909 25283 14943
rect 25792 14940 25820 14971
rect 25225 14903 25283 14909
rect 25700 14912 25820 14940
rect 23198 14832 23204 14884
rect 23256 14872 23262 14884
rect 23256 14844 24256 14872
rect 23256 14832 23262 14844
rect 20088 14776 20668 14804
rect 19797 14767 19855 14773
rect 20714 14764 20720 14816
rect 20772 14764 20778 14816
rect 21082 14764 21088 14816
rect 21140 14764 21146 14816
rect 21358 14764 21364 14816
rect 21416 14804 21422 14816
rect 22278 14804 22284 14816
rect 21416 14776 22284 14804
rect 21416 14764 21422 14776
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23750 14764 23756 14816
rect 23808 14764 23814 14816
rect 24228 14804 24256 14844
rect 25700 14804 25728 14912
rect 24228 14776 25728 14804
rect 27264 14804 27292 14980
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 27540 14952 27568 15116
rect 30024 15088 30052 15116
rect 30098 15104 30104 15156
rect 30156 15104 30162 15156
rect 27706 15036 27712 15088
rect 27764 15076 27770 15088
rect 27985 15079 28043 15085
rect 27985 15076 27997 15079
rect 27764 15048 27997 15076
rect 27764 15036 27770 15048
rect 27985 15045 27997 15048
rect 28031 15076 28043 15079
rect 28534 15076 28540 15088
rect 28031 15048 28540 15076
rect 28031 15045 28043 15048
rect 27985 15039 28043 15045
rect 28534 15036 28540 15048
rect 28592 15036 28598 15088
rect 30006 15036 30012 15088
rect 30064 15036 30070 15088
rect 28813 15011 28871 15017
rect 28813 15008 28825 15011
rect 28460 14980 28825 15008
rect 27522 14900 27528 14952
rect 27580 14900 27586 14952
rect 28460 14949 28488 14980
rect 28813 14977 28825 14980
rect 28859 14977 28871 15011
rect 28813 14971 28871 14977
rect 28994 14968 29000 15020
rect 29052 14968 29058 15020
rect 29914 14968 29920 15020
rect 29972 14968 29978 15020
rect 30116 15017 30144 15104
rect 30101 15011 30159 15017
rect 30101 14977 30113 15011
rect 30147 14977 30159 15011
rect 30101 14971 30159 14977
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 28718 14900 28724 14952
rect 28776 14940 28782 14952
rect 29638 14940 29644 14952
rect 28776 14912 29644 14940
rect 28776 14900 28782 14912
rect 29638 14900 29644 14912
rect 29696 14900 29702 14952
rect 30009 14943 30067 14949
rect 30009 14909 30021 14943
rect 30055 14940 30067 14943
rect 30650 14940 30656 14952
rect 30055 14912 30656 14940
rect 30055 14909 30067 14912
rect 30009 14903 30067 14909
rect 30650 14900 30656 14912
rect 30708 14900 30714 14952
rect 28258 14832 28264 14884
rect 28316 14832 28322 14884
rect 28350 14832 28356 14884
rect 28408 14872 28414 14884
rect 28902 14872 28908 14884
rect 28408 14844 28908 14872
rect 28408 14832 28414 14844
rect 28902 14832 28908 14844
rect 28960 14832 28966 14884
rect 28368 14804 28396 14832
rect 27264 14776 28396 14804
rect 28810 14764 28816 14816
rect 28868 14764 28874 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 14090 14600 14096 14612
rect 12406 14572 14096 14600
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14464 9643 14467
rect 10042 14464 10048 14476
rect 9631 14436 10048 14464
rect 9631 14433 9643 14436
rect 9585 14427 9643 14433
rect 10042 14424 10048 14436
rect 10100 14464 10106 14476
rect 10318 14464 10324 14476
rect 10100 14436 10324 14464
rect 10100 14424 10106 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 11514 14424 11520 14476
rect 11572 14424 11578 14476
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14464 12311 14467
rect 12406 14464 12434 14572
rect 14090 14560 14096 14572
rect 14148 14600 14154 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 14148 14572 14197 14600
rect 14148 14560 14154 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 16724 14572 16773 14600
rect 16724 14560 16730 14572
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 16761 14563 16819 14569
rect 17586 14560 17592 14612
rect 17644 14560 17650 14612
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 18049 14603 18107 14609
rect 18049 14600 18061 14603
rect 18012 14572 18061 14600
rect 18012 14560 18018 14572
rect 18049 14569 18061 14572
rect 18095 14569 18107 14603
rect 18049 14563 18107 14569
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20070 14560 20076 14612
rect 20128 14560 20134 14612
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21140 14572 22094 14600
rect 21140 14560 21146 14572
rect 13722 14492 13728 14544
rect 13780 14492 13786 14544
rect 14918 14492 14924 14544
rect 14976 14492 14982 14544
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 19334 14532 19340 14544
rect 15252 14504 15976 14532
rect 15252 14492 15258 14504
rect 13740 14464 13768 14492
rect 12299 14436 12434 14464
rect 13004 14436 13768 14464
rect 14936 14464 14964 14492
rect 14936 14436 15884 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8619 14368 8984 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 8956 14269 8984 14368
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 11204 14368 11437 14396
rect 11204 14356 11210 14368
rect 11425 14365 11437 14368
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 12618 14356 12624 14408
rect 12676 14396 12682 14408
rect 13004 14405 13032 14436
rect 12805 14399 12863 14405
rect 12805 14396 12817 14399
rect 12676 14368 12817 14396
rect 12676 14356 12682 14368
rect 12805 14365 12817 14368
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13170 14356 13176 14408
rect 13228 14356 13234 14408
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13964 14368 14105 14396
rect 13964 14356 13970 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14936 14396 14964 14436
rect 15105 14399 15163 14405
rect 15105 14396 15117 14399
rect 14936 14368 15117 14396
rect 14093 14359 14151 14365
rect 15105 14365 15117 14368
rect 15151 14365 15163 14399
rect 15105 14359 15163 14365
rect 15194 14356 15200 14408
rect 15252 14356 15258 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15746 14396 15752 14408
rect 15427 14368 15752 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 15856 14405 15884 14436
rect 15948 14405 15976 14504
rect 16224 14504 19340 14532
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15933 14399 15991 14405
rect 15933 14365 15945 14399
rect 15979 14365 15991 14399
rect 15933 14359 15991 14365
rect 16114 14356 16120 14408
rect 16172 14356 16178 14408
rect 16224 14405 16252 14504
rect 19334 14492 19340 14504
rect 19392 14532 19398 14544
rect 19613 14535 19671 14541
rect 19613 14532 19625 14535
rect 19392 14504 19625 14532
rect 19392 14492 19398 14504
rect 19613 14501 19625 14504
rect 19659 14501 19671 14535
rect 19613 14495 19671 14501
rect 19996 14532 20024 14560
rect 21821 14535 21879 14541
rect 21821 14532 21833 14535
rect 19996 14504 21833 14532
rect 16942 14424 16948 14476
rect 17000 14424 17006 14476
rect 17954 14424 17960 14476
rect 18012 14424 18018 14476
rect 19889 14467 19947 14473
rect 18248 14436 19472 14464
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17126 14396 17132 14408
rect 17083 14368 17132 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14396 17463 14399
rect 17451 14368 17724 14396
rect 17451 14365 17463 14368
rect 17405 14359 17463 14365
rect 17696 14340 17724 14368
rect 17770 14356 17776 14408
rect 17828 14356 17834 14408
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14396 17923 14399
rect 17972 14396 18000 14424
rect 18248 14408 18276 14436
rect 17911 14368 18000 14396
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 18432 14368 18521 14396
rect 9324 14300 12434 14328
rect 9324 14269 9352 14300
rect 8389 14263 8447 14269
rect 8389 14260 8401 14263
rect 8352 14232 8401 14260
rect 8352 14220 8358 14232
rect 8389 14229 8401 14232
rect 8435 14229 8447 14263
rect 8389 14223 8447 14229
rect 8941 14263 8999 14269
rect 8941 14229 8953 14263
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14229 9367 14263
rect 9309 14223 9367 14229
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 9674 14260 9680 14272
rect 9447 14232 9680 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 12406 14260 12434 14300
rect 12894 14288 12900 14340
rect 12952 14288 12958 14340
rect 14826 14328 14832 14340
rect 13004 14300 14832 14328
rect 13004 14272 13032 14300
rect 14826 14288 14832 14300
rect 14884 14288 14890 14340
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 15611 14300 17264 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 12621 14263 12679 14269
rect 12621 14260 12633 14263
rect 12406 14232 12633 14260
rect 12621 14229 12633 14232
rect 12667 14229 12679 14263
rect 12621 14223 12679 14229
rect 12986 14220 12992 14272
rect 13044 14220 13050 14272
rect 14550 14220 14556 14272
rect 14608 14220 14614 14272
rect 15654 14220 15660 14272
rect 15712 14220 15718 14272
rect 17236 14260 17264 14300
rect 17310 14288 17316 14340
rect 17368 14288 17374 14340
rect 17586 14288 17592 14340
rect 17644 14288 17650 14340
rect 17678 14288 17684 14340
rect 17736 14288 17742 14340
rect 18432 14328 18460 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 18598 14356 18604 14408
rect 18656 14356 18662 14408
rect 19058 14356 19064 14408
rect 19116 14356 19122 14408
rect 19150 14356 19156 14408
rect 19208 14396 19214 14408
rect 19444 14405 19472 14436
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 19996 14464 20024 14504
rect 19935 14436 20024 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 19208 14368 19257 14396
rect 19208 14356 19214 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19429 14399 19487 14405
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 18969 14331 19027 14337
rect 18432 14300 18828 14328
rect 18800 14272 18828 14300
rect 18969 14297 18981 14331
rect 19015 14328 19027 14331
rect 19337 14331 19395 14337
rect 19337 14328 19349 14331
rect 19015 14300 19349 14328
rect 19015 14297 19027 14300
rect 18969 14291 19027 14297
rect 19337 14297 19349 14300
rect 19383 14328 19395 14331
rect 20180 14328 20208 14359
rect 19383 14300 20208 14328
rect 19383 14297 19395 14300
rect 19337 14291 19395 14297
rect 18414 14260 18420 14272
rect 17236 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18782 14220 18788 14272
rect 18840 14220 18846 14272
rect 18877 14263 18935 14269
rect 18877 14229 18889 14263
rect 18923 14260 18935 14263
rect 20622 14260 20628 14272
rect 18923 14232 20628 14260
rect 18923 14229 18935 14232
rect 18877 14223 18935 14229
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 21468 14260 21496 14504
rect 21821 14501 21833 14504
rect 21867 14501 21879 14535
rect 22066 14532 22094 14572
rect 22462 14560 22468 14612
rect 22520 14560 22526 14612
rect 26142 14600 26148 14612
rect 23032 14572 26148 14600
rect 22066 14504 22784 14532
rect 21821 14495 21879 14501
rect 21542 14424 21548 14476
rect 21600 14464 21606 14476
rect 22097 14467 22155 14473
rect 22097 14464 22109 14467
rect 21600 14436 22109 14464
rect 21600 14424 21606 14436
rect 22097 14433 22109 14436
rect 22143 14433 22155 14467
rect 22097 14427 22155 14433
rect 22189 14399 22247 14405
rect 22189 14396 22201 14399
rect 22112 14368 22201 14396
rect 22112 14340 22140 14368
rect 22189 14365 22201 14368
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22278 14356 22284 14408
rect 22336 14356 22342 14408
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 22649 14399 22707 14405
rect 22649 14396 22661 14399
rect 22428 14368 22661 14396
rect 22428 14356 22434 14368
rect 22649 14365 22661 14368
rect 22695 14365 22707 14399
rect 22756 14396 22784 14504
rect 23032 14408 23060 14572
rect 26142 14560 26148 14572
rect 26200 14600 26206 14612
rect 26878 14600 26884 14612
rect 26200 14572 26884 14600
rect 26200 14560 26206 14572
rect 26878 14560 26884 14572
rect 26936 14560 26942 14612
rect 27249 14603 27307 14609
rect 27249 14569 27261 14603
rect 27295 14600 27307 14603
rect 27338 14600 27344 14612
rect 27295 14572 27344 14600
rect 27295 14569 27307 14572
rect 27249 14563 27307 14569
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 28810 14560 28816 14612
rect 28868 14560 28874 14612
rect 28997 14603 29055 14609
rect 28997 14569 29009 14603
rect 29043 14600 29055 14603
rect 29086 14600 29092 14612
rect 29043 14572 29092 14600
rect 29043 14569 29055 14572
rect 28997 14563 29055 14569
rect 29086 14560 29092 14572
rect 29144 14560 29150 14612
rect 29178 14560 29184 14612
rect 29236 14600 29242 14612
rect 29730 14600 29736 14612
rect 29236 14572 29736 14600
rect 29236 14560 29242 14572
rect 29730 14560 29736 14572
rect 29788 14560 29794 14612
rect 31110 14560 31116 14612
rect 31168 14560 31174 14612
rect 31570 14560 31576 14612
rect 31628 14560 31634 14612
rect 27433 14535 27491 14541
rect 27433 14501 27445 14535
rect 27479 14532 27491 14535
rect 28718 14532 28724 14544
rect 27479 14504 28724 14532
rect 27479 14501 27491 14504
rect 27433 14495 27491 14501
rect 28718 14492 28724 14504
rect 28776 14492 28782 14544
rect 28828 14532 28856 14560
rect 28828 14504 32076 14532
rect 23290 14424 23296 14476
rect 23348 14464 23354 14476
rect 23474 14464 23480 14476
rect 23348 14436 23480 14464
rect 23348 14424 23354 14436
rect 23474 14424 23480 14436
rect 23532 14464 23538 14476
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23532 14436 23857 14464
rect 23532 14424 23538 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 28626 14464 28632 14476
rect 23845 14427 23903 14433
rect 26804 14436 28632 14464
rect 22833 14399 22891 14405
rect 22833 14396 22845 14399
rect 22756 14368 22845 14396
rect 22649 14359 22707 14365
rect 22833 14365 22845 14368
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 23014 14356 23020 14408
rect 23072 14356 23078 14408
rect 24394 14356 24400 14408
rect 24452 14356 24458 14408
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 24912 14368 25237 14396
rect 24912 14356 24918 14368
rect 25225 14365 25237 14368
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 22094 14288 22100 14340
rect 22152 14288 22158 14340
rect 22296 14328 22324 14356
rect 22738 14328 22744 14340
rect 22296 14300 22744 14328
rect 22738 14288 22744 14300
rect 22796 14288 22802 14340
rect 25240 14328 25268 14359
rect 25498 14356 25504 14408
rect 25556 14356 25562 14408
rect 26804 14405 26832 14436
rect 28626 14424 28632 14436
rect 28684 14424 28690 14476
rect 30929 14467 30987 14473
rect 30929 14464 30941 14467
rect 28828 14436 30941 14464
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14365 26847 14399
rect 26789 14359 26847 14365
rect 26878 14356 26884 14408
rect 26936 14356 26942 14408
rect 27062 14356 27068 14408
rect 27120 14356 27126 14408
rect 27617 14399 27675 14405
rect 27617 14396 27629 14399
rect 27540 14368 27629 14396
rect 25240 14300 27292 14328
rect 27264 14272 27292 14300
rect 27540 14272 27568 14368
rect 27617 14365 27629 14368
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14365 27767 14399
rect 27709 14359 27767 14365
rect 27893 14399 27951 14405
rect 27893 14365 27905 14399
rect 27939 14365 27951 14399
rect 27893 14359 27951 14365
rect 27724 14328 27752 14359
rect 27632 14300 27752 14328
rect 27632 14272 27660 14300
rect 22186 14260 22192 14272
rect 21468 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 23290 14220 23296 14272
rect 23348 14220 23354 14272
rect 23658 14220 23664 14272
rect 23716 14220 23722 14272
rect 23750 14220 23756 14272
rect 23808 14220 23814 14272
rect 27246 14220 27252 14272
rect 27304 14220 27310 14272
rect 27522 14220 27528 14272
rect 27580 14220 27586 14272
rect 27614 14220 27620 14272
rect 27672 14220 27678 14272
rect 27908 14260 27936 14359
rect 27982 14356 27988 14408
rect 28040 14356 28046 14408
rect 28629 14331 28687 14337
rect 28629 14297 28641 14331
rect 28675 14328 28687 14331
rect 28718 14328 28724 14340
rect 28675 14300 28724 14328
rect 28675 14297 28687 14300
rect 28629 14291 28687 14297
rect 28718 14288 28724 14300
rect 28776 14288 28782 14340
rect 28828 14337 28856 14436
rect 30929 14433 30941 14436
rect 30975 14433 30987 14467
rect 30929 14427 30987 14433
rect 31404 14436 31708 14464
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14365 30251 14399
rect 30193 14359 30251 14365
rect 28813 14331 28871 14337
rect 28813 14297 28825 14331
rect 28859 14297 28871 14331
rect 28813 14291 28871 14297
rect 28828 14260 28856 14291
rect 27908 14232 28856 14260
rect 28902 14220 28908 14272
rect 28960 14260 28966 14272
rect 30208 14260 30236 14359
rect 30834 14356 30840 14408
rect 30892 14396 30898 14408
rect 31404 14405 31432 14436
rect 31680 14405 31708 14436
rect 32048 14408 32076 14504
rect 32122 14492 32128 14544
rect 32180 14532 32186 14544
rect 32677 14535 32735 14541
rect 32677 14532 32689 14535
rect 32180 14504 32689 14532
rect 32180 14492 32186 14504
rect 32232 14473 32260 14504
rect 32677 14501 32689 14504
rect 32723 14501 32735 14535
rect 32677 14495 32735 14501
rect 32217 14467 32275 14473
rect 32217 14433 32229 14467
rect 32263 14433 32275 14467
rect 32217 14427 32275 14433
rect 32490 14424 32496 14476
rect 32548 14424 32554 14476
rect 32784 14436 35664 14464
rect 31389 14399 31447 14405
rect 30892 14368 31340 14396
rect 30892 14356 30898 14368
rect 31312 14328 31340 14368
rect 31389 14365 31401 14399
rect 31435 14365 31447 14399
rect 31389 14359 31447 14365
rect 31481 14399 31539 14405
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31665 14399 31723 14405
rect 31665 14396 31677 14399
rect 31623 14368 31677 14396
rect 31481 14359 31539 14365
rect 31665 14365 31677 14368
rect 31711 14396 31723 14399
rect 31846 14396 31852 14408
rect 31711 14368 31852 14396
rect 31711 14365 31723 14368
rect 31665 14359 31723 14365
rect 31496 14328 31524 14359
rect 31846 14356 31852 14368
rect 31904 14356 31910 14408
rect 32030 14356 32036 14408
rect 32088 14396 32094 14408
rect 32125 14399 32183 14405
rect 32125 14396 32137 14399
rect 32088 14368 32137 14396
rect 32088 14356 32094 14368
rect 32125 14365 32137 14368
rect 32171 14396 32183 14399
rect 32585 14399 32643 14405
rect 32585 14396 32597 14399
rect 32171 14368 32597 14396
rect 32171 14365 32183 14368
rect 32125 14359 32183 14365
rect 32585 14365 32597 14368
rect 32631 14365 32643 14399
rect 32585 14359 32643 14365
rect 31312 14300 31524 14328
rect 31570 14288 31576 14340
rect 31628 14328 31634 14340
rect 32784 14328 32812 14436
rect 35636 14408 35664 14436
rect 32861 14399 32919 14405
rect 32861 14365 32873 14399
rect 32907 14365 32919 14399
rect 32861 14359 32919 14365
rect 31628 14300 32812 14328
rect 31628 14288 31634 14300
rect 28960 14232 30236 14260
rect 30285 14263 30343 14269
rect 28960 14220 28966 14232
rect 30285 14229 30297 14263
rect 30331 14260 30343 14263
rect 30374 14260 30380 14272
rect 30331 14232 30380 14260
rect 30331 14229 30343 14232
rect 30285 14223 30343 14229
rect 30374 14220 30380 14232
rect 30432 14220 30438 14272
rect 31386 14220 31392 14272
rect 31444 14260 31450 14272
rect 32876 14260 32904 14359
rect 35618 14356 35624 14408
rect 35676 14356 35682 14408
rect 31444 14232 32904 14260
rect 31444 14220 31450 14232
rect 33042 14220 33048 14272
rect 33100 14220 33106 14272
rect 1104 14170 38824 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 38824 14170
rect 1104 14096 38824 14118
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 8938 14056 8944 14068
rect 7800 14028 8944 14056
rect 7800 14016 7806 14028
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9674 14056 9680 14068
rect 9539 14028 9680 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11514 14056 11520 14068
rect 11379 14028 11520 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14056 12403 14059
rect 12618 14056 12624 14068
rect 12391 14028 12624 14056
rect 12391 14025 12403 14028
rect 12345 14019 12403 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13814 14016 13820 14068
rect 13872 14016 13878 14068
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 14148 14028 14228 14056
rect 14148 14016 14154 14028
rect 7760 13929 7788 14016
rect 8021 13991 8079 13997
rect 8021 13957 8033 13991
rect 8067 13988 8079 13991
rect 8294 13988 8300 14000
rect 8067 13960 8300 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8662 13948 8668 14000
rect 8720 13948 8726 14000
rect 9692 13988 9720 14016
rect 13832 13988 13860 14016
rect 9692 13960 11008 13988
rect 13832 13960 14136 13988
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9858 13920 9864 13932
rect 9723 13892 9864 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10980 13929 11008 13960
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13889 11023 13923
rect 10965 13883 11023 13889
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 11977 13923 12035 13929
rect 11977 13920 11989 13923
rect 11940 13892 11989 13920
rect 11940 13880 11946 13892
rect 11977 13889 11989 13892
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 13998 13880 14004 13932
rect 14056 13880 14062 13932
rect 14108 13929 14136 13960
rect 14200 13929 14228 14028
rect 14918 14016 14924 14068
rect 14976 14016 14982 14068
rect 15654 14016 15660 14068
rect 15712 14016 15718 14068
rect 17770 14016 17776 14068
rect 17828 14016 17834 14068
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19058 14056 19064 14068
rect 18739 14028 19064 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19610 14016 19616 14068
rect 19668 14016 19674 14068
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 19760 14028 20821 14056
rect 19760 14016 19766 14028
rect 20809 14025 20821 14028
rect 20855 14025 20867 14059
rect 20809 14019 20867 14025
rect 23290 14016 23296 14068
rect 23348 14016 23354 14068
rect 23566 14016 23572 14068
rect 23624 14016 23630 14068
rect 23658 14016 23664 14068
rect 23716 14016 23722 14068
rect 27062 14016 27068 14068
rect 27120 14016 27126 14068
rect 27246 14016 27252 14068
rect 27304 14056 27310 14068
rect 27304 14028 31340 14056
rect 27304 14016 27310 14028
rect 14458 13988 14464 14000
rect 14292 13960 14464 13988
rect 14292 13929 14320 13960
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 14936 13988 14964 14016
rect 14936 13960 15424 13988
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14921 13923 14979 13929
rect 14921 13920 14933 13923
rect 14323 13892 14933 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 14921 13889 14933 13892
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 15396 13929 15424 13960
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10704 13824 11069 13852
rect 10704 13793 10732 13824
rect 11057 13821 11069 13824
rect 11103 13852 11115 13855
rect 11900 13852 11928 13880
rect 11103 13824 11928 13852
rect 11103 13821 11115 13824
rect 11057 13815 11115 13821
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 14550 13852 14556 13864
rect 14292 13824 14556 13852
rect 10689 13787 10747 13793
rect 10689 13753 10701 13787
rect 10735 13753 10747 13787
rect 10689 13747 10747 13753
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 14292 13716 14320 13824
rect 14550 13812 14556 13824
rect 14608 13852 14614 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14608 13824 14749 13852
rect 14608 13812 14614 13824
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 14826 13812 14832 13864
rect 14884 13812 14890 13864
rect 14461 13787 14519 13793
rect 14461 13753 14473 13787
rect 14507 13784 14519 13787
rect 15212 13784 15240 13880
rect 15672 13852 15700 14016
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17368 13960 18092 13988
rect 17368 13948 17374 13960
rect 17604 13929 17632 13960
rect 18064 13932 18092 13960
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17770 13880 17776 13932
rect 17828 13880 17834 13932
rect 18046 13880 18052 13932
rect 18104 13880 18110 13932
rect 18432 13920 18460 14016
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 18432 13892 18613 13920
rect 18601 13889 18613 13892
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18782 13880 18788 13932
rect 18840 13920 18846 13932
rect 19628 13929 19656 14016
rect 19904 13960 23244 13988
rect 19613 13923 19671 13929
rect 18840 13892 19472 13920
rect 18840 13880 18846 13892
rect 15672 13824 19288 13852
rect 14507 13756 15240 13784
rect 19260 13784 19288 13824
rect 19334 13812 19340 13864
rect 19392 13812 19398 13864
rect 19444 13861 19472 13892
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19904 13852 19932 13960
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22572 13892 22845 13920
rect 19429 13815 19487 13821
rect 19536 13824 19932 13852
rect 19536 13784 19564 13824
rect 20806 13812 20812 13864
rect 20864 13812 20870 13864
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 21324 13824 22109 13852
rect 21324 13812 21330 13824
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 22572 13793 22600 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13920 22983 13923
rect 23014 13920 23020 13932
rect 22971 13892 23020 13920
rect 22971 13889 22983 13892
rect 22925 13883 22983 13889
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 23106 13880 23112 13932
rect 23164 13880 23170 13932
rect 19260 13756 19564 13784
rect 19797 13787 19855 13793
rect 14507 13753 14519 13756
rect 14461 13747 14519 13753
rect 19797 13753 19809 13787
rect 19843 13784 19855 13787
rect 22557 13787 22615 13793
rect 19843 13756 22094 13784
rect 19843 13753 19855 13756
rect 19797 13747 19855 13753
rect 13320 13688 14320 13716
rect 13320 13676 13326 13688
rect 14550 13676 14556 13728
rect 14608 13676 14614 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 14884 13688 15301 13716
rect 14884 13676 14890 13688
rect 15289 13685 15301 13688
rect 15335 13685 15347 13719
rect 15289 13679 15347 13685
rect 20990 13676 20996 13728
rect 21048 13676 21054 13728
rect 22066 13716 22094 13756
rect 22557 13753 22569 13787
rect 22603 13753 22615 13787
rect 23216 13784 23244 13960
rect 23308 13920 23336 14016
rect 23385 13923 23443 13929
rect 23385 13920 23397 13923
rect 23308 13892 23397 13920
rect 23385 13889 23397 13892
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13852 23351 13855
rect 23676 13852 23704 14016
rect 27522 13988 27528 14000
rect 25608 13960 27528 13988
rect 25608 13932 25636 13960
rect 27522 13948 27528 13960
rect 27580 13988 27586 14000
rect 29546 13988 29552 14000
rect 27580 13960 27844 13988
rect 27580 13948 27586 13960
rect 23750 13880 23756 13932
rect 23808 13920 23814 13932
rect 24857 13923 24915 13929
rect 24857 13920 24869 13923
rect 23808 13892 24869 13920
rect 23808 13880 23814 13892
rect 24857 13889 24869 13892
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25424 13852 25452 13883
rect 25590 13880 25596 13932
rect 25648 13880 25654 13932
rect 27246 13880 27252 13932
rect 27304 13880 27310 13932
rect 27614 13920 27620 13932
rect 27356 13892 27620 13920
rect 27356 13852 27384 13892
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 27816 13929 27844 13960
rect 28000 13960 29552 13988
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 23339 13824 23704 13852
rect 23768 13824 27384 13852
rect 23339 13821 23351 13824
rect 23293 13815 23351 13821
rect 23768 13784 23796 13824
rect 27430 13812 27436 13864
rect 27488 13852 27494 13864
rect 27525 13855 27583 13861
rect 27525 13852 27537 13855
rect 27488 13824 27537 13852
rect 27488 13812 27494 13824
rect 27525 13821 27537 13824
rect 27571 13852 27583 13855
rect 28000 13852 28028 13960
rect 29546 13948 29552 13960
rect 29604 13948 29610 14000
rect 29730 13948 29736 14000
rect 29788 13988 29794 14000
rect 30009 13991 30067 13997
rect 30009 13988 30021 13991
rect 29788 13960 30021 13988
rect 29788 13948 29794 13960
rect 30009 13957 30021 13960
rect 30055 13957 30067 13991
rect 30009 13951 30067 13957
rect 30101 13991 30159 13997
rect 30101 13957 30113 13991
rect 30147 13988 30159 13991
rect 31312 13988 31340 14028
rect 31478 14016 31484 14068
rect 31536 14016 31542 14068
rect 31570 14016 31576 14068
rect 31628 14016 31634 14068
rect 31849 14059 31907 14065
rect 31849 14025 31861 14059
rect 31895 14056 31907 14059
rect 32030 14056 32036 14068
rect 31895 14028 32036 14056
rect 31895 14025 31907 14028
rect 31849 14019 31907 14025
rect 32030 14016 32036 14028
rect 32088 14016 32094 14068
rect 33042 14016 33048 14068
rect 33100 14016 33106 14068
rect 31588 13988 31616 14016
rect 33060 13988 33088 14016
rect 30147 13960 31248 13988
rect 31312 13960 31616 13988
rect 31680 13960 33088 13988
rect 30147 13957 30159 13960
rect 30101 13951 30159 13957
rect 31220 13932 31248 13960
rect 28442 13920 28448 13932
rect 27571 13824 28028 13852
rect 28092 13892 28448 13920
rect 27571 13821 27583 13824
rect 27525 13815 27583 13821
rect 25590 13784 25596 13796
rect 23216 13756 23796 13784
rect 24872 13756 25596 13784
rect 22557 13747 22615 13753
rect 24872 13716 24900 13756
rect 25590 13744 25596 13756
rect 25648 13744 25654 13796
rect 26970 13744 26976 13796
rect 27028 13784 27034 13796
rect 28092 13784 28120 13892
rect 28442 13880 28448 13892
rect 28500 13920 28506 13932
rect 28500 13892 29224 13920
rect 28500 13880 28506 13892
rect 28626 13812 28632 13864
rect 28684 13852 28690 13864
rect 29196 13852 29224 13892
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 29871 13923 29929 13929
rect 29871 13920 29883 13923
rect 29328 13892 29883 13920
rect 29328 13880 29334 13892
rect 29871 13889 29883 13892
rect 29917 13889 29929 13923
rect 29871 13883 29929 13889
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13920 30251 13923
rect 30558 13920 30564 13932
rect 30239 13892 30564 13920
rect 30239 13889 30251 13892
rect 30193 13883 30251 13889
rect 30558 13880 30564 13892
rect 30616 13880 30622 13932
rect 31202 13880 31208 13932
rect 31260 13880 31266 13932
rect 31386 13880 31392 13932
rect 31444 13880 31450 13932
rect 31680 13929 31708 13960
rect 31665 13923 31723 13929
rect 31665 13889 31677 13923
rect 31711 13889 31723 13923
rect 31665 13883 31723 13889
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13920 31999 13923
rect 32030 13920 32036 13932
rect 31987 13892 32036 13920
rect 31987 13889 31999 13892
rect 31941 13883 31999 13889
rect 32030 13880 32036 13892
rect 32088 13880 32094 13932
rect 32214 13880 32220 13932
rect 32272 13920 32278 13932
rect 32490 13920 32496 13932
rect 32272 13892 32496 13920
rect 32272 13880 32278 13892
rect 32490 13880 32496 13892
rect 32548 13880 32554 13932
rect 29733 13855 29791 13861
rect 29733 13852 29745 13855
rect 28684 13824 29132 13852
rect 29196 13824 29745 13852
rect 28684 13812 28690 13824
rect 27028 13756 28120 13784
rect 29104 13784 29132 13824
rect 29733 13821 29745 13824
rect 29779 13821 29791 13855
rect 31297 13855 31355 13861
rect 29733 13815 29791 13821
rect 29840 13824 31248 13852
rect 29840 13784 29868 13824
rect 29104 13756 29868 13784
rect 31220 13784 31248 13824
rect 31297 13821 31309 13855
rect 31343 13852 31355 13855
rect 32401 13855 32459 13861
rect 32401 13852 32413 13855
rect 31343 13824 32413 13852
rect 31343 13821 31355 13824
rect 31297 13815 31355 13821
rect 32401 13821 32413 13824
rect 32447 13821 32459 13855
rect 32401 13815 32459 13821
rect 32125 13787 32183 13793
rect 32125 13784 32137 13787
rect 31220 13756 32137 13784
rect 27028 13744 27034 13756
rect 32125 13753 32137 13756
rect 32171 13753 32183 13787
rect 32125 13747 32183 13753
rect 22066 13688 24900 13716
rect 24946 13676 24952 13728
rect 25004 13676 25010 13728
rect 25498 13676 25504 13728
rect 25556 13676 25562 13728
rect 27433 13719 27491 13725
rect 27433 13685 27445 13719
rect 27479 13716 27491 13719
rect 27614 13716 27620 13728
rect 27479 13688 27620 13716
rect 27479 13685 27491 13688
rect 27433 13679 27491 13685
rect 27614 13676 27620 13688
rect 27672 13676 27678 13728
rect 27890 13676 27896 13728
rect 27948 13716 27954 13728
rect 27985 13719 28043 13725
rect 27985 13716 27997 13719
rect 27948 13688 27997 13716
rect 27948 13676 27954 13688
rect 27985 13685 27997 13688
rect 28031 13685 28043 13719
rect 27985 13679 28043 13685
rect 30377 13719 30435 13725
rect 30377 13685 30389 13719
rect 30423 13716 30435 13719
rect 30466 13716 30472 13728
rect 30423 13688 30472 13716
rect 30423 13685 30435 13688
rect 30377 13679 30435 13685
rect 30466 13676 30472 13688
rect 30524 13676 30530 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 4062 13472 4068 13524
rect 4120 13472 4126 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 9950 13512 9956 13524
rect 9048 13484 9956 13512
rect 4080 13444 4108 13472
rect 9048 13453 9076 13484
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 13722 13512 13728 13524
rect 13004 13484 13728 13512
rect 13004 13456 13032 13484
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13814 13472 13820 13524
rect 13872 13472 13878 13524
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 13998 13512 14004 13524
rect 13955 13484 14004 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14185 13515 14243 13521
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 14458 13512 14464 13524
rect 14231 13484 14464 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 18230 13472 18236 13524
rect 18288 13472 18294 13524
rect 22370 13512 22376 13524
rect 22020 13484 22376 13512
rect 9033 13447 9091 13453
rect 9033 13444 9045 13447
rect 4080 13416 9045 13444
rect 9033 13413 9045 13416
rect 9079 13413 9091 13447
rect 9033 13407 9091 13413
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 11882 13444 11888 13456
rect 11287 13416 11888 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 12986 13404 12992 13456
rect 13044 13404 13050 13456
rect 13354 13404 13360 13456
rect 13412 13404 13418 13456
rect 13832 13444 13860 13472
rect 22020 13453 22048 13484
rect 22370 13472 22376 13484
rect 22428 13472 22434 13524
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23293 13515 23351 13521
rect 23293 13512 23305 13515
rect 23164 13484 23305 13512
rect 23164 13472 23170 13484
rect 23293 13481 23305 13484
rect 23339 13481 23351 13515
rect 27246 13512 27252 13524
rect 23293 13475 23351 13481
rect 24228 13484 27252 13512
rect 15105 13447 15163 13453
rect 15105 13444 15117 13447
rect 13832 13416 15117 13444
rect 15105 13413 15117 13416
rect 15151 13413 15163 13447
rect 15105 13407 15163 13413
rect 22005 13447 22063 13453
rect 22005 13413 22017 13447
rect 22051 13413 22063 13447
rect 22005 13407 22063 13413
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 14553 13379 14611 13385
rect 11379 13348 13860 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 8772 13240 8800 13271
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9732 13280 9781 13308
rect 9732 13268 9738 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 9122 13240 9128 13252
rect 8772 13212 9128 13240
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9784 13240 9812 13271
rect 9858 13268 9864 13320
rect 9916 13308 9922 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9916 13280 10057 13308
rect 9916 13268 9922 13280
rect 10045 13277 10057 13280
rect 10091 13308 10103 13311
rect 10318 13308 10324 13320
rect 10091 13280 10324 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 13262 13308 13268 13320
rect 13127 13280 13268 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13556 13317 13584 13348
rect 13541 13311 13599 13317
rect 13452 13289 13510 13295
rect 10873 13243 10931 13249
rect 10873 13240 10885 13243
rect 9784 13212 10885 13240
rect 10873 13209 10885 13212
rect 10919 13209 10931 13243
rect 10873 13203 10931 13209
rect 12250 13200 12256 13252
rect 12308 13200 12314 13252
rect 12437 13243 12495 13249
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 12894 13240 12900 13252
rect 12483 13212 12900 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 13004 13240 13032 13268
rect 13452 13255 13464 13289
rect 13498 13255 13510 13289
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 13722 13268 13728 13320
rect 13780 13268 13786 13320
rect 13832 13308 13860 13348
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 14599 13348 15056 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13832 13280 14473 13308
rect 14461 13277 14473 13280
rect 14507 13308 14519 13311
rect 14921 13311 14979 13317
rect 14921 13308 14933 13311
rect 14507 13280 14933 13308
rect 14507 13277 14519 13280
rect 14461 13271 14519 13277
rect 14921 13277 14933 13280
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 13452 13252 13510 13255
rect 13173 13243 13231 13249
rect 13173 13240 13185 13243
rect 13004 13212 13185 13240
rect 13173 13209 13185 13212
rect 13219 13209 13231 13243
rect 13173 13203 13231 13209
rect 13357 13243 13415 13249
rect 13357 13209 13369 13243
rect 13403 13209 13415 13243
rect 13357 13203 13415 13209
rect 13372 13172 13400 13203
rect 13446 13200 13452 13252
rect 13504 13240 13510 13252
rect 14737 13243 14795 13249
rect 14737 13240 14749 13243
rect 13504 13212 14749 13240
rect 13504 13200 13510 13212
rect 14737 13209 14749 13212
rect 14783 13240 14795 13243
rect 15028 13240 15056 13348
rect 18046 13336 18052 13388
rect 18104 13336 18110 13388
rect 21082 13336 21088 13388
rect 21140 13376 21146 13388
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 21140 13348 21557 13376
rect 21140 13336 21146 13348
rect 21545 13345 21557 13348
rect 21591 13345 21603 13379
rect 24228 13376 24256 13484
rect 27246 13472 27252 13484
rect 27304 13472 27310 13524
rect 27525 13515 27583 13521
rect 27525 13481 27537 13515
rect 27571 13512 27583 13515
rect 27614 13512 27620 13524
rect 27571 13484 27620 13512
rect 27571 13481 27583 13484
rect 27525 13475 27583 13481
rect 27614 13472 27620 13484
rect 27672 13472 27678 13524
rect 27982 13472 27988 13524
rect 28040 13512 28046 13524
rect 28077 13515 28135 13521
rect 28077 13512 28089 13515
rect 28040 13484 28089 13512
rect 28040 13472 28046 13484
rect 28077 13481 28089 13484
rect 28123 13481 28135 13515
rect 28077 13475 28135 13481
rect 28169 13515 28227 13521
rect 28169 13481 28181 13515
rect 28215 13512 28227 13515
rect 30834 13512 30840 13524
rect 28215 13484 30840 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 31202 13472 31208 13524
rect 31260 13512 31266 13524
rect 31481 13515 31539 13521
rect 31481 13512 31493 13515
rect 31260 13484 31493 13512
rect 31260 13472 31266 13484
rect 31481 13481 31493 13484
rect 31527 13481 31539 13515
rect 31481 13475 31539 13481
rect 31846 13472 31852 13524
rect 31904 13472 31910 13524
rect 24302 13404 24308 13456
rect 24360 13444 24366 13456
rect 24360 13416 25360 13444
rect 24360 13404 24366 13416
rect 21545 13339 21603 13345
rect 22756 13348 24256 13376
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 17770 13308 17776 13320
rect 17276 13280 17776 13308
rect 17276 13268 17282 13280
rect 17770 13268 17776 13280
rect 17828 13308 17834 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17828 13280 17969 13308
rect 17828 13268 17834 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 18064 13308 18092 13336
rect 22756 13320 22784 13348
rect 23124 13320 23152 13348
rect 24394 13336 24400 13388
rect 24452 13376 24458 13388
rect 24673 13379 24731 13385
rect 24673 13376 24685 13379
rect 24452 13348 24685 13376
rect 24452 13336 24458 13348
rect 24673 13345 24685 13348
rect 24719 13345 24731 13379
rect 24673 13339 24731 13345
rect 21266 13308 21272 13320
rect 18064 13280 21272 13308
rect 17957 13271 18015 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21637 13311 21695 13317
rect 21637 13277 21649 13311
rect 21683 13308 21695 13311
rect 22094 13308 22100 13320
rect 21683 13280 22100 13308
rect 21683 13277 21695 13280
rect 21637 13271 21695 13277
rect 22094 13268 22100 13280
rect 22152 13308 22158 13320
rect 22554 13308 22560 13320
rect 22152 13280 22560 13308
rect 22152 13268 22158 13280
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 22738 13268 22744 13320
rect 22796 13268 22802 13320
rect 22830 13268 22836 13320
rect 22888 13268 22894 13320
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23106 13268 23112 13320
rect 23164 13268 23170 13320
rect 14783 13212 15056 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 19702 13200 19708 13252
rect 19760 13240 19766 13252
rect 22756 13240 22784 13268
rect 19760 13212 22784 13240
rect 24688 13240 24716 13339
rect 24946 13336 24952 13388
rect 25004 13336 25010 13388
rect 24762 13268 24768 13320
rect 24820 13268 24826 13320
rect 24964 13308 24992 13336
rect 25332 13317 25360 13416
rect 28261 13379 28319 13385
rect 28261 13345 28273 13379
rect 28307 13376 28319 13379
rect 30852 13376 30880 13472
rect 28307 13348 28764 13376
rect 30852 13348 31432 13376
rect 28307 13345 28319 13348
rect 28261 13339 28319 13345
rect 28736 13320 28764 13348
rect 25225 13311 25283 13317
rect 25225 13308 25237 13311
rect 24964 13280 25237 13308
rect 25225 13277 25237 13280
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 25317 13311 25375 13317
rect 25317 13277 25329 13311
rect 25363 13277 25375 13311
rect 25317 13271 25375 13277
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 27525 13311 27583 13317
rect 27525 13277 27537 13311
rect 27571 13308 27583 13311
rect 27706 13308 27712 13320
rect 27571 13280 27712 13308
rect 27571 13277 27583 13280
rect 27525 13271 27583 13277
rect 25516 13240 25544 13271
rect 27706 13268 27712 13280
rect 27764 13268 27770 13320
rect 27798 13268 27804 13320
rect 27856 13268 27862 13320
rect 27890 13268 27896 13320
rect 27948 13308 27954 13320
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 27948 13280 27997 13308
rect 27948 13268 27954 13280
rect 27985 13277 27997 13280
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28000 13240 28028 13271
rect 28718 13268 28724 13320
rect 28776 13268 28782 13320
rect 29546 13268 29552 13320
rect 29604 13268 29610 13320
rect 31404 13317 31432 13348
rect 32214 13336 32220 13388
rect 32272 13336 32278 13388
rect 31389 13311 31447 13317
rect 31389 13277 31401 13311
rect 31435 13277 31447 13311
rect 31389 13271 31447 13277
rect 31573 13311 31631 13317
rect 31573 13277 31585 13311
rect 31619 13308 31631 13311
rect 31938 13308 31944 13320
rect 31619 13280 31944 13308
rect 31619 13277 31631 13280
rect 31573 13271 31631 13277
rect 31938 13268 31944 13280
rect 31996 13308 32002 13320
rect 32033 13311 32091 13317
rect 32033 13308 32045 13311
rect 31996 13280 32045 13308
rect 31996 13268 32002 13280
rect 32033 13277 32045 13280
rect 32079 13277 32091 13311
rect 32033 13271 32091 13277
rect 28074 13240 28080 13252
rect 24688 13212 25544 13240
rect 27632 13212 28080 13240
rect 19760 13200 19766 13212
rect 27632 13184 27660 13212
rect 28074 13200 28080 13212
rect 28132 13200 28138 13252
rect 29822 13200 29828 13252
rect 29880 13200 29886 13252
rect 30374 13200 30380 13252
rect 30432 13200 30438 13252
rect 31312 13212 31754 13240
rect 14458 13172 14464 13184
rect 13372 13144 14464 13172
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 25130 13132 25136 13184
rect 25188 13132 25194 13184
rect 25682 13132 25688 13184
rect 25740 13132 25746 13184
rect 27614 13132 27620 13184
rect 27672 13132 27678 13184
rect 27709 13175 27767 13181
rect 27709 13141 27721 13175
rect 27755 13172 27767 13175
rect 27890 13172 27896 13184
rect 27755 13144 27896 13172
rect 27755 13141 27767 13144
rect 27709 13135 27767 13141
rect 27890 13132 27896 13144
rect 27948 13132 27954 13184
rect 30098 13132 30104 13184
rect 30156 13172 30162 13184
rect 31312 13181 31340 13212
rect 31726 13184 31754 13212
rect 31297 13175 31355 13181
rect 31297 13172 31309 13175
rect 30156 13144 31309 13172
rect 30156 13132 30162 13144
rect 31297 13141 31309 13144
rect 31343 13141 31355 13175
rect 31726 13144 31760 13184
rect 31297 13135 31355 13141
rect 31754 13132 31760 13144
rect 31812 13132 31818 13184
rect 1104 13082 38824 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 38824 13082
rect 1104 13008 38824 13030
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12342 12968 12348 12980
rect 12032 12940 12348 12968
rect 12032 12928 12038 12940
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12584 12940 12633 12968
rect 12584 12928 12590 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 12894 12928 12900 12980
rect 12952 12928 12958 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 9769 12903 9827 12909
rect 9769 12869 9781 12903
rect 9815 12900 9827 12903
rect 13096 12900 13124 12931
rect 13354 12928 13360 12980
rect 13412 12928 13418 12980
rect 14550 12928 14556 12980
rect 14608 12928 14614 12980
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 17184 12940 17325 12968
rect 17184 12928 17190 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21183 12971 21241 12977
rect 21183 12968 21195 12971
rect 21048 12940 21195 12968
rect 21048 12928 21054 12940
rect 21183 12937 21195 12940
rect 21229 12937 21241 12971
rect 21183 12931 21241 12937
rect 22554 12928 22560 12980
rect 22612 12928 22618 12980
rect 22734 12971 22792 12977
rect 22734 12937 22746 12971
rect 22780 12968 22792 12971
rect 22922 12968 22928 12980
rect 22780 12940 22928 12968
rect 22780 12937 22792 12940
rect 22734 12931 22792 12937
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 24762 12928 24768 12980
rect 24820 12928 24826 12980
rect 24946 12928 24952 12980
rect 25004 12928 25010 12980
rect 25590 12928 25596 12980
rect 25648 12968 25654 12980
rect 27617 12971 27675 12977
rect 27617 12968 27629 12971
rect 25648 12940 27629 12968
rect 25648 12928 25654 12940
rect 27617 12937 27629 12940
rect 27663 12937 27675 12971
rect 27617 12931 27675 12937
rect 27706 12928 27712 12980
rect 27764 12928 27770 12980
rect 27982 12928 27988 12980
rect 28040 12968 28046 12980
rect 28353 12971 28411 12977
rect 28353 12968 28365 12971
rect 28040 12940 28365 12968
rect 28040 12928 28046 12940
rect 28353 12937 28365 12940
rect 28399 12937 28411 12971
rect 28353 12931 28411 12937
rect 29270 12928 29276 12980
rect 29328 12928 29334 12980
rect 29549 12971 29607 12977
rect 29549 12937 29561 12971
rect 29595 12968 29607 12971
rect 29822 12968 29828 12980
rect 29595 12940 29828 12968
rect 29595 12937 29607 12940
rect 29549 12931 29607 12937
rect 29822 12928 29828 12940
rect 29880 12928 29886 12980
rect 30009 12971 30067 12977
rect 30009 12937 30021 12971
rect 30055 12968 30067 12971
rect 30466 12968 30472 12980
rect 30055 12940 30472 12968
rect 30055 12937 30067 12940
rect 30009 12931 30067 12937
rect 30466 12928 30472 12940
rect 30524 12928 30530 12980
rect 13372 12900 13400 12928
rect 9815 12872 13124 12900
rect 13280 12872 13400 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 12529 12835 12587 12841
rect 12529 12832 12541 12835
rect 11808 12804 12541 12832
rect 11808 12776 11836 12804
rect 12529 12801 12541 12804
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 9858 12724 9864 12776
rect 9916 12724 9922 12776
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 11882 12724 11888 12776
rect 11940 12724 11946 12776
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12158 12764 12164 12776
rect 12115 12736 12164 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 12158 12724 12164 12736
rect 12216 12764 12222 12776
rect 12728 12764 12756 12795
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 13280 12841 13308 12872
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 14568 12832 14596 12928
rect 21085 12903 21143 12909
rect 20640 12872 20944 12900
rect 13403 12804 14596 12832
rect 15657 12835 15715 12841
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 15657 12801 15669 12835
rect 15703 12832 15715 12835
rect 16666 12832 16672 12844
rect 15703 12804 16672 12832
rect 15703 12801 15715 12804
rect 15657 12795 15715 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 17773 12835 17831 12841
rect 17773 12832 17785 12835
rect 16908 12804 17785 12832
rect 16908 12792 16914 12804
rect 17773 12801 17785 12804
rect 17819 12801 17831 12835
rect 17773 12795 17831 12801
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 18288 12804 18797 12832
rect 18288 12792 18294 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 19794 12792 19800 12844
rect 19852 12832 19858 12844
rect 20530 12832 20536 12844
rect 19852 12804 20536 12832
rect 19852 12792 19858 12804
rect 20530 12792 20536 12804
rect 20588 12832 20594 12844
rect 20640 12841 20668 12872
rect 20916 12866 20944 12872
rect 21085 12869 21097 12903
rect 21131 12869 21143 12903
rect 22572 12900 22600 12928
rect 22649 12903 22707 12909
rect 22649 12900 22661 12903
rect 22572 12872 22661 12900
rect 21085 12866 21143 12869
rect 20916 12863 21143 12866
rect 22649 12869 22661 12872
rect 22695 12869 22707 12903
rect 22833 12903 22891 12909
rect 22833 12900 22845 12903
rect 22649 12863 22707 12869
rect 22756 12872 22845 12900
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20588 12804 20637 12832
rect 20588 12792 20594 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 20806 12792 20812 12844
rect 20864 12792 20870 12844
rect 20916 12838 21128 12863
rect 22756 12844 22784 12872
rect 22833 12869 22845 12872
rect 22879 12900 22891 12903
rect 24302 12900 24308 12912
rect 22879 12872 24308 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 24302 12860 24308 12872
rect 24360 12860 24366 12912
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 12216 12736 12756 12764
rect 12820 12764 12848 12792
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 12820 12736 13645 12764
rect 12216 12724 12222 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 13722 12724 13728 12776
rect 13780 12724 13786 12776
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12764 17003 12767
rect 18877 12767 18935 12773
rect 16991 12736 17448 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 11900 12696 11928 12724
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 11900 12668 12357 12696
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 12345 12659 12403 12665
rect 17218 12656 17224 12708
rect 17276 12656 17282 12708
rect 17420 12705 17448 12736
rect 18877 12733 18889 12767
rect 18923 12764 18935 12767
rect 19058 12764 19064 12776
rect 18923 12736 19064 12764
rect 18923 12733 18935 12736
rect 18877 12727 18935 12733
rect 19058 12724 19064 12736
rect 19116 12724 19122 12776
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 18414 12696 18420 12708
rect 17451 12668 18420 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 19153 12699 19211 12705
rect 19153 12665 19165 12699
rect 19199 12696 19211 12699
rect 19794 12696 19800 12708
rect 19199 12668 19800 12696
rect 19199 12665 19211 12668
rect 19153 12659 19211 12665
rect 19794 12656 19800 12668
rect 19852 12656 19858 12708
rect 20806 12656 20812 12708
rect 20864 12696 20870 12708
rect 21284 12696 21312 12795
rect 21358 12792 21364 12844
rect 21416 12792 21422 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22066 12804 22569 12832
rect 20864 12668 21312 12696
rect 20864 12656 20870 12668
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8904 12600 9413 12628
rect 8904 12588 8910 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12434 12628 12440 12640
rect 12299 12600 12440 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 20990 12588 20996 12640
rect 21048 12588 21054 12640
rect 21082 12588 21088 12640
rect 21140 12628 21146 12640
rect 22066 12628 22094 12804
rect 22557 12801 22569 12804
rect 22603 12801 22615 12835
rect 22557 12795 22615 12801
rect 22738 12792 22744 12844
rect 22796 12792 22802 12844
rect 24320 12832 24348 12860
rect 24762 12832 24768 12844
rect 24320 12804 24768 12832
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 24964 12841 24992 12928
rect 25222 12860 25228 12912
rect 25280 12900 25286 12912
rect 25682 12900 25688 12912
rect 25280 12872 25688 12900
rect 25280 12860 25286 12872
rect 25682 12860 25688 12872
rect 25740 12860 25746 12912
rect 27341 12903 27399 12909
rect 27341 12869 27353 12903
rect 27387 12900 27399 12903
rect 27430 12900 27436 12912
rect 27387 12872 27436 12900
rect 27387 12869 27399 12872
rect 27341 12863 27399 12869
rect 27430 12860 27436 12872
rect 27488 12860 27494 12912
rect 30098 12860 30104 12912
rect 30156 12860 30162 12912
rect 30653 12903 30711 12909
rect 30653 12869 30665 12903
rect 30699 12900 30711 12903
rect 31938 12900 31944 12912
rect 30699 12872 31944 12900
rect 30699 12869 30711 12872
rect 30653 12863 30711 12869
rect 31938 12860 31944 12872
rect 31996 12860 32002 12912
rect 32030 12860 32036 12912
rect 32088 12900 32094 12912
rect 32088 12872 32352 12900
rect 32088 12860 32094 12872
rect 24949 12835 25007 12841
rect 24949 12801 24961 12835
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 25130 12792 25136 12844
rect 25188 12832 25194 12844
rect 25317 12835 25375 12841
rect 25188 12804 25268 12832
rect 25188 12792 25194 12804
rect 25240 12773 25268 12804
rect 25317 12801 25329 12835
rect 25363 12832 25375 12835
rect 25498 12832 25504 12844
rect 25363 12804 25504 12832
rect 25363 12801 25375 12804
rect 25317 12795 25375 12801
rect 25498 12792 25504 12804
rect 25556 12792 25562 12844
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12764 25283 12767
rect 25958 12764 25964 12776
rect 25271 12736 25964 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 25958 12724 25964 12736
rect 26016 12764 26022 12776
rect 26145 12767 26203 12773
rect 26145 12764 26157 12767
rect 26016 12736 26157 12764
rect 26016 12724 26022 12736
rect 26145 12733 26157 12736
rect 26191 12733 26203 12767
rect 26252 12764 26280 12795
rect 27522 12792 27528 12844
rect 27580 12792 27586 12844
rect 27982 12792 27988 12844
rect 28040 12792 28046 12844
rect 28166 12792 28172 12844
rect 28224 12792 28230 12844
rect 28905 12835 28963 12841
rect 28905 12801 28917 12835
rect 28951 12801 28963 12835
rect 28905 12795 28963 12801
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12832 29423 12835
rect 29411 12804 29684 12832
rect 29411 12801 29423 12804
rect 29365 12795 29423 12801
rect 27614 12764 27620 12776
rect 26252 12736 27620 12764
rect 26145 12727 26203 12733
rect 27614 12724 27620 12736
rect 27672 12724 27678 12776
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28258 12764 28264 12776
rect 27856 12736 28264 12764
rect 27856 12724 27862 12736
rect 28258 12724 28264 12736
rect 28316 12764 28322 12776
rect 28813 12767 28871 12773
rect 28813 12764 28825 12767
rect 28316 12736 28825 12764
rect 28316 12724 28322 12736
rect 28813 12733 28825 12736
rect 28859 12733 28871 12767
rect 28813 12727 28871 12733
rect 28920 12764 28948 12795
rect 29454 12764 29460 12776
rect 28920 12736 29460 12764
rect 25866 12656 25872 12708
rect 25924 12656 25930 12708
rect 27890 12656 27896 12708
rect 27948 12696 27954 12708
rect 28920 12696 28948 12736
rect 29454 12724 29460 12736
rect 29512 12724 29518 12776
rect 29656 12705 29684 12804
rect 30834 12792 30840 12844
rect 30892 12792 30898 12844
rect 32122 12792 32128 12844
rect 32180 12792 32186 12844
rect 32324 12841 32352 12872
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12832 32367 12835
rect 32582 12832 32588 12844
rect 32355 12804 32588 12832
rect 32355 12801 32367 12804
rect 32309 12795 32367 12801
rect 32582 12792 32588 12804
rect 32640 12792 32646 12844
rect 30190 12724 30196 12776
rect 30248 12724 30254 12776
rect 30469 12767 30527 12773
rect 30469 12733 30481 12767
rect 30515 12764 30527 12767
rect 30558 12764 30564 12776
rect 30515 12736 30564 12764
rect 30515 12733 30527 12736
rect 30469 12727 30527 12733
rect 30558 12724 30564 12736
rect 30616 12724 30622 12776
rect 27948 12668 28948 12696
rect 29641 12699 29699 12705
rect 27948 12656 27954 12668
rect 29641 12665 29653 12699
rect 29687 12665 29699 12699
rect 29641 12659 29699 12665
rect 21140 12600 22094 12628
rect 21140 12588 21146 12600
rect 25038 12588 25044 12640
rect 25096 12588 25102 12640
rect 31846 12588 31852 12640
rect 31904 12628 31910 12640
rect 32493 12631 32551 12637
rect 32493 12628 32505 12631
rect 31904 12600 32505 12628
rect 31904 12588 31910 12600
rect 32493 12597 32505 12600
rect 32539 12597 32551 12631
rect 32493 12591 32551 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 12250 12384 12256 12436
rect 12308 12424 12314 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12308 12396 12633 12424
rect 12308 12384 12314 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13722 12424 13728 12436
rect 13035 12396 13728 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 16761 12427 16819 12433
rect 16761 12393 16773 12427
rect 16807 12424 16819 12427
rect 16850 12424 16856 12436
rect 16807 12396 16856 12424
rect 16807 12393 16819 12396
rect 16761 12387 16819 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 18322 12424 18328 12436
rect 16960 12396 18328 12424
rect 12345 12359 12403 12365
rect 12345 12325 12357 12359
rect 12391 12356 12403 12359
rect 13446 12356 13452 12368
rect 12391 12328 13452 12356
rect 12391 12325 12403 12328
rect 12345 12319 12403 12325
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11848 12260 11897 12288
rect 11848 12248 11854 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 15286 12248 15292 12300
rect 15344 12248 15350 12300
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8846 12220 8852 12232
rect 8619 12192 8852 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 10704 12192 11989 12220
rect 9217 12155 9275 12161
rect 9217 12152 9229 12155
rect 8772 12124 9229 12152
rect 8772 12093 8800 12124
rect 9217 12121 9229 12124
rect 9263 12121 9275 12155
rect 9217 12115 9275 12121
rect 9674 12112 9680 12164
rect 9732 12112 9738 12164
rect 10704 12096 10732 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12526 12180 12532 12232
rect 12584 12180 12590 12232
rect 13630 12180 13636 12232
rect 13688 12220 13694 12232
rect 15010 12220 15016 12232
rect 13688 12192 15016 12220
rect 13688 12180 13694 12192
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 16298 12112 16304 12164
rect 16356 12112 16362 12164
rect 16868 12152 16896 12384
rect 16960 12297 16988 12396
rect 18064 12297 18092 12396
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 19061 12427 19119 12433
rect 19061 12424 19073 12427
rect 18472 12396 19073 12424
rect 18472 12384 18478 12396
rect 19061 12393 19073 12396
rect 19107 12424 19119 12427
rect 19107 12396 19334 12424
rect 19107 12393 19119 12396
rect 19061 12387 19119 12393
rect 16945 12291 17003 12297
rect 16945 12257 16957 12291
rect 16991 12257 17003 12291
rect 16945 12251 17003 12257
rect 18049 12291 18107 12297
rect 18049 12257 18061 12291
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 17221 12223 17279 12229
rect 17221 12189 17233 12223
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 18371 12192 18736 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 17126 12152 17132 12164
rect 16868 12124 17132 12152
rect 17126 12112 17132 12124
rect 17184 12152 17190 12164
rect 17236 12152 17264 12183
rect 17184 12124 17264 12152
rect 17184 12112 17190 12124
rect 18708 12096 18736 12192
rect 19306 12152 19334 12396
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21358 12424 21364 12436
rect 20772 12396 21364 12424
rect 20772 12384 20778 12396
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 22738 12384 22744 12436
rect 22796 12384 22802 12436
rect 22922 12384 22928 12436
rect 22980 12424 22986 12436
rect 25498 12424 25504 12436
rect 22980 12396 25504 12424
rect 22980 12384 22986 12396
rect 25498 12384 25504 12396
rect 25556 12384 25562 12436
rect 26050 12384 26056 12436
rect 26108 12424 26114 12436
rect 27154 12424 27160 12436
rect 26108 12396 27160 12424
rect 26108 12384 26114 12396
rect 27154 12384 27160 12396
rect 27212 12424 27218 12436
rect 28810 12424 28816 12436
rect 27212 12396 28816 12424
rect 27212 12384 27218 12396
rect 28810 12384 28816 12396
rect 28868 12384 28874 12436
rect 31297 12427 31355 12433
rect 31297 12393 31309 12427
rect 31343 12424 31355 12427
rect 31386 12424 31392 12436
rect 31343 12396 31392 12424
rect 31343 12393 31355 12396
rect 31297 12387 31355 12393
rect 31386 12384 31392 12396
rect 31444 12384 31450 12436
rect 31941 12427 31999 12433
rect 31941 12393 31953 12427
rect 31987 12424 31999 12427
rect 32122 12424 32128 12436
rect 31987 12396 32128 12424
rect 31987 12393 31999 12396
rect 31941 12387 31999 12393
rect 32122 12384 32128 12396
rect 32180 12384 32186 12436
rect 20349 12359 20407 12365
rect 20349 12325 20361 12359
rect 20395 12356 20407 12359
rect 22002 12356 22008 12368
rect 20395 12328 22008 12356
rect 20395 12325 20407 12328
rect 20349 12319 20407 12325
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 20211 12260 20760 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 20732 12232 20760 12260
rect 20990 12248 20996 12300
rect 21048 12248 21054 12300
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20088 12152 20116 12183
rect 20530 12180 20536 12232
rect 20588 12180 20594 12232
rect 20714 12180 20720 12232
rect 20772 12180 20778 12232
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 20898 12180 20904 12232
rect 20956 12180 20962 12232
rect 21008 12220 21036 12248
rect 21836 12229 21864 12328
rect 22002 12316 22008 12328
rect 22060 12316 22066 12368
rect 22756 12356 22784 12384
rect 22388 12328 22784 12356
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21008 12192 21281 12220
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12189 21879 12223
rect 21821 12183 21879 12189
rect 22005 12223 22063 12229
rect 22005 12189 22017 12223
rect 22051 12220 22063 12223
rect 22388 12220 22416 12328
rect 22940 12297 22968 12384
rect 23201 12359 23259 12365
rect 23201 12325 23213 12359
rect 23247 12325 23259 12359
rect 23201 12319 23259 12325
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 22051 12192 22416 12220
rect 22051 12189 22063 12192
rect 22005 12183 22063 12189
rect 22830 12180 22836 12232
rect 22888 12180 22894 12232
rect 20625 12155 20683 12161
rect 20625 12152 20637 12155
rect 19306 12124 20637 12152
rect 20625 12121 20637 12124
rect 20671 12152 20683 12155
rect 20824 12152 20852 12180
rect 20671 12124 20852 12152
rect 20993 12155 21051 12161
rect 20671 12121 20683 12124
rect 20625 12115 20683 12121
rect 20993 12121 21005 12155
rect 21039 12121 21051 12155
rect 20993 12115 21051 12121
rect 21361 12155 21419 12161
rect 21361 12121 21373 12155
rect 21407 12152 21419 12155
rect 21637 12155 21695 12161
rect 21637 12152 21649 12155
rect 21407 12124 21649 12152
rect 21407 12121 21419 12124
rect 21361 12115 21419 12121
rect 21637 12121 21649 12124
rect 21683 12121 21695 12155
rect 21637 12115 21695 12121
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12053 8815 12087
rect 8757 12047 8815 12053
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10686 12084 10692 12096
rect 9916 12056 10692 12084
rect 9916 12044 9922 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 12250 12044 12256 12096
rect 12308 12084 12314 12096
rect 17862 12084 17868 12096
rect 12308 12056 17868 12084
rect 12308 12044 12314 12056
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18690 12084 18696 12096
rect 18003 12056 18696 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 19610 12044 19616 12096
rect 19668 12084 19674 12096
rect 19705 12087 19763 12093
rect 19705 12084 19717 12087
rect 19668 12056 19717 12084
rect 19668 12044 19674 12056
rect 19705 12053 19717 12056
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 21008 12084 21036 12115
rect 20864 12056 21036 12084
rect 21177 12087 21235 12093
rect 20864 12044 20870 12056
rect 21177 12053 21189 12087
rect 21223 12084 21235 12087
rect 21450 12084 21456 12096
rect 21223 12056 21456 12084
rect 21223 12053 21235 12056
rect 21177 12047 21235 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 21545 12087 21603 12093
rect 21545 12053 21557 12087
rect 21591 12084 21603 12087
rect 22940 12084 22968 12251
rect 23106 12180 23112 12232
rect 23164 12180 23170 12232
rect 23216 12220 23244 12319
rect 31754 12316 31760 12368
rect 31812 12356 31818 12368
rect 33045 12359 33103 12365
rect 31812 12328 31984 12356
rect 31812 12316 31818 12328
rect 25038 12248 25044 12300
rect 25096 12248 25102 12300
rect 25314 12248 25320 12300
rect 25372 12248 25378 12300
rect 25884 12260 26188 12288
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 23216 12192 23489 12220
rect 23477 12189 23489 12192
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23750 12180 23756 12232
rect 23808 12220 23814 12232
rect 23845 12223 23903 12229
rect 23845 12220 23857 12223
rect 23808 12192 23857 12220
rect 23808 12180 23814 12192
rect 23845 12189 23857 12192
rect 23891 12189 23903 12223
rect 23845 12183 23903 12189
rect 24949 12223 25007 12229
rect 24949 12189 24961 12223
rect 24995 12220 25007 12223
rect 25884 12220 25912 12260
rect 26160 12232 26188 12260
rect 29454 12248 29460 12300
rect 29512 12288 29518 12300
rect 31481 12291 31539 12297
rect 31481 12288 31493 12291
rect 29512 12260 31493 12288
rect 29512 12248 29518 12260
rect 24995 12192 25912 12220
rect 24995 12189 25007 12192
rect 24949 12183 25007 12189
rect 25958 12180 25964 12232
rect 26016 12180 26022 12232
rect 26142 12180 26148 12232
rect 26200 12180 26206 12232
rect 27617 12223 27675 12229
rect 27617 12189 27629 12223
rect 27663 12220 27675 12223
rect 28074 12220 28080 12232
rect 27663 12192 28080 12220
rect 27663 12189 27675 12192
rect 27617 12183 27675 12189
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12189 31263 12223
rect 31205 12183 31263 12189
rect 23124 12152 23152 12180
rect 23569 12155 23627 12161
rect 23569 12152 23581 12155
rect 23124 12124 23581 12152
rect 23569 12121 23581 12124
rect 23615 12121 23627 12155
rect 23569 12115 23627 12121
rect 23661 12155 23719 12161
rect 23661 12121 23673 12155
rect 23707 12152 23719 12155
rect 25866 12152 25872 12164
rect 23707 12124 25872 12152
rect 23707 12121 23719 12124
rect 23661 12115 23719 12121
rect 25866 12112 25872 12124
rect 25924 12112 25930 12164
rect 26053 12155 26111 12161
rect 26053 12121 26065 12155
rect 26099 12152 26111 12155
rect 27798 12152 27804 12164
rect 26099 12124 27804 12152
rect 26099 12121 26111 12124
rect 26053 12115 26111 12121
rect 27798 12112 27804 12124
rect 27856 12112 27862 12164
rect 31220 12096 31248 12183
rect 21591 12056 22968 12084
rect 21591 12053 21603 12056
rect 21545 12047 21603 12053
rect 23290 12044 23296 12096
rect 23348 12044 23354 12096
rect 25406 12044 25412 12096
rect 25464 12084 25470 12096
rect 25590 12084 25596 12096
rect 25464 12056 25596 12084
rect 25464 12044 25470 12056
rect 25590 12044 25596 12056
rect 25648 12044 25654 12096
rect 27430 12044 27436 12096
rect 27488 12044 27494 12096
rect 31202 12044 31208 12096
rect 31260 12044 31266 12096
rect 31312 12084 31340 12260
rect 31481 12257 31493 12260
rect 31527 12257 31539 12291
rect 31481 12251 31539 12257
rect 31846 12248 31852 12300
rect 31904 12248 31910 12300
rect 31389 12223 31447 12229
rect 31389 12189 31401 12223
rect 31435 12220 31447 12223
rect 31864 12220 31892 12248
rect 31435 12192 31892 12220
rect 31435 12189 31447 12192
rect 31389 12183 31447 12189
rect 31956 12152 31984 12328
rect 33045 12325 33057 12359
rect 33091 12325 33103 12359
rect 33045 12319 33103 12325
rect 32033 12223 32091 12229
rect 32033 12189 32045 12223
rect 32079 12220 32091 12223
rect 32214 12220 32220 12232
rect 32079 12192 32220 12220
rect 32079 12189 32091 12192
rect 32033 12183 32091 12189
rect 32214 12180 32220 12192
rect 32272 12180 32278 12232
rect 32309 12223 32367 12229
rect 32309 12189 32321 12223
rect 32355 12189 32367 12223
rect 33060 12220 33088 12319
rect 33873 12223 33931 12229
rect 33873 12220 33885 12223
rect 33060 12192 33885 12220
rect 32309 12183 32367 12189
rect 33873 12189 33885 12192
rect 33919 12189 33931 12223
rect 33873 12183 33931 12189
rect 32122 12152 32128 12164
rect 31956 12124 32128 12152
rect 32122 12112 32128 12124
rect 32180 12152 32186 12164
rect 32324 12152 32352 12183
rect 32180 12124 32352 12152
rect 33888 12152 33916 12183
rect 34146 12180 34152 12232
rect 34204 12180 34210 12232
rect 34514 12180 34520 12232
rect 34572 12180 34578 12232
rect 34532 12152 34560 12180
rect 33888 12124 34560 12152
rect 32180 12112 32186 12124
rect 31662 12084 31668 12096
rect 31312 12056 31668 12084
rect 31662 12044 31668 12056
rect 31720 12084 31726 12096
rect 33137 12087 33195 12093
rect 33137 12084 33149 12087
rect 31720 12056 33149 12084
rect 31720 12044 31726 12056
rect 33137 12053 33149 12056
rect 33183 12053 33195 12087
rect 33137 12047 33195 12053
rect 1104 11994 38824 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 38824 11994
rect 1104 11920 38824 11942
rect 9033 11883 9091 11889
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 9674 11880 9680 11892
rect 9079 11852 9680 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11790 11880 11796 11892
rect 11379 11852 11796 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 16298 11840 16304 11892
rect 16356 11840 16362 11892
rect 16666 11840 16672 11892
rect 16724 11840 16730 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 17083 11852 19441 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 20349 11883 20407 11889
rect 19429 11843 19487 11849
rect 19536 11852 20300 11880
rect 9232 11784 10640 11812
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 8956 11676 8984 11707
rect 9122 11676 9128 11688
rect 8956 11648 9128 11676
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 9232 11617 9260 11784
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10612 11753 10640 11784
rect 17126 11772 17132 11824
rect 17184 11772 17190 11824
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 19536 11812 19564 11852
rect 17920 11784 19564 11812
rect 17920 11772 17926 11784
rect 19702 11772 19708 11824
rect 19760 11772 19766 11824
rect 19794 11772 19800 11824
rect 19852 11772 19858 11824
rect 20272 11812 20300 11852
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 20714 11880 20720 11892
rect 20395 11852 20720 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 20898 11840 20904 11892
rect 20956 11840 20962 11892
rect 20990 11840 20996 11892
rect 21048 11889 21054 11892
rect 21048 11883 21067 11889
rect 21055 11849 21067 11883
rect 21048 11843 21067 11849
rect 21048 11840 21054 11843
rect 21174 11840 21180 11892
rect 21232 11840 21238 11892
rect 25501 11883 25559 11889
rect 25501 11849 25513 11883
rect 25547 11880 25559 11883
rect 26050 11880 26056 11892
rect 25547 11852 26056 11880
rect 25547 11849 25559 11852
rect 25501 11843 25559 11849
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 26142 11840 26148 11892
rect 26200 11880 26206 11892
rect 26237 11883 26295 11889
rect 26237 11880 26249 11883
rect 26200 11852 26249 11880
rect 26200 11840 26206 11852
rect 26237 11849 26249 11852
rect 26283 11849 26295 11883
rect 26237 11843 26295 11849
rect 26602 11840 26608 11892
rect 26660 11880 26666 11892
rect 27249 11883 27307 11889
rect 27249 11880 27261 11883
rect 26660 11852 27261 11880
rect 26660 11840 26666 11852
rect 27249 11849 27261 11852
rect 27295 11880 27307 11883
rect 27295 11852 29040 11880
rect 27295 11849 27307 11852
rect 27249 11843 27307 11849
rect 20806 11812 20812 11824
rect 20272 11784 20812 11812
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9916 11716 9965 11744
rect 9916 11704 9922 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11744 16451 11747
rect 17402 11744 17408 11756
rect 16439 11716 17408 11744
rect 16439 11713 16451 11716
rect 16393 11707 16451 11713
rect 17402 11704 17408 11716
rect 17460 11704 17466 11756
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 19978 11704 19984 11756
rect 20036 11704 20042 11756
rect 20732 11753 20760 11784
rect 20806 11772 20812 11784
rect 20864 11772 20870 11824
rect 20916 11812 20944 11840
rect 27632 11821 27660 11852
rect 25593 11815 25651 11821
rect 25593 11812 25605 11815
rect 20916 11784 25605 11812
rect 25593 11781 25605 11784
rect 25639 11781 25651 11815
rect 25593 11775 25651 11781
rect 25777 11815 25835 11821
rect 25777 11781 25789 11815
rect 25823 11812 25835 11815
rect 27617 11815 27675 11821
rect 25823 11784 27568 11812
rect 25823 11781 25835 11784
rect 25777 11775 25835 11781
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 20456 11716 20545 11744
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10318 11676 10324 11688
rect 10275 11648 10324 11676
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 17310 11636 17316 11688
rect 17368 11636 17374 11688
rect 20456 11676 20484 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 24854 11704 24860 11756
rect 24912 11744 24918 11756
rect 25225 11747 25283 11753
rect 25225 11744 25237 11747
rect 24912 11716 25237 11744
rect 24912 11704 24918 11716
rect 25225 11713 25237 11716
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 25409 11747 25467 11753
rect 25409 11713 25421 11747
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 18984 11648 20484 11676
rect 9217 11611 9275 11617
rect 9217 11608 9229 11611
rect 4120 11580 9229 11608
rect 4120 11568 4126 11580
rect 9217 11577 9229 11580
rect 9263 11577 9275 11611
rect 9217 11571 9275 11577
rect 18984 11552 19012 11648
rect 18966 11500 18972 11552
rect 19024 11500 19030 11552
rect 20364 11540 20392 11648
rect 25424 11620 25452 11707
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 26053 11747 26111 11753
rect 26053 11744 26065 11747
rect 25740 11716 26065 11744
rect 25740 11704 25746 11716
rect 26053 11713 26065 11716
rect 26099 11713 26111 11747
rect 26053 11707 26111 11713
rect 26142 11704 26148 11756
rect 26200 11744 26206 11756
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 26200 11716 27169 11744
rect 26200 11704 26206 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11713 27399 11747
rect 27540 11744 27568 11784
rect 27617 11781 27629 11815
rect 27663 11781 27675 11815
rect 27817 11815 27875 11821
rect 27817 11812 27829 11815
rect 27617 11775 27675 11781
rect 27724 11784 27829 11812
rect 27724 11744 27752 11784
rect 27817 11781 27829 11784
rect 27863 11781 27875 11815
rect 27817 11775 27875 11781
rect 29012 11753 29040 11852
rect 31662 11840 31668 11892
rect 31720 11880 31726 11892
rect 31720 11852 32260 11880
rect 31720 11840 31726 11852
rect 32122 11772 32128 11824
rect 32180 11772 32186 11824
rect 28813 11747 28871 11753
rect 28813 11744 28825 11747
rect 27540 11716 28825 11744
rect 27341 11707 27399 11713
rect 28813 11713 28825 11716
rect 28859 11713 28871 11747
rect 28813 11707 28871 11713
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11713 29055 11747
rect 28997 11707 29055 11713
rect 31481 11747 31539 11753
rect 31481 11713 31493 11747
rect 31527 11744 31539 11747
rect 31846 11744 31852 11756
rect 31527 11716 31852 11744
rect 31527 11713 31539 11716
rect 31481 11707 31539 11713
rect 25866 11636 25872 11688
rect 25924 11636 25930 11688
rect 27356 11676 27384 11707
rect 31846 11704 31852 11716
rect 31904 11704 31910 11756
rect 27356 11648 27844 11676
rect 25406 11568 25412 11620
rect 25464 11608 25470 11620
rect 26973 11611 27031 11617
rect 26973 11608 26985 11611
rect 25464 11580 26985 11608
rect 25464 11568 25470 11580
rect 26973 11577 26985 11580
rect 27019 11577 27031 11611
rect 26973 11571 27031 11577
rect 27522 11568 27528 11620
rect 27580 11568 27586 11620
rect 27816 11608 27844 11648
rect 31386 11636 31392 11688
rect 31444 11636 31450 11688
rect 31849 11611 31907 11617
rect 27816 11580 30512 11608
rect 20993 11543 21051 11549
rect 20993 11540 21005 11543
rect 20364 11512 21005 11540
rect 20993 11509 21005 11512
rect 21039 11540 21051 11543
rect 21450 11540 21456 11552
rect 21039 11512 21456 11540
rect 21039 11509 21051 11512
rect 20993 11503 21051 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 27816 11549 27844 11580
rect 30484 11552 30512 11580
rect 31849 11577 31861 11611
rect 31895 11608 31907 11611
rect 31938 11608 31944 11620
rect 31895 11580 31944 11608
rect 31895 11577 31907 11580
rect 31849 11571 31907 11577
rect 31938 11568 31944 11580
rect 31996 11568 32002 11620
rect 32232 11608 32260 11852
rect 32582 11840 32588 11892
rect 32640 11840 32646 11892
rect 32401 11611 32459 11617
rect 32401 11608 32413 11611
rect 32232 11580 32413 11608
rect 32401 11577 32413 11580
rect 32447 11577 32459 11611
rect 32401 11571 32459 11577
rect 27801 11543 27859 11549
rect 27801 11509 27813 11543
rect 27847 11509 27859 11543
rect 27801 11503 27859 11509
rect 27985 11543 28043 11549
rect 27985 11509 27997 11543
rect 28031 11540 28043 11543
rect 28258 11540 28264 11552
rect 28031 11512 28264 11540
rect 28031 11509 28043 11512
rect 27985 11503 28043 11509
rect 28258 11500 28264 11512
rect 28316 11540 28322 11552
rect 28626 11540 28632 11552
rect 28316 11512 28632 11540
rect 28316 11500 28322 11512
rect 28626 11500 28632 11512
rect 28684 11500 28690 11552
rect 28902 11500 28908 11552
rect 28960 11500 28966 11552
rect 30466 11500 30472 11552
rect 30524 11500 30530 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 15933 11339 15991 11345
rect 15933 11305 15945 11339
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 12069 11271 12127 11277
rect 12069 11237 12081 11271
rect 12115 11268 12127 11271
rect 12342 11268 12348 11280
rect 12115 11240 12348 11268
rect 12115 11237 12127 11240
rect 12069 11231 12127 11237
rect 12342 11228 12348 11240
rect 12400 11268 12406 11280
rect 15948 11268 15976 11299
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 23290 11336 23296 11348
rect 22664 11308 23296 11336
rect 12400 11240 15240 11268
rect 15948 11240 16160 11268
rect 12400 11228 12406 11240
rect 14292 11209 14320 11240
rect 13633 11203 13691 11209
rect 11900 11172 12664 11200
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 11333 11135 11391 11141
rect 11333 11132 11345 11135
rect 10744 11104 11345 11132
rect 10744 11092 10750 11104
rect 11333 11101 11345 11104
rect 11379 11132 11391 11135
rect 11609 11135 11667 11141
rect 11609 11132 11621 11135
rect 11379 11104 11621 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11609 11101 11621 11104
rect 11655 11101 11667 11135
rect 11609 11095 11667 11101
rect 11698 11092 11704 11144
rect 11756 11092 11762 11144
rect 11900 11141 11928 11172
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 12032 11104 12173 11132
rect 12032 11092 12038 11104
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12434 11092 12440 11144
rect 12492 11092 12498 11144
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 10778 11064 10784 11076
rect 9180 11036 10784 11064
rect 9180 11024 9186 11036
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 12636 11073 12664 11172
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13679 11172 14105 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14366 11160 14372 11212
rect 14424 11200 14430 11212
rect 14826 11200 14832 11212
rect 14424 11172 14832 11200
rect 14424 11160 14430 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 15212 11141 15240 11240
rect 16132 11212 16160 11240
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 17402 11160 17408 11212
rect 17460 11200 17466 11212
rect 17460 11172 17816 11200
rect 17460 11160 17466 11172
rect 15013 11135 15071 11141
rect 15013 11134 15025 11135
rect 14936 11132 15025 11134
rect 13596 11106 15025 11132
rect 13596 11104 14964 11106
rect 13596 11092 13602 11104
rect 15013 11101 15025 11106
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11132 15255 11135
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 15243 11104 15485 11132
rect 15243 11101 15255 11104
rect 15197 11095 15255 11101
rect 15473 11101 15485 11104
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 11425 11067 11483 11073
rect 11425 11033 11437 11067
rect 11471 11064 11483 11067
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 11471 11036 12265 11064
rect 11471 11033 11483 11036
rect 11425 11027 11483 11033
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 12621 11067 12679 11073
rect 12621 11033 12633 11067
rect 12667 11064 12679 11067
rect 12667 11036 14320 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 14292 11008 14320 11036
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 13998 10996 14004 11008
rect 13955 10968 14004 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 14332 10968 14749 10996
rect 14332 10956 14338 10968
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 14737 10959 14795 10965
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 15120 10996 15148 11095
rect 15562 11092 15568 11144
rect 15620 11132 15626 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15620 11104 15761 11132
rect 15620 11092 15626 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 15948 11064 15976 11095
rect 17218 11092 17224 11144
rect 17276 11132 17282 11144
rect 17788 11141 17816 11172
rect 17972 11172 18460 11200
rect 17972 11141 18000 11172
rect 18432 11144 18460 11172
rect 17681 11135 17739 11141
rect 17681 11132 17693 11135
rect 17276 11104 17693 11132
rect 17276 11092 17282 11104
rect 17681 11101 17693 11104
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 17862 11064 17868 11076
rect 15948 11036 17868 11064
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 18064 11064 18092 11095
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 22664 11141 22692 11308
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23382 11296 23388 11348
rect 23440 11336 23446 11348
rect 24302 11336 24308 11348
rect 23440 11308 24308 11336
rect 23440 11296 23446 11308
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 24394 11296 24400 11348
rect 24452 11296 24458 11348
rect 25682 11336 25688 11348
rect 24780 11308 25688 11336
rect 23661 11271 23719 11277
rect 23661 11268 23673 11271
rect 23492 11240 23673 11268
rect 22925 11203 22983 11209
rect 22925 11169 22937 11203
rect 22971 11200 22983 11203
rect 23382 11200 23388 11212
rect 22971 11172 23388 11200
rect 22971 11169 22983 11172
rect 22925 11163 22983 11169
rect 23382 11160 23388 11172
rect 23440 11160 23446 11212
rect 22649 11135 22707 11141
rect 22649 11101 22661 11135
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 18064 11036 18552 11064
rect 18524 11008 18552 11036
rect 22830 11024 22836 11076
rect 22888 11064 22894 11076
rect 23382 11064 23388 11076
rect 22888 11036 23388 11064
rect 22888 11024 22894 11036
rect 23382 11024 23388 11036
rect 23440 11024 23446 11076
rect 14884 10968 15148 10996
rect 14884 10956 14890 10968
rect 15378 10956 15384 11008
rect 15436 10956 15442 11008
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 18233 10999 18291 11005
rect 18233 10996 18245 10999
rect 18104 10968 18245 10996
rect 18104 10956 18110 10968
rect 18233 10965 18245 10968
rect 18279 10965 18291 10999
rect 18233 10959 18291 10965
rect 18506 10956 18512 11008
rect 18564 10956 18570 11008
rect 22278 10956 22284 11008
rect 22336 10956 22342 11008
rect 22738 10956 22744 11008
rect 22796 10996 22802 11008
rect 23492 10996 23520 11240
rect 23661 11237 23673 11240
rect 23707 11237 23719 11271
rect 23661 11231 23719 11237
rect 24780 11212 24808 11308
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 25866 11296 25872 11348
rect 25924 11296 25930 11348
rect 28718 11296 28724 11348
rect 28776 11296 28782 11348
rect 28902 11296 28908 11348
rect 28960 11296 28966 11348
rect 32214 11296 32220 11348
rect 32272 11336 32278 11348
rect 38194 11336 38200 11348
rect 32272 11308 38200 11336
rect 32272 11296 32278 11308
rect 38194 11296 38200 11308
rect 38252 11296 38258 11348
rect 25884 11268 25912 11296
rect 25148 11240 25912 11268
rect 26988 11240 28304 11268
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 23891 11172 24440 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24412 11141 24440 11172
rect 24762 11160 24768 11212
rect 24820 11160 24826 11212
rect 25148 11209 25176 11240
rect 26988 11212 27016 11240
rect 25133 11203 25191 11209
rect 25133 11169 25145 11203
rect 25179 11169 25191 11203
rect 25133 11163 25191 11169
rect 25222 11160 25228 11212
rect 25280 11160 25286 11212
rect 25409 11203 25467 11209
rect 25409 11169 25421 11203
rect 25455 11200 25467 11203
rect 26970 11200 26976 11212
rect 25455 11172 26976 11200
rect 25455 11169 25467 11172
rect 25409 11163 25467 11169
rect 26970 11160 26976 11172
rect 27028 11160 27034 11212
rect 28276 11209 28304 11240
rect 27801 11203 27859 11209
rect 27801 11169 27813 11203
rect 27847 11200 27859 11203
rect 28261 11203 28319 11209
rect 27847 11172 28028 11200
rect 27847 11169 27859 11172
rect 27801 11163 27859 11169
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24670 11132 24676 11144
rect 24627 11104 24676 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 24670 11092 24676 11104
rect 24728 11132 24734 11144
rect 28000 11141 28028 11172
rect 28261 11169 28273 11203
rect 28307 11169 28319 11203
rect 28920 11200 28948 11296
rect 28920 11172 29408 11200
rect 28261 11163 28319 11169
rect 25685 11135 25743 11141
rect 25685 11132 25697 11135
rect 24728 11104 25697 11132
rect 24728 11092 24734 11104
rect 25685 11101 25697 11104
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 27893 11135 27951 11141
rect 27893 11101 27905 11135
rect 27939 11101 27951 11135
rect 27893 11095 27951 11101
rect 27985 11135 28043 11141
rect 27985 11101 27997 11135
rect 28031 11101 28043 11135
rect 27985 11095 28043 11101
rect 25222 11024 25228 11076
rect 25280 11064 25286 11076
rect 25501 11067 25559 11073
rect 25501 11064 25513 11067
rect 25280 11036 25513 11064
rect 25280 11024 25286 11036
rect 25501 11033 25513 11036
rect 25547 11033 25559 11067
rect 27908 11064 27936 11095
rect 28166 11092 28172 11144
rect 28224 11092 28230 11144
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 28276 11104 28365 11132
rect 28074 11064 28080 11076
rect 27908 11036 28080 11064
rect 25501 11027 25559 11033
rect 28074 11024 28080 11036
rect 28132 11024 28138 11076
rect 28276 11008 28304 11104
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28552 11064 28580 11095
rect 28626 11092 28632 11144
rect 28684 11132 28690 11144
rect 29380 11141 29408 11172
rect 29089 11135 29147 11141
rect 29089 11132 29101 11135
rect 28684 11104 29101 11132
rect 28684 11092 28690 11104
rect 29089 11101 29101 11104
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 29365 11135 29423 11141
rect 29365 11101 29377 11135
rect 29411 11101 29423 11135
rect 29365 11095 29423 11101
rect 30466 11092 30472 11144
rect 30524 11092 30530 11144
rect 30484 11064 30512 11092
rect 32122 11064 32128 11076
rect 28552 11036 28856 11064
rect 30484 11036 32128 11064
rect 22796 10968 23520 10996
rect 22796 10956 22802 10968
rect 28258 10956 28264 11008
rect 28316 10956 28322 11008
rect 28350 10956 28356 11008
rect 28408 10996 28414 11008
rect 28552 10996 28580 11036
rect 28828 11008 28856 11036
rect 32122 11024 32128 11036
rect 32180 11024 32186 11076
rect 28408 10968 28580 10996
rect 28408 10956 28414 10968
rect 28810 10956 28816 11008
rect 28868 10956 28874 11008
rect 28902 10956 28908 11008
rect 28960 10956 28966 11008
rect 29273 10999 29331 11005
rect 29273 10965 29285 10999
rect 29319 10996 29331 10999
rect 30377 10999 30435 11005
rect 30377 10996 30389 10999
rect 29319 10968 30389 10996
rect 29319 10965 29331 10968
rect 29273 10959 29331 10965
rect 30377 10965 30389 10968
rect 30423 10996 30435 10999
rect 30926 10996 30932 11008
rect 30423 10968 30932 10996
rect 30423 10965 30435 10968
rect 30377 10959 30435 10965
rect 30926 10956 30932 10968
rect 30984 10956 30990 11008
rect 1104 10906 38824 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 38824 10906
rect 1104 10832 38824 10854
rect 11698 10752 11704 10804
rect 11756 10752 11762 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 14415 10764 15332 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 12434 10724 12440 10736
rect 11624 10696 12440 10724
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10502 10656 10508 10668
rect 10183 10628 10508 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10060 10520 10088 10619
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 11624 10665 11652 10696
rect 12434 10684 12440 10696
rect 12492 10684 12498 10736
rect 14108 10696 14688 10724
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10704 10588 10732 10619
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 14108 10665 14136 10696
rect 14660 10668 14688 10696
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 14093 10659 14151 10665
rect 12299 10628 14044 10656
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 10778 10588 10784 10600
rect 10704 10560 10784 10588
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 12342 10548 12348 10600
rect 12400 10548 12406 10600
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10557 13783 10591
rect 14016 10588 14044 10628
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14274 10656 14280 10668
rect 14231 10628 14280 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14366 10616 14372 10668
rect 14424 10616 14430 10668
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 14384 10588 14412 10616
rect 14016 10560 14412 10588
rect 13725 10551 13783 10557
rect 12526 10520 12532 10532
rect 10060 10492 12532 10520
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9766 10452 9772 10464
rect 9723 10424 9772 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 12618 10412 12624 10464
rect 12676 10412 12682 10464
rect 13556 10452 13584 10548
rect 13740 10520 13768 10551
rect 13906 10520 13912 10532
rect 13740 10492 13912 10520
rect 13906 10480 13912 10492
rect 13964 10520 13970 10532
rect 14476 10520 14504 10619
rect 14642 10616 14648 10668
rect 14700 10616 14706 10668
rect 15304 10588 15332 10764
rect 15378 10752 15384 10804
rect 15436 10792 15442 10804
rect 16041 10795 16099 10801
rect 16041 10792 16053 10795
rect 15436 10764 16053 10792
rect 15436 10752 15442 10764
rect 16041 10761 16053 10764
rect 16087 10761 16099 10795
rect 16041 10755 16099 10761
rect 16209 10795 16267 10801
rect 16209 10761 16221 10795
rect 16255 10761 16267 10795
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 16209 10755 16267 10761
rect 17512 10764 18245 10792
rect 15396 10656 15424 10752
rect 15841 10727 15899 10733
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 15887 10696 15921 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15396 10628 15485 10656
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15749 10659 15807 10665
rect 15611 10628 15700 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15672 10588 15700 10628
rect 15749 10625 15761 10659
rect 15795 10656 15807 10659
rect 15856 10656 15884 10687
rect 16114 10656 16120 10668
rect 15795 10628 16120 10656
rect 15795 10625 15807 10628
rect 15749 10619 15807 10625
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16224 10656 16252 10755
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16224 10628 16313 10656
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10656 16543 10659
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16531 10628 16957 10656
rect 16531 10625 16543 10628
rect 16485 10619 16543 10625
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 16500 10588 16528 10619
rect 17218 10616 17224 10668
rect 17276 10616 17282 10668
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 17512 10665 17540 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24670 10792 24676 10804
rect 24075 10764 24676 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 24762 10752 24768 10804
rect 24820 10752 24826 10804
rect 27430 10752 27436 10804
rect 27488 10752 27494 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 28353 10795 28411 10801
rect 28353 10792 28365 10795
rect 28224 10764 28365 10792
rect 28224 10752 28230 10764
rect 28353 10761 28365 10764
rect 28399 10761 28411 10795
rect 28902 10792 28908 10804
rect 28353 10755 28411 10761
rect 28618 10764 28908 10792
rect 18046 10724 18052 10736
rect 17696 10696 18052 10724
rect 17696 10665 17724 10696
rect 18046 10684 18052 10696
rect 18104 10684 18110 10736
rect 18340 10696 19012 10724
rect 17497 10659 17555 10665
rect 17497 10625 17509 10659
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 17957 10659 18015 10665
rect 17957 10656 17969 10659
rect 17920 10628 17969 10656
rect 17920 10616 17926 10628
rect 17957 10625 17969 10628
rect 18003 10656 18015 10659
rect 18340 10656 18368 10696
rect 18003 10628 18368 10656
rect 18003 10625 18015 10628
rect 17957 10619 18015 10625
rect 18414 10616 18420 10668
rect 18472 10616 18478 10668
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 18984 10665 19012 10696
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18564 10628 18613 10656
rect 18564 10616 18570 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 18969 10659 19027 10665
rect 18969 10625 18981 10659
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22278 10656 22284 10668
rect 22051 10628 22284 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 24688 10665 24716 10752
rect 26050 10724 26056 10736
rect 25976 10696 26056 10724
rect 24673 10659 24731 10665
rect 24673 10625 24685 10659
rect 24719 10625 24731 10659
rect 24673 10619 24731 10625
rect 24857 10659 24915 10665
rect 24857 10625 24869 10659
rect 24903 10656 24915 10659
rect 25222 10656 25228 10668
rect 24903 10628 25228 10656
rect 24903 10625 24915 10628
rect 24857 10619 24915 10625
rect 25222 10616 25228 10628
rect 25280 10616 25286 10668
rect 25406 10616 25412 10668
rect 25464 10616 25470 10668
rect 25498 10616 25504 10668
rect 25556 10616 25562 10668
rect 25976 10665 26004 10696
rect 26050 10684 26056 10696
rect 26108 10684 26114 10736
rect 26970 10684 26976 10736
rect 27028 10684 27034 10736
rect 27065 10727 27123 10733
rect 27065 10693 27077 10727
rect 27111 10724 27123 10727
rect 27448 10724 27476 10752
rect 28618 10733 28646 10764
rect 28902 10752 28908 10764
rect 28960 10752 28966 10804
rect 29917 10795 29975 10801
rect 29917 10792 29929 10795
rect 29748 10764 29929 10792
rect 27111 10696 27476 10724
rect 27111 10693 27123 10696
rect 27065 10687 27123 10693
rect 25777 10659 25835 10665
rect 25777 10656 25789 10659
rect 25700 10628 25789 10656
rect 15304 10560 15700 10588
rect 13964 10492 14504 10520
rect 13964 10480 13970 10492
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 13556 10424 14565 10452
rect 14553 10421 14565 10424
rect 14599 10452 14611 10455
rect 15562 10452 15568 10464
rect 14599 10424 15568 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 15672 10452 15700 10560
rect 15764 10560 16528 10588
rect 16761 10591 16819 10597
rect 15764 10529 15792 10560
rect 16761 10557 16773 10591
rect 16807 10588 16819 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 16807 10560 18889 10588
rect 16807 10557 16819 10560
rect 16761 10551 16819 10557
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 22738 10548 22744 10600
rect 22796 10588 22802 10600
rect 23569 10591 23627 10597
rect 23569 10588 23581 10591
rect 22796 10560 23581 10588
rect 22796 10548 22802 10560
rect 23569 10557 23581 10560
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 15749 10523 15807 10529
rect 15749 10489 15761 10523
rect 15795 10489 15807 10523
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 15749 10483 15807 10489
rect 16040 10492 17785 10520
rect 16040 10461 16068 10492
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 17773 10483 17831 10489
rect 17862 10480 17868 10532
rect 17920 10480 17926 10532
rect 18141 10523 18199 10529
rect 18141 10489 18153 10523
rect 18187 10520 18199 10523
rect 18782 10520 18788 10532
rect 18187 10492 18788 10520
rect 18187 10489 18199 10492
rect 18141 10483 18199 10489
rect 18782 10480 18788 10492
rect 18840 10480 18846 10532
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 23937 10523 23995 10529
rect 23937 10520 23949 10523
rect 23440 10492 23949 10520
rect 23440 10480 23446 10492
rect 23937 10489 23949 10492
rect 23983 10520 23995 10523
rect 24026 10520 24032 10532
rect 23983 10492 24032 10520
rect 23983 10489 23995 10492
rect 23937 10483 23995 10489
rect 24026 10480 24032 10492
rect 24084 10520 24090 10532
rect 25424 10520 25452 10616
rect 24084 10492 25452 10520
rect 24084 10480 24090 10492
rect 16025 10455 16083 10461
rect 16025 10452 16037 10455
rect 15672 10424 16037 10452
rect 16025 10421 16037 10424
rect 16071 10421 16083 10455
rect 16025 10415 16083 10421
rect 16298 10412 16304 10464
rect 16356 10412 16362 10464
rect 19337 10455 19395 10461
rect 19337 10421 19349 10455
rect 19383 10452 19395 10455
rect 19886 10452 19892 10464
rect 19383 10424 19892 10452
rect 19383 10421 19395 10424
rect 19337 10415 19395 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 21692 10424 21833 10452
rect 21692 10412 21698 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 25406 10412 25412 10464
rect 25464 10452 25470 10464
rect 25700 10461 25728 10628
rect 25777 10625 25789 10628
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 25961 10659 26019 10665
rect 25961 10625 25973 10659
rect 26007 10625 26019 10659
rect 26988 10656 27016 10684
rect 27448 10665 27476 10696
rect 28603 10727 28661 10733
rect 28603 10693 28615 10727
rect 28649 10693 28661 10727
rect 28603 10687 28661 10693
rect 28813 10727 28871 10733
rect 28813 10693 28825 10727
rect 28859 10724 28871 10727
rect 29181 10727 29239 10733
rect 29181 10724 29193 10727
rect 28859 10696 29193 10724
rect 28859 10693 28871 10696
rect 28813 10687 28871 10693
rect 29181 10693 29193 10696
rect 29227 10693 29239 10727
rect 29181 10687 29239 10693
rect 29748 10668 29776 10764
rect 29917 10761 29929 10764
rect 29963 10761 29975 10795
rect 31297 10795 31355 10801
rect 31297 10792 31309 10795
rect 29917 10755 29975 10761
rect 30852 10764 31309 10792
rect 30852 10733 30880 10764
rect 31297 10761 31309 10764
rect 31343 10792 31355 10795
rect 31386 10792 31392 10804
rect 31343 10764 31392 10792
rect 31343 10761 31355 10764
rect 31297 10755 31355 10761
rect 31386 10752 31392 10764
rect 31444 10752 31450 10804
rect 32122 10752 32128 10804
rect 32180 10752 32186 10804
rect 30621 10727 30679 10733
rect 30621 10724 30633 10727
rect 29840 10696 30633 10724
rect 27249 10659 27307 10665
rect 27249 10656 27261 10659
rect 26988 10628 27261 10656
rect 25961 10619 26019 10625
rect 27249 10625 27261 10628
rect 27295 10625 27307 10659
rect 27249 10619 27307 10625
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10625 27399 10659
rect 27341 10619 27399 10625
rect 27433 10659 27491 10665
rect 27433 10625 27445 10659
rect 27479 10625 27491 10659
rect 27433 10619 27491 10625
rect 27264 10520 27292 10619
rect 27356 10588 27384 10619
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 27709 10659 27767 10665
rect 27709 10625 27721 10659
rect 27755 10656 27767 10659
rect 27982 10656 27988 10668
rect 27755 10628 27988 10656
rect 27755 10625 27767 10628
rect 27709 10619 27767 10625
rect 27724 10588 27752 10619
rect 27982 10616 27988 10628
rect 28040 10616 28046 10668
rect 28169 10659 28227 10665
rect 28169 10625 28181 10659
rect 28215 10656 28227 10659
rect 28350 10656 28356 10668
rect 28215 10628 28356 10656
rect 28215 10625 28227 10628
rect 28169 10619 28227 10625
rect 28350 10616 28356 10628
rect 28408 10616 28414 10668
rect 28442 10616 28448 10668
rect 28500 10616 28506 10668
rect 28718 10616 28724 10668
rect 28776 10616 28782 10668
rect 28902 10616 28908 10668
rect 28960 10616 28966 10668
rect 29365 10659 29423 10665
rect 29365 10656 29377 10659
rect 29012 10628 29377 10656
rect 27356 10560 27752 10588
rect 27522 10520 27528 10532
rect 27264 10492 27528 10520
rect 27522 10480 27528 10492
rect 27580 10480 27586 10532
rect 29012 10520 29040 10628
rect 29365 10625 29377 10628
rect 29411 10625 29423 10659
rect 29365 10619 29423 10625
rect 29457 10659 29515 10665
rect 29457 10625 29469 10659
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10625 29699 10659
rect 29641 10619 29699 10625
rect 29472 10588 29500 10619
rect 27908 10492 29040 10520
rect 29196 10560 29500 10588
rect 27908 10464 27936 10492
rect 29196 10464 29224 10560
rect 29656 10464 29684 10619
rect 29730 10616 29736 10668
rect 29788 10616 29794 10668
rect 29840 10600 29868 10696
rect 30621 10693 30633 10696
rect 30667 10693 30679 10727
rect 30621 10687 30679 10693
rect 30837 10727 30895 10733
rect 30837 10693 30849 10727
rect 30883 10693 30895 10727
rect 30837 10687 30895 10693
rect 30193 10659 30251 10665
rect 30193 10625 30205 10659
rect 30239 10656 30251 10659
rect 30852 10656 30880 10687
rect 30926 10684 30932 10736
rect 30984 10684 30990 10736
rect 30239 10628 30880 10656
rect 31113 10659 31171 10665
rect 30239 10625 30251 10628
rect 30193 10619 30251 10625
rect 31113 10625 31125 10659
rect 31159 10656 31171 10659
rect 31294 10656 31300 10668
rect 31159 10628 31300 10656
rect 31159 10625 31171 10628
rect 31113 10619 31171 10625
rect 31294 10616 31300 10628
rect 31352 10616 31358 10668
rect 32858 10616 32864 10668
rect 32916 10656 32922 10668
rect 35342 10656 35348 10668
rect 32916 10628 35348 10656
rect 32916 10616 32922 10628
rect 35342 10616 35348 10628
rect 35400 10616 35406 10668
rect 29822 10548 29828 10600
rect 29880 10548 29886 10600
rect 30374 10548 30380 10600
rect 30432 10588 30438 10600
rect 33137 10591 33195 10597
rect 30432 10560 30696 10588
rect 30432 10548 30438 10560
rect 25685 10455 25743 10461
rect 25685 10452 25697 10455
rect 25464 10424 25697 10452
rect 25464 10412 25470 10424
rect 25685 10421 25697 10424
rect 25731 10421 25743 10455
rect 25685 10415 25743 10421
rect 25866 10412 25872 10464
rect 25924 10412 25930 10464
rect 27338 10412 27344 10464
rect 27396 10412 27402 10464
rect 27890 10412 27896 10464
rect 27948 10412 27954 10464
rect 28074 10412 28080 10464
rect 28132 10412 28138 10464
rect 29086 10412 29092 10464
rect 29144 10412 29150 10464
rect 29178 10412 29184 10464
rect 29236 10412 29242 10464
rect 29638 10412 29644 10464
rect 29696 10452 29702 10464
rect 30668 10461 30696 10560
rect 33137 10557 33149 10591
rect 33183 10588 33195 10591
rect 34146 10588 34152 10600
rect 33183 10560 34152 10588
rect 33183 10557 33195 10560
rect 33137 10551 33195 10557
rect 30469 10455 30527 10461
rect 30469 10452 30481 10455
rect 29696 10424 30481 10452
rect 29696 10412 29702 10424
rect 30469 10421 30481 10424
rect 30515 10421 30527 10455
rect 30469 10415 30527 10421
rect 30653 10455 30711 10461
rect 30653 10421 30665 10455
rect 30699 10421 30711 10455
rect 30653 10415 30711 10421
rect 30834 10412 30840 10464
rect 30892 10452 30898 10464
rect 33152 10452 33180 10551
rect 34146 10548 34152 10560
rect 34204 10548 34210 10600
rect 30892 10424 33180 10452
rect 30892 10412 30898 10424
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10560 10220 10701 10248
rect 10560 10208 10566 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 12434 10248 12440 10260
rect 10689 10211 10747 10217
rect 11348 10220 12440 10248
rect 8938 10072 8944 10124
rect 8996 10072 9002 10124
rect 10594 10044 10600 10056
rect 10350 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 10704 10044 10732 10211
rect 11348 10189 11376 10220
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12526 10208 12532 10260
rect 12584 10208 12590 10260
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 13817 10251 13875 10257
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 13906 10248 13912 10260
rect 13863 10220 13912 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14461 10251 14519 10257
rect 14461 10217 14473 10251
rect 14507 10248 14519 10251
rect 14642 10248 14648 10260
rect 14507 10220 14648 10248
rect 14507 10217 14519 10220
rect 14461 10211 14519 10217
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16448 10220 17049 10248
rect 16448 10208 16454 10220
rect 17037 10217 17049 10220
rect 17083 10248 17095 10251
rect 17862 10248 17868 10260
rect 17083 10220 17868 10248
rect 17083 10217 17095 10220
rect 17037 10211 17095 10217
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 21266 10248 21272 10260
rect 20947 10220 21272 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 21440 10251 21498 10257
rect 21440 10217 21452 10251
rect 21486 10248 21498 10251
rect 21634 10248 21640 10260
rect 21486 10220 21640 10248
rect 21486 10217 21498 10220
rect 21440 10211 21498 10217
rect 21634 10208 21640 10220
rect 21692 10208 21698 10260
rect 22738 10208 22744 10260
rect 22796 10248 22802 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 22796 10220 22937 10248
rect 22796 10208 22802 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 11333 10183 11391 10189
rect 11333 10149 11345 10183
rect 11379 10149 11391 10183
rect 11333 10143 11391 10149
rect 11701 10183 11759 10189
rect 11701 10149 11713 10183
rect 11747 10149 11759 10183
rect 11701 10143 11759 10149
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11514 10112 11520 10124
rect 11103 10084 11520 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11514 10072 11520 10084
rect 11572 10112 11578 10124
rect 11716 10112 11744 10143
rect 11572 10084 11744 10112
rect 12636 10112 12664 10208
rect 13188 10152 17632 10180
rect 12636 10084 12940 10112
rect 11572 10072 11578 10084
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10704 10016 10977 10044
rect 10965 10013 10977 10016
rect 11011 10044 11023 10047
rect 11425 10047 11483 10053
rect 11425 10044 11437 10047
rect 11011 10016 11437 10044
rect 11011 10013 11023 10016
rect 10965 10007 11023 10013
rect 11425 10013 11437 10016
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 12912 10053 12940 10084
rect 13188 10056 13216 10152
rect 13648 10084 14964 10112
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13170 10044 13176 10056
rect 13127 10016 13176 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 9214 9936 9220 9988
rect 9272 9936 9278 9988
rect 12820 9976 12848 10004
rect 13648 9976 13676 10084
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10044 13967 10047
rect 13955 10016 14320 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 12820 9948 13676 9976
rect 13740 9976 13768 10007
rect 14292 9988 14320 10016
rect 14093 9979 14151 9985
rect 14093 9976 14105 9979
rect 13740 9948 14105 9976
rect 11885 9911 11943 9917
rect 11885 9877 11897 9911
rect 11931 9908 11943 9911
rect 13740 9908 13768 9948
rect 14093 9945 14105 9948
rect 14139 9945 14151 9979
rect 14093 9939 14151 9945
rect 14274 9936 14280 9988
rect 14332 9936 14338 9988
rect 14936 9976 14964 10084
rect 16224 10053 16252 10152
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17218 10112 17224 10124
rect 16908 10084 17224 10112
rect 16908 10072 16914 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 16393 10047 16451 10053
rect 16393 10044 16405 10047
rect 16356 10016 16405 10044
rect 16356 10004 16362 10016
rect 16393 10013 16405 10016
rect 16439 10013 16451 10047
rect 16393 10007 16451 10013
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16942 10044 16948 10056
rect 16623 10016 16948 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10044 17371 10047
rect 17494 10044 17500 10056
rect 17359 10016 17500 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 16485 9979 16543 9985
rect 16485 9976 16497 9979
rect 14936 9948 16497 9976
rect 16485 9945 16497 9948
rect 16531 9945 16543 9979
rect 17604 9976 17632 10152
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 17828 10152 18797 10180
rect 17828 10140 17834 10152
rect 18785 10149 18797 10152
rect 18831 10149 18843 10183
rect 18785 10143 18843 10149
rect 20073 10183 20131 10189
rect 20073 10149 20085 10183
rect 20119 10149 20131 10183
rect 20073 10143 20131 10149
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 18012 10084 18337 10112
rect 18012 10072 18018 10084
rect 18325 10081 18337 10084
rect 18371 10112 18383 10115
rect 18506 10112 18512 10124
rect 18371 10084 18512 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 18414 10004 18420 10056
rect 18472 10044 18478 10056
rect 20088 10044 20116 10143
rect 20349 10115 20407 10121
rect 20349 10081 20361 10115
rect 20395 10081 20407 10115
rect 21177 10115 21235 10121
rect 20349 10075 20407 10081
rect 20456 10084 21128 10112
rect 18472 10016 20116 10044
rect 18472 10004 18478 10016
rect 19978 9976 19984 9988
rect 17604 9948 19984 9976
rect 16485 9939 16543 9945
rect 19978 9936 19984 9948
rect 20036 9936 20042 9988
rect 20364 9976 20392 10075
rect 20456 10053 20484 10084
rect 21100 10056 21128 10084
rect 21177 10081 21189 10115
rect 21223 10112 21235 10115
rect 21818 10112 21824 10124
rect 21223 10084 21824 10112
rect 21223 10081 21235 10084
rect 21177 10075 21235 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10013 20499 10047
rect 20990 10044 20996 10056
rect 20441 10007 20499 10013
rect 20640 10016 20996 10044
rect 20640 9976 20668 10016
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 21082 10004 21088 10056
rect 21140 10004 21146 10056
rect 22940 10044 22968 10211
rect 28074 10208 28080 10260
rect 28132 10208 28138 10260
rect 28902 10208 28908 10260
rect 28960 10208 28966 10260
rect 30285 10251 30343 10257
rect 30285 10217 30297 10251
rect 30331 10248 30343 10251
rect 30374 10248 30380 10260
rect 30331 10220 30380 10248
rect 30331 10217 30343 10220
rect 30285 10211 30343 10217
rect 30374 10208 30380 10220
rect 30432 10208 30438 10260
rect 30926 10208 30932 10260
rect 30984 10208 30990 10260
rect 31849 10251 31907 10257
rect 31849 10217 31861 10251
rect 31895 10248 31907 10251
rect 32858 10248 32864 10260
rect 31895 10220 32864 10248
rect 31895 10217 31907 10220
rect 31849 10211 31907 10217
rect 32858 10208 32864 10220
rect 32916 10208 32922 10260
rect 28092 10180 28120 10208
rect 29181 10183 29239 10189
rect 29181 10180 29193 10183
rect 25702 10152 26924 10180
rect 28092 10152 29193 10180
rect 23753 10047 23811 10053
rect 23753 10044 23765 10047
rect 22940 10016 23765 10044
rect 23753 10013 23765 10016
rect 23799 10013 23811 10047
rect 24029 10047 24087 10053
rect 24029 10044 24041 10047
rect 23753 10007 23811 10013
rect 23952 10016 24041 10044
rect 23952 9988 23980 10016
rect 24029 10013 24041 10016
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 25314 10004 25320 10056
rect 25372 10004 25378 10056
rect 25702 10053 25730 10152
rect 25866 10072 25872 10124
rect 25924 10112 25930 10124
rect 26896 10121 26924 10152
rect 29181 10149 29193 10152
rect 29227 10180 29239 10183
rect 29730 10180 29736 10192
rect 29227 10152 29736 10180
rect 29227 10149 29239 10152
rect 29181 10143 29239 10149
rect 29730 10140 29736 10152
rect 29788 10140 29794 10192
rect 30944 10180 30972 10208
rect 30208 10152 30972 10180
rect 26237 10115 26295 10121
rect 26237 10112 26249 10115
rect 25924 10084 26249 10112
rect 25924 10072 25930 10084
rect 25685 10047 25743 10053
rect 25685 10013 25697 10047
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 25774 10004 25780 10056
rect 25832 10004 25838 10056
rect 25976 10053 26004 10084
rect 26237 10081 26249 10084
rect 26283 10081 26295 10115
rect 26237 10075 26295 10081
rect 26697 10115 26755 10121
rect 26697 10081 26709 10115
rect 26743 10081 26755 10115
rect 26697 10075 26755 10081
rect 26881 10115 26939 10121
rect 26881 10081 26893 10115
rect 26927 10112 26939 10115
rect 28442 10112 28448 10124
rect 26927 10084 28448 10112
rect 26927 10081 26939 10084
rect 26881 10075 26939 10081
rect 25961 10047 26019 10053
rect 25961 10013 25973 10047
rect 26007 10013 26019 10047
rect 25961 10007 26019 10013
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10044 26387 10047
rect 26602 10044 26608 10056
rect 26375 10016 26608 10044
rect 26375 10013 26387 10016
rect 26329 10007 26387 10013
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 20364 9948 20668 9976
rect 22186 9936 22192 9988
rect 22244 9936 22250 9988
rect 23934 9936 23940 9988
rect 23992 9936 23998 9988
rect 25409 9979 25467 9985
rect 25409 9945 25421 9979
rect 25455 9945 25467 9979
rect 25409 9939 25467 9945
rect 25501 9979 25559 9985
rect 25501 9945 25513 9979
rect 25547 9976 25559 9979
rect 25869 9979 25927 9985
rect 25869 9976 25881 9979
rect 25547 9948 25881 9976
rect 25547 9945 25559 9948
rect 25501 9939 25559 9945
rect 25869 9945 25881 9948
rect 25915 9945 25927 9979
rect 26712 9976 26740 10075
rect 28442 10072 28448 10084
rect 28500 10072 28506 10124
rect 28810 10072 28816 10124
rect 28868 10112 28874 10124
rect 28868 10084 29316 10112
rect 28868 10072 28874 10084
rect 27154 10004 27160 10056
rect 27212 10004 27218 10056
rect 27338 10004 27344 10056
rect 27396 10004 27402 10056
rect 28905 10047 28963 10053
rect 28905 10013 28917 10047
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 28997 10047 29055 10053
rect 28997 10013 29009 10047
rect 29043 10044 29055 10047
rect 29178 10044 29184 10056
rect 29043 10016 29184 10044
rect 29043 10013 29055 10016
rect 28997 10007 29055 10013
rect 27019 9979 27077 9985
rect 27019 9976 27031 9979
rect 26712 9948 27031 9976
rect 25869 9939 25927 9945
rect 27019 9945 27031 9948
rect 27065 9945 27077 9979
rect 27019 9939 27077 9945
rect 27249 9979 27307 9985
rect 27249 9945 27261 9979
rect 27295 9976 27307 9979
rect 27890 9976 27896 9988
rect 27295 9948 27896 9976
rect 27295 9945 27307 9948
rect 27249 9939 27307 9945
rect 11931 9880 13768 9908
rect 11931 9877 11943 9880
rect 11885 9871 11943 9877
rect 16758 9868 16764 9920
rect 16816 9868 16822 9920
rect 23017 9911 23075 9917
rect 23017 9877 23029 9911
rect 23063 9908 23075 9911
rect 23290 9908 23296 9920
rect 23063 9880 23296 9908
rect 23063 9877 23075 9880
rect 23017 9871 23075 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 25130 9868 25136 9920
rect 25188 9868 25194 9920
rect 25314 9868 25320 9920
rect 25372 9908 25378 9920
rect 25424 9908 25452 9939
rect 27890 9936 27896 9948
rect 27948 9976 27954 9988
rect 28920 9976 28948 10007
rect 27948 9948 28948 9976
rect 27948 9936 27954 9948
rect 25958 9908 25964 9920
rect 25372 9880 25964 9908
rect 25372 9868 25378 9880
rect 25958 9868 25964 9880
rect 26016 9868 26022 9920
rect 27522 9868 27528 9920
rect 27580 9868 27586 9920
rect 28258 9868 28264 9920
rect 28316 9908 28322 9920
rect 29012 9908 29040 10007
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 29288 10053 29316 10084
rect 29638 10072 29644 10124
rect 29696 10072 29702 10124
rect 29273 10047 29331 10053
rect 29273 10013 29285 10047
rect 29319 10044 29331 10047
rect 29656 10044 29684 10072
rect 30208 10053 30236 10152
rect 30834 10072 30840 10124
rect 30892 10072 30898 10124
rect 29319 10016 29684 10044
rect 30193 10047 30251 10053
rect 29319 10013 29331 10016
rect 29273 10007 29331 10013
rect 30193 10013 30205 10047
rect 30239 10013 30251 10047
rect 30193 10007 30251 10013
rect 30374 10004 30380 10056
rect 30432 10046 30438 10056
rect 31113 10047 31171 10053
rect 30432 10018 30475 10046
rect 30432 10004 30438 10018
rect 31113 10013 31125 10047
rect 31159 10044 31171 10047
rect 31159 10016 31340 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 31312 9988 31340 10016
rect 31294 9936 31300 9988
rect 31352 9936 31358 9988
rect 28316 9880 29040 9908
rect 28316 9868 28322 9880
rect 1104 9818 38824 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 38824 9818
rect 1104 9744 38824 9766
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 9272 9676 9321 9704
rect 9272 9664 9278 9676
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9309 9667 9367 9673
rect 9766 9664 9772 9716
rect 9824 9664 9830 9716
rect 10502 9664 10508 9716
rect 10560 9664 10566 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 12434 9704 12440 9716
rect 10836 9676 12440 9704
rect 10836 9664 10842 9676
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 12529 9707 12587 9713
rect 12529 9673 12541 9707
rect 12575 9704 12587 9707
rect 12710 9704 12716 9716
rect 12575 9676 12716 9704
rect 12575 9673 12587 9676
rect 12529 9667 12587 9673
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 22186 9664 22192 9716
rect 22244 9664 22250 9716
rect 24026 9664 24032 9716
rect 24084 9664 24090 9716
rect 25774 9664 25780 9716
rect 25832 9664 25838 9716
rect 25958 9664 25964 9716
rect 26016 9704 26022 9716
rect 26016 9676 27936 9704
rect 26016 9664 26022 9676
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9784 9568 9812 9664
rect 9539 9540 9812 9568
rect 10137 9571 10195 9577
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 10137 9537 10149 9571
rect 10183 9568 10195 9571
rect 10520 9568 10548 9664
rect 14645 9639 14703 9645
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 19797 9639 19855 9645
rect 19797 9636 19809 9639
rect 14691 9608 19809 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 19797 9605 19809 9608
rect 19843 9605 19855 9639
rect 19797 9599 19855 9605
rect 23032 9608 23980 9636
rect 10183 9540 10548 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 12161 9571 12219 9577
rect 12161 9568 12173 9571
rect 11572 9540 12173 9568
rect 11572 9528 11578 9540
rect 12161 9537 12173 9540
rect 12207 9568 12219 9571
rect 12207 9540 12434 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9876 9364 9904 9463
rect 12250 9460 12256 9512
rect 12308 9460 12314 9512
rect 12406 9432 12434 9540
rect 13998 9528 14004 9580
rect 14056 9568 14062 9580
rect 14553 9571 14611 9577
rect 14553 9568 14565 9571
rect 14056 9540 14565 9568
rect 14056 9528 14062 9540
rect 14553 9537 14565 9540
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 14752 9500 14780 9531
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 14976 9540 19533 9568
rect 14976 9528 14982 9540
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19702 9528 19708 9580
rect 19760 9528 19766 9580
rect 15930 9500 15936 9512
rect 14752 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 19812 9500 19840 9599
rect 23032 9580 23060 9608
rect 23952 9580 23980 9608
rect 25406 9596 25412 9648
rect 25464 9596 25470 9648
rect 25593 9639 25651 9645
rect 25593 9605 25605 9639
rect 25639 9636 25651 9639
rect 26050 9636 26056 9648
rect 25639 9608 26056 9636
rect 25639 9605 25651 9608
rect 25593 9599 25651 9605
rect 26050 9596 26056 9608
rect 26108 9596 26114 9648
rect 27908 9636 27936 9676
rect 27982 9664 27988 9716
rect 28040 9664 28046 9716
rect 28994 9704 29000 9716
rect 28092 9676 29000 9704
rect 28092 9636 28120 9676
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 29086 9664 29092 9716
rect 29144 9704 29150 9716
rect 30193 9707 30251 9713
rect 30193 9704 30205 9707
rect 29144 9676 30205 9704
rect 29144 9664 29150 9676
rect 30193 9673 30205 9676
rect 30239 9673 30251 9707
rect 30193 9667 30251 9673
rect 30374 9664 30380 9716
rect 30432 9704 30438 9716
rect 31294 9704 31300 9716
rect 30432 9676 31300 9704
rect 30432 9664 30438 9676
rect 31294 9664 31300 9676
rect 31352 9664 31358 9716
rect 30285 9639 30343 9645
rect 27908 9608 28120 9636
rect 28368 9608 29960 9636
rect 19886 9528 19892 9580
rect 19944 9528 19950 9580
rect 22002 9528 22008 9580
rect 22060 9568 22066 9580
rect 22097 9571 22155 9577
rect 22097 9568 22109 9571
rect 22060 9540 22109 9568
rect 22060 9528 22066 9540
rect 22097 9537 22109 9540
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 23014 9528 23020 9580
rect 23072 9528 23078 9580
rect 23290 9528 23296 9580
rect 23348 9528 23354 9580
rect 23934 9528 23940 9580
rect 23992 9528 23998 9580
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9537 28043 9571
rect 27985 9531 28043 9537
rect 28000 9500 28028 9531
rect 28166 9528 28172 9580
rect 28224 9528 28230 9580
rect 28258 9500 28264 9512
rect 19812 9472 22094 9500
rect 28000 9472 28264 9500
rect 14550 9432 14556 9444
rect 12406 9404 14556 9432
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 10318 9364 10324 9376
rect 9876 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9364 10382 9376
rect 10686 9364 10692 9376
rect 10376 9336 10692 9364
rect 10376 9324 10382 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 10873 9367 10931 9373
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 10962 9364 10968 9376
rect 10919 9336 10968 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 14366 9324 14372 9376
rect 14424 9324 14430 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 18046 9364 18052 9376
rect 15528 9336 18052 9364
rect 15528 9324 15534 9336
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 20070 9324 20076 9376
rect 20128 9324 20134 9376
rect 22066 9364 22094 9472
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 28368 9432 28396 9608
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 29595 9540 29868 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 29840 9441 29868 9540
rect 29932 9500 29960 9608
rect 30285 9605 30297 9639
rect 30331 9636 30343 9639
rect 30392 9636 30420 9664
rect 30331 9608 30420 9636
rect 30331 9605 30343 9608
rect 30285 9599 30343 9605
rect 30377 9503 30435 9509
rect 30377 9500 30389 9503
rect 29932 9472 30389 9500
rect 30377 9469 30389 9472
rect 30423 9469 30435 9503
rect 30377 9463 30435 9469
rect 27396 9404 28396 9432
rect 29825 9435 29883 9441
rect 27396 9392 27402 9404
rect 29825 9401 29837 9435
rect 29871 9401 29883 9435
rect 29825 9395 29883 9401
rect 25314 9364 25320 9376
rect 22066 9336 25320 9364
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 29638 9324 29644 9376
rect 29696 9364 29702 9376
rect 29733 9367 29791 9373
rect 29733 9364 29745 9367
rect 29696 9336 29745 9364
rect 29696 9324 29702 9336
rect 29733 9333 29745 9336
rect 29779 9333 29791 9367
rect 29733 9327 29791 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 11514 9120 11520 9172
rect 11572 9120 11578 9172
rect 14550 9120 14556 9172
rect 14608 9120 14614 9172
rect 15289 9163 15347 9169
rect 15289 9129 15301 9163
rect 15335 9160 15347 9163
rect 15470 9160 15476 9172
rect 15335 9132 15476 9160
rect 15335 9129 15347 9132
rect 15289 9123 15347 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 15930 9120 15936 9172
rect 15988 9120 15994 9172
rect 16942 9120 16948 9172
rect 17000 9120 17006 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 18417 9163 18475 9169
rect 17276 9132 18368 9160
rect 17276 9120 17282 9132
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 10686 8956 10692 8968
rect 10551 8928 10692 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10827 8928 11008 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10980 8832 11008 8928
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 14568 8965 14596 9120
rect 14737 9095 14795 9101
rect 14737 9061 14749 9095
rect 14783 9061 14795 9095
rect 17865 9095 17923 9101
rect 17865 9092 17877 9095
rect 14737 9055 14795 9061
rect 15672 9064 17877 9092
rect 14752 9024 14780 9055
rect 14752 8996 15608 9024
rect 15580 8965 15608 8996
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 12308 8928 14473 8956
rect 12308 8916 12314 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8956 14611 8959
rect 15565 8959 15623 8965
rect 14599 8928 14872 8956
rect 14599 8925 14611 8928
rect 14553 8919 14611 8925
rect 10962 8780 10968 8832
rect 11020 8780 11026 8832
rect 14476 8820 14504 8919
rect 14734 8848 14740 8900
rect 14792 8848 14798 8900
rect 14844 8888 14872 8928
rect 15565 8925 15577 8959
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 15105 8891 15163 8897
rect 15105 8888 15117 8891
rect 14844 8860 15117 8888
rect 15105 8857 15117 8860
rect 15151 8888 15163 8891
rect 15672 8888 15700 9064
rect 17865 9061 17877 9064
rect 17911 9061 17923 9095
rect 18340 9092 18368 9132
rect 18417 9129 18429 9163
rect 18463 9160 18475 9163
rect 18966 9160 18972 9172
rect 18463 9132 18972 9160
rect 18463 9129 18475 9132
rect 18417 9123 18475 9129
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19061 9163 19119 9169
rect 19061 9129 19073 9163
rect 19107 9160 19119 9163
rect 19702 9160 19708 9172
rect 19107 9132 19708 9160
rect 19107 9129 19119 9132
rect 19061 9123 19119 9129
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 20070 9120 20076 9172
rect 20128 9120 20134 9172
rect 25608 9132 26280 9160
rect 18340 9064 19656 9092
rect 17865 9055 17923 9061
rect 19628 9033 19656 9064
rect 17221 9027 17279 9033
rect 16408 8996 17172 9024
rect 16408 8965 16436 8996
rect 17144 8965 17172 8996
rect 17221 8993 17233 9027
rect 17267 9024 17279 9027
rect 18601 9027 18659 9033
rect 18601 9024 18613 9027
rect 17267 8996 18613 9024
rect 17267 8993 17279 8996
rect 17221 8987 17279 8993
rect 18601 8993 18613 8996
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 8993 19671 9027
rect 19613 8987 19671 8993
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15795 8928 16405 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16393 8925 16405 8928
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16807 8928 16865 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 17129 8959 17187 8965
rect 17129 8925 17141 8959
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 15151 8860 15700 8888
rect 15151 8857 15163 8860
rect 15105 8851 15163 8857
rect 15305 8823 15363 8829
rect 15305 8820 15317 8823
rect 14476 8792 15317 8820
rect 15305 8789 15317 8792
rect 15351 8789 15363 8823
rect 15305 8783 15363 8789
rect 15473 8823 15531 8829
rect 15473 8789 15485 8823
rect 15519 8820 15531 8823
rect 15764 8820 15792 8919
rect 16577 8891 16635 8897
rect 16577 8857 16589 8891
rect 16623 8857 16635 8891
rect 17052 8888 17080 8919
rect 17236 8888 17264 8987
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17678 8956 17684 8968
rect 17635 8928 17684 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17052 8860 17264 8888
rect 17328 8888 17356 8919
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 17770 8916 17776 8968
rect 17828 8916 17834 8968
rect 18046 8916 18052 8968
rect 18104 8916 18110 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18693 8959 18751 8965
rect 18693 8956 18705 8959
rect 18279 8928 18705 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18693 8925 18705 8928
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20088 8956 20116 9120
rect 20254 9052 20260 9104
rect 20312 9052 20318 9104
rect 24397 9095 24455 9101
rect 24397 9061 24409 9095
rect 24443 9061 24455 9095
rect 24397 9055 24455 9061
rect 21082 8984 21088 9036
rect 21140 8984 21146 9036
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 23014 9024 23020 9036
rect 22152 8996 23020 9024
rect 22152 8984 22158 8996
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 19935 8928 20116 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 18138 8888 18144 8900
rect 17328 8860 18144 8888
rect 16577 8851 16635 8857
rect 15519 8792 15792 8820
rect 16592 8820 16620 8851
rect 17328 8820 17356 8860
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 16592 8792 17356 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17552 8792 17693 8820
rect 17552 8780 17558 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 18708 8820 18736 8919
rect 19797 8891 19855 8897
rect 19797 8857 19809 8891
rect 19843 8888 19855 8891
rect 21100 8888 21128 8984
rect 21821 8959 21879 8965
rect 21821 8956 21833 8959
rect 19843 8860 21128 8888
rect 21284 8928 21833 8956
rect 19843 8857 19855 8860
rect 19797 8851 19855 8857
rect 21284 8832 21312 8928
rect 21821 8925 21833 8928
rect 21867 8925 21879 8959
rect 21821 8919 21879 8925
rect 23385 8959 23443 8965
rect 23385 8925 23397 8959
rect 23431 8956 23443 8959
rect 24412 8956 24440 9055
rect 25222 9052 25228 9104
rect 25280 9052 25286 9104
rect 24486 8984 24492 9036
rect 24544 9024 24550 9036
rect 25041 9027 25099 9033
rect 25041 9024 25053 9027
rect 24544 8996 25053 9024
rect 24544 8984 24550 8996
rect 25041 8993 25053 8996
rect 25087 9024 25099 9027
rect 25608 9024 25636 9132
rect 26050 9092 26056 9104
rect 25700 9064 26056 9092
rect 25700 9033 25728 9064
rect 26050 9052 26056 9064
rect 26108 9092 26114 9104
rect 26145 9095 26203 9101
rect 26145 9092 26157 9095
rect 26108 9064 26157 9092
rect 26108 9052 26114 9064
rect 26145 9061 26157 9064
rect 26191 9061 26203 9095
rect 26145 9055 26203 9061
rect 25087 8996 25636 9024
rect 25685 9027 25743 9033
rect 25087 8993 25099 8996
rect 25041 8987 25099 8993
rect 25685 8993 25697 9027
rect 25731 8993 25743 9027
rect 26252 9024 26280 9132
rect 28166 9120 28172 9172
rect 28224 9160 28230 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 28224 9132 28457 9160
rect 28224 9120 28230 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 28445 9123 28503 9129
rect 29638 9120 29644 9172
rect 29696 9120 29702 9172
rect 31294 9120 31300 9172
rect 31352 9120 31358 9172
rect 26602 9052 26608 9104
rect 26660 9092 26666 9104
rect 27430 9092 27436 9104
rect 26660 9064 27436 9092
rect 26660 9052 26666 9064
rect 27430 9052 27436 9064
rect 27488 9092 27494 9104
rect 28626 9092 28632 9104
rect 27488 9064 28632 9092
rect 27488 9052 27494 9064
rect 28626 9052 28632 9064
rect 28684 9092 28690 9104
rect 29181 9095 29239 9101
rect 29181 9092 29193 9095
rect 28684 9064 29193 9092
rect 28684 9052 28690 9064
rect 29181 9061 29193 9064
rect 29227 9061 29239 9095
rect 29181 9055 29239 9061
rect 27338 9024 27344 9036
rect 26252 8996 27344 9024
rect 25685 8987 25743 8993
rect 27338 8984 27344 8996
rect 27396 8984 27402 9036
rect 29656 9024 29684 9120
rect 29825 9027 29883 9033
rect 29825 9024 29837 9027
rect 27908 8996 28580 9024
rect 29656 8996 29837 9024
rect 23431 8928 24440 8956
rect 24765 8959 24823 8965
rect 23431 8925 23443 8928
rect 23385 8919 23443 8925
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 25130 8956 25136 8968
rect 24811 8928 25136 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 27065 8959 27123 8965
rect 27065 8925 27077 8959
rect 27111 8956 27123 8959
rect 27522 8956 27528 8968
rect 27111 8928 27528 8956
rect 27111 8925 27123 8928
rect 27065 8919 27123 8925
rect 25608 8888 25636 8919
rect 27522 8916 27528 8928
rect 27580 8916 27586 8968
rect 27908 8897 27936 8996
rect 28258 8916 28264 8968
rect 28316 8916 28322 8968
rect 28552 8965 28580 8996
rect 29825 8993 29837 8996
rect 29871 8993 29883 9027
rect 29825 8987 29883 8993
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 28537 8959 28595 8965
rect 28537 8925 28549 8959
rect 28583 8925 28595 8959
rect 28537 8919 28595 8925
rect 25869 8891 25927 8897
rect 25869 8888 25881 8891
rect 24872 8860 25881 8888
rect 20990 8820 20996 8832
rect 18708 8792 20996 8820
rect 17681 8783 17739 8789
rect 20990 8780 20996 8792
rect 21048 8820 21054 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 21048 8792 21097 8820
rect 21048 8780 21054 8792
rect 21085 8789 21097 8792
rect 21131 8789 21143 8823
rect 21085 8783 21143 8789
rect 21266 8780 21272 8832
rect 21324 8780 21330 8832
rect 23198 8780 23204 8832
rect 23256 8780 23262 8832
rect 24670 8780 24676 8832
rect 24728 8820 24734 8832
rect 24872 8829 24900 8860
rect 25869 8857 25881 8860
rect 25915 8857 25927 8891
rect 27893 8891 27951 8897
rect 27893 8888 27905 8891
rect 25869 8851 25927 8857
rect 26344 8860 27905 8888
rect 26344 8829 26372 8860
rect 27893 8857 27905 8860
rect 27939 8857 27951 8891
rect 27893 8851 27951 8857
rect 28077 8891 28135 8897
rect 28077 8857 28089 8891
rect 28123 8888 28135 8891
rect 28368 8888 28396 8919
rect 28994 8916 29000 8968
rect 29052 8956 29058 8968
rect 29546 8956 29552 8968
rect 29052 8928 29552 8956
rect 29052 8916 29058 8928
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 28123 8860 28396 8888
rect 28123 8857 28135 8860
rect 28077 8851 28135 8857
rect 24857 8823 24915 8829
rect 24857 8820 24869 8823
rect 24728 8792 24869 8820
rect 24728 8780 24734 8792
rect 24857 8789 24869 8792
rect 24903 8789 24915 8823
rect 24857 8783 24915 8789
rect 26329 8823 26387 8829
rect 26329 8789 26341 8823
rect 26375 8789 26387 8823
rect 26329 8783 26387 8789
rect 26694 8780 26700 8832
rect 26752 8780 26758 8832
rect 27157 8823 27215 8829
rect 27157 8789 27169 8823
rect 27203 8820 27215 8823
rect 27614 8820 27620 8832
rect 27203 8792 27620 8820
rect 27203 8789 27215 8792
rect 27157 8783 27215 8789
rect 27614 8780 27620 8792
rect 27672 8780 27678 8832
rect 27982 8780 27988 8832
rect 28040 8820 28046 8832
rect 28092 8820 28120 8851
rect 28902 8848 28908 8900
rect 28960 8848 28966 8900
rect 30098 8848 30104 8900
rect 30156 8888 30162 8900
rect 30156 8860 30314 8888
rect 30156 8848 30162 8860
rect 28040 8792 28120 8820
rect 29365 8823 29423 8829
rect 28040 8780 28046 8792
rect 29365 8789 29377 8823
rect 29411 8820 29423 8823
rect 29822 8820 29828 8832
rect 29411 8792 29828 8820
rect 29411 8789 29423 8792
rect 29365 8783 29423 8789
rect 29822 8780 29828 8792
rect 29880 8780 29886 8832
rect 1104 8730 38824 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 38824 8730
rect 1104 8656 38824 8678
rect 15010 8616 15016 8628
rect 11624 8588 15016 8616
rect 11624 8489 11652 8588
rect 15010 8576 15016 8588
rect 15068 8616 15074 8628
rect 15562 8616 15568 8628
rect 15068 8588 15568 8616
rect 15068 8576 15074 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 16758 8576 16764 8628
rect 16816 8616 16822 8628
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 16816 8588 17049 8616
rect 16816 8576 16822 8588
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 17828 8588 18337 8616
rect 17828 8576 17834 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 19536 8588 21864 8616
rect 12618 8508 12624 8560
rect 12676 8508 12682 8560
rect 13817 8551 13875 8557
rect 13817 8517 13829 8551
rect 13863 8548 13875 8551
rect 14366 8548 14372 8560
rect 13863 8520 14372 8548
rect 13863 8517 13875 8520
rect 13817 8511 13875 8517
rect 14366 8508 14372 8520
rect 14424 8508 14430 8560
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 18785 8551 18843 8557
rect 18785 8548 18797 8551
rect 18196 8520 18797 8548
rect 18196 8508 18202 8520
rect 18785 8517 18797 8520
rect 18831 8517 18843 8551
rect 19536 8548 19564 8588
rect 21361 8551 21419 8557
rect 21361 8548 21373 8551
rect 18785 8511 18843 8517
rect 19444 8520 19564 8548
rect 20930 8520 21373 8548
rect 19444 8489 19472 8520
rect 21361 8517 21373 8520
rect 21407 8517 21419 8551
rect 21361 8511 21419 8517
rect 21836 8492 21864 8588
rect 23198 8576 23204 8628
rect 23256 8576 23262 8628
rect 26050 8576 26056 8628
rect 26108 8616 26114 8628
rect 26513 8619 26571 8625
rect 26513 8616 26525 8619
rect 26108 8588 26525 8616
rect 26108 8576 26114 8588
rect 26513 8585 26525 8588
rect 26559 8585 26571 8619
rect 26513 8579 26571 8585
rect 26694 8576 26700 8628
rect 26752 8576 26758 8628
rect 27893 8619 27951 8625
rect 27893 8585 27905 8619
rect 27939 8616 27951 8619
rect 27982 8616 27988 8628
rect 27939 8588 27988 8616
rect 27939 8585 27951 8588
rect 27893 8579 27951 8585
rect 27982 8576 27988 8588
rect 28040 8576 28046 8628
rect 28626 8576 28632 8628
rect 28684 8576 28690 8628
rect 30098 8576 30104 8628
rect 30156 8576 30162 8628
rect 22833 8551 22891 8557
rect 22833 8517 22845 8551
rect 22879 8548 22891 8551
rect 23216 8548 23244 8576
rect 22879 8520 23244 8548
rect 22879 8517 22891 8520
rect 22833 8511 22891 8517
rect 23566 8508 23572 8560
rect 23624 8508 23630 8560
rect 25590 8548 25596 8560
rect 24228 8520 25596 8548
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8449 11667 8483
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 11609 8443 11667 8449
rect 13924 8452 14657 8480
rect 11882 8372 11888 8424
rect 11940 8372 11946 8424
rect 13924 8421 13952 8452
rect 14645 8449 14657 8452
rect 14691 8480 14703 8483
rect 14921 8483 14979 8489
rect 14921 8480 14933 8483
rect 14691 8452 14933 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 14921 8449 14933 8452
rect 14967 8449 14979 8483
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 14921 8443 14979 8449
rect 17144 8452 18245 8480
rect 17144 8424 17172 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13740 8384 13921 8412
rect 13446 8304 13452 8356
rect 13504 8304 13510 8356
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 13357 8279 13415 8285
rect 13357 8276 13369 8279
rect 13228 8248 13369 8276
rect 13228 8236 13234 8248
rect 13357 8245 13369 8248
rect 13403 8276 13415 8279
rect 13740 8276 13768 8384
rect 13909 8381 13921 8384
rect 13955 8381 13967 8415
rect 13909 8375 13967 8381
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8412 14151 8415
rect 14139 8384 14688 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14274 8304 14280 8356
rect 14332 8304 14338 8356
rect 14660 8344 14688 8384
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 15381 8415 15439 8421
rect 14792 8384 15332 8412
rect 14792 8372 14798 8384
rect 15304 8353 15332 8384
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 16850 8412 16856 8424
rect 15427 8384 16856 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 16850 8372 16856 8384
rect 16908 8372 16914 8424
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17218 8372 17224 8424
rect 17276 8372 17282 8424
rect 17678 8372 17684 8424
rect 17736 8412 17742 8424
rect 17773 8415 17831 8421
rect 17773 8412 17785 8415
rect 17736 8384 17785 8412
rect 17736 8372 17742 8384
rect 17773 8381 17785 8384
rect 17819 8412 17831 8415
rect 17954 8412 17960 8424
rect 17819 8384 17960 8412
rect 17819 8381 17831 8384
rect 17773 8375 17831 8381
rect 17954 8372 17960 8384
rect 18012 8372 18018 8424
rect 15289 8347 15347 8353
rect 14660 8316 15240 8344
rect 13403 8248 13768 8276
rect 15212 8276 15240 8316
rect 15289 8313 15301 8347
rect 15335 8344 15347 8347
rect 15470 8344 15476 8356
rect 15335 8316 15476 8344
rect 15335 8313 15347 8316
rect 15289 8307 15347 8313
rect 15470 8304 15476 8316
rect 15528 8304 15534 8356
rect 17236 8344 17264 8372
rect 15580 8316 17264 8344
rect 17865 8347 17923 8353
rect 15580 8276 15608 8316
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 18138 8344 18144 8356
rect 17911 8316 18144 8344
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 18248 8344 18276 8443
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 21818 8440 21824 8492
rect 21876 8480 21882 8492
rect 22557 8483 22615 8489
rect 22557 8480 22569 8483
rect 21876 8452 22569 8480
rect 21876 8440 21882 8452
rect 22557 8449 22569 8452
rect 22603 8449 22615 8483
rect 22557 8443 22615 8449
rect 19702 8372 19708 8424
rect 19760 8372 19766 8424
rect 21100 8412 21128 8440
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 21100 8384 21189 8412
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 21468 8412 21496 8440
rect 22002 8412 22008 8424
rect 21468 8384 22008 8412
rect 21177 8375 21235 8381
rect 22002 8372 22008 8384
rect 22060 8412 22066 8424
rect 23474 8412 23480 8424
rect 22060 8384 23480 8412
rect 22060 8372 22066 8384
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 18417 8347 18475 8353
rect 18417 8344 18429 8347
rect 18248 8316 18429 8344
rect 18417 8313 18429 8316
rect 18463 8313 18475 8347
rect 24228 8344 24256 8520
rect 25590 8508 25596 8520
rect 25648 8548 25654 8560
rect 25648 8520 26648 8548
rect 25648 8508 25654 8520
rect 24670 8480 24676 8492
rect 24320 8452 24676 8480
rect 24320 8421 24348 8452
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 25777 8483 25835 8489
rect 25777 8480 25789 8483
rect 25424 8452 25789 8480
rect 24305 8415 24363 8421
rect 24305 8381 24317 8415
rect 24351 8381 24363 8415
rect 24305 8375 24363 8381
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8381 24455 8415
rect 24397 8375 24455 8381
rect 24412 8344 24440 8375
rect 24228 8316 24440 8344
rect 18417 8307 18475 8313
rect 25130 8304 25136 8356
rect 25188 8344 25194 8356
rect 25424 8353 25452 8452
rect 25777 8449 25789 8452
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 25498 8372 25504 8424
rect 25556 8372 25562 8424
rect 25409 8347 25467 8353
rect 25409 8344 25421 8347
rect 25188 8316 25421 8344
rect 25188 8304 25194 8316
rect 25409 8313 25421 8316
rect 25455 8313 25467 8347
rect 26620 8344 26648 8520
rect 26712 8480 26740 8576
rect 30466 8548 30472 8560
rect 29012 8520 30472 8548
rect 26789 8483 26847 8489
rect 26789 8480 26801 8483
rect 26712 8452 26801 8480
rect 26789 8449 26801 8452
rect 26835 8449 26847 8483
rect 26789 8443 26847 8449
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8480 27583 8483
rect 27614 8480 27620 8492
rect 27571 8452 27620 8480
rect 27571 8449 27583 8452
rect 27525 8443 27583 8449
rect 27614 8440 27620 8452
rect 27672 8480 27678 8492
rect 28902 8480 28908 8492
rect 27672 8452 28908 8480
rect 27672 8440 27678 8452
rect 28902 8440 28908 8452
rect 28960 8440 28966 8492
rect 27430 8372 27436 8424
rect 27488 8372 27494 8424
rect 29012 8412 29040 8520
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 29656 8489 29684 8520
rect 30466 8508 30472 8520
rect 30524 8508 30530 8560
rect 29365 8483 29423 8489
rect 29365 8480 29377 8483
rect 29236 8452 29377 8480
rect 29236 8440 29242 8452
rect 29365 8449 29377 8452
rect 29411 8449 29423 8483
rect 29365 8443 29423 8449
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 29641 8443 29699 8449
rect 29730 8440 29736 8492
rect 29788 8480 29794 8492
rect 30009 8483 30067 8489
rect 30009 8480 30021 8483
rect 29788 8452 30021 8480
rect 29788 8440 29794 8452
rect 30009 8449 30021 8452
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 38194 8440 38200 8492
rect 38252 8440 38258 8492
rect 28000 8384 29040 8412
rect 28000 8356 28028 8384
rect 27982 8344 27988 8356
rect 26620 8316 27988 8344
rect 25409 8307 25467 8313
rect 27982 8304 27988 8316
rect 28040 8304 28046 8356
rect 38378 8304 38384 8356
rect 38436 8304 38442 8356
rect 15212 8248 15608 8276
rect 13403 8245 13415 8248
rect 13357 8239 13415 8245
rect 16666 8236 16672 8288
rect 16724 8236 16730 8288
rect 26602 8236 26608 8288
rect 26660 8236 26666 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11940 8044 12265 8072
rect 11940 8032 11946 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 12618 8032 12624 8084
rect 12676 8032 12682 8084
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 15470 8072 15476 8084
rect 15243 8044 15476 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17184 8044 17325 8072
rect 17184 8032 17190 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18138 8072 18144 8084
rect 18003 8044 18144 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18432 8044 19656 8072
rect 10686 7964 10692 8016
rect 10744 8004 10750 8016
rect 18432 8004 18460 8044
rect 10744 7976 12940 8004
rect 10744 7964 10750 7976
rect 12413 7867 12471 7873
rect 12413 7833 12425 7867
rect 12459 7864 12471 7867
rect 12537 7871 12595 7877
rect 12459 7833 12472 7864
rect 12413 7827 12472 7833
rect 12537 7837 12549 7871
rect 12583 7868 12595 7871
rect 12710 7868 12716 7880
rect 12583 7840 12716 7868
rect 12583 7837 12595 7840
rect 12537 7831 12595 7837
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12912 7877 12940 7976
rect 17604 7976 18460 8004
rect 19628 8004 19656 8044
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 19981 8075 20039 8081
rect 19981 8072 19993 8075
rect 19760 8044 19993 8072
rect 19760 8032 19766 8044
rect 19981 8041 19993 8044
rect 20027 8041 20039 8075
rect 21450 8072 21456 8084
rect 19981 8035 20039 8041
rect 20732 8044 21456 8072
rect 20732 8004 20760 8044
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 23566 8032 23572 8084
rect 23624 8032 23630 8084
rect 28994 8072 29000 8084
rect 26252 8044 29000 8072
rect 19628 7976 20760 8004
rect 15562 7896 15568 7948
rect 15620 7896 15626 7948
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12444 7800 12472 7827
rect 12912 7800 12940 7831
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 17604 7877 17632 7976
rect 20625 7939 20683 7945
rect 20625 7936 20637 7939
rect 18984 7908 20637 7936
rect 18984 7877 19012 7908
rect 20625 7905 20637 7908
rect 20671 7905 20683 7939
rect 22094 7936 22100 7948
rect 20625 7899 20683 7905
rect 21192 7908 22100 7936
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13280 7840 14197 7868
rect 13280 7800 13308 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7837 17647 7871
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 17589 7831 17647 7837
rect 18064 7840 18705 7868
rect 12444 7772 12572 7800
rect 12912 7772 13308 7800
rect 12544 7732 12572 7772
rect 13446 7760 13452 7812
rect 13504 7760 13510 7812
rect 14476 7800 14504 7831
rect 14200 7772 14504 7800
rect 13464 7732 13492 7760
rect 14200 7744 14228 7772
rect 15838 7760 15844 7812
rect 15896 7760 15902 7812
rect 17497 7803 17555 7809
rect 17497 7800 17509 7803
rect 17066 7772 17509 7800
rect 17497 7769 17509 7772
rect 17543 7769 17555 7803
rect 17497 7763 17555 7769
rect 18064 7744 18092 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7837 19027 7871
rect 18969 7831 19027 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20254 7868 20260 7880
rect 20211 7840 20260 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 18322 7760 18328 7812
rect 18380 7800 18386 7812
rect 18984 7800 19012 7831
rect 20254 7828 20260 7840
rect 20312 7828 20318 7880
rect 18380 7772 19012 7800
rect 18380 7760 18386 7772
rect 12544 7704 13492 7732
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 14182 7732 14188 7744
rect 13955 7704 14188 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 20640 7732 20668 7899
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 20947 7840 21128 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 21100 7812 21128 7840
rect 21082 7760 21088 7812
rect 21140 7760 21146 7812
rect 21192 7732 21220 7908
rect 22094 7896 22100 7908
rect 22152 7896 22158 7948
rect 26252 7945 26280 8044
rect 28994 8032 29000 8044
rect 29052 8032 29058 8084
rect 26237 7939 26295 7945
rect 26237 7905 26249 7939
rect 26283 7905 26295 7939
rect 26237 7899 26295 7905
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 26602 7936 26608 7948
rect 26559 7908 26608 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 26602 7896 26608 7908
rect 26660 7896 26666 7948
rect 27982 7896 27988 7948
rect 28040 7936 28046 7948
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 28040 7908 28089 7936
rect 28040 7896 28046 7908
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28077 7899 28135 7905
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 28353 7871 28411 7877
rect 28353 7837 28365 7871
rect 28399 7868 28411 7871
rect 28902 7868 28908 7880
rect 28399 7840 28908 7868
rect 28399 7837 28411 7840
rect 28353 7831 28411 7837
rect 27246 7760 27252 7812
rect 27304 7760 27310 7812
rect 20640 7704 21220 7732
rect 21266 7692 21272 7744
rect 21324 7732 21330 7744
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21324 7704 21649 7732
rect 21324 7692 21330 7704
rect 21637 7701 21649 7704
rect 21683 7701 21695 7735
rect 21637 7695 21695 7701
rect 27985 7735 28043 7741
rect 27985 7701 27997 7735
rect 28031 7732 28043 7735
rect 28368 7732 28396 7831
rect 28902 7828 28908 7840
rect 28960 7828 28966 7880
rect 28031 7704 28396 7732
rect 28031 7701 28043 7704
rect 27985 7695 28043 7701
rect 28994 7692 29000 7744
rect 29052 7732 29058 7744
rect 29089 7735 29147 7741
rect 29089 7732 29101 7735
rect 29052 7704 29101 7732
rect 29052 7692 29058 7704
rect 29089 7701 29101 7704
rect 29135 7732 29147 7735
rect 29178 7732 29184 7744
rect 29135 7704 29184 7732
rect 29135 7701 29147 7704
rect 29089 7695 29147 7701
rect 29178 7692 29184 7704
rect 29236 7692 29242 7744
rect 1104 7642 38824 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 38824 7642
rect 1104 7568 38824 7590
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 16025 7531 16083 7537
rect 16025 7528 16037 7531
rect 15896 7500 16037 7528
rect 15896 7488 15902 7500
rect 16025 7497 16037 7500
rect 16071 7497 16083 7531
rect 16025 7491 16083 7497
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 17126 7488 17132 7540
rect 17184 7488 17190 7540
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 27341 7531 27399 7537
rect 27341 7528 27353 7531
rect 27304 7500 27353 7528
rect 27304 7488 27310 7500
rect 27341 7497 27353 7500
rect 27387 7497 27399 7531
rect 27341 7491 27399 7497
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16684 7392 16712 7488
rect 16255 7364 16712 7392
rect 17144 7392 17172 7488
rect 17589 7395 17647 7401
rect 17589 7392 17601 7395
rect 17144 7364 17601 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 17589 7361 17601 7364
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 18322 7352 18328 7404
rect 18380 7352 18386 7404
rect 23492 7392 23520 7488
rect 27249 7395 27307 7401
rect 27249 7392 27261 7395
rect 23492 7364 27261 7392
rect 27249 7361 27261 7364
rect 27295 7392 27307 7395
rect 29730 7392 29736 7404
rect 27295 7364 29736 7392
rect 27295 7361 27307 7364
rect 27249 7355 27307 7361
rect 29730 7352 29736 7364
rect 29788 7352 29794 7404
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17328 7256 17356 7287
rect 18340 7256 18368 7352
rect 17328 7228 17448 7256
rect 17420 7188 17448 7228
rect 17972 7228 18368 7256
rect 17972 7188 18000 7228
rect 17420 7160 18000 7188
rect 18046 7148 18052 7200
rect 18104 7188 18110 7200
rect 18325 7191 18383 7197
rect 18325 7188 18337 7191
rect 18104 7160 18337 7188
rect 18104 7148 18110 7160
rect 18325 7157 18337 7160
rect 18371 7157 18383 7191
rect 18325 7151 18383 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1104 5466 38824 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1104 2202 38824 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 15476 37408 15528 37460
rect 17408 37408 17460 37460
rect 19340 37408 19392 37460
rect 21916 37408 21968 37460
rect 15660 37179 15712 37188
rect 15660 37145 15669 37179
rect 15669 37145 15703 37179
rect 15703 37145 15712 37179
rect 15660 37136 15712 37145
rect 17316 37136 17368 37188
rect 19524 37179 19576 37188
rect 19524 37145 19533 37179
rect 19533 37145 19567 37179
rect 19567 37145 19576 37179
rect 19524 37136 19576 37145
rect 22376 37179 22428 37188
rect 22376 37145 22385 37179
rect 22385 37145 22419 37179
rect 22419 37145 22428 37179
rect 22376 37136 22428 37145
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 7564 31263 7616 31272
rect 7564 31229 7573 31263
rect 7573 31229 7607 31263
rect 7607 31229 7616 31263
rect 7564 31220 7616 31229
rect 8208 31127 8260 31136
rect 8208 31093 8217 31127
rect 8217 31093 8251 31127
rect 8251 31093 8260 31127
rect 8208 31084 8260 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7564 30880 7616 30932
rect 8208 30880 8260 30932
rect 7840 30744 7892 30796
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 7196 30676 7248 30685
rect 7472 30719 7524 30728
rect 7472 30685 7481 30719
rect 7481 30685 7515 30719
rect 7515 30685 7524 30719
rect 7472 30676 7524 30685
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 10600 30676 10652 30685
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 12256 30719 12308 30728
rect 12256 30685 12265 30719
rect 12265 30685 12299 30719
rect 12299 30685 12308 30719
rect 12256 30676 12308 30685
rect 15568 30676 15620 30728
rect 6368 30583 6420 30592
rect 6368 30549 6377 30583
rect 6377 30549 6411 30583
rect 6411 30549 6420 30583
rect 6368 30540 6420 30549
rect 7104 30540 7156 30592
rect 8392 30583 8444 30592
rect 8392 30549 8401 30583
rect 8401 30549 8435 30583
rect 8435 30549 8444 30583
rect 8392 30540 8444 30549
rect 8484 30540 8536 30592
rect 10784 30583 10836 30592
rect 10784 30549 10793 30583
rect 10793 30549 10827 30583
rect 10827 30549 10836 30583
rect 10784 30540 10836 30549
rect 11244 30583 11296 30592
rect 11244 30549 11253 30583
rect 11253 30549 11287 30583
rect 11287 30549 11296 30583
rect 11244 30540 11296 30549
rect 12900 30583 12952 30592
rect 12900 30549 12909 30583
rect 12909 30549 12943 30583
rect 12943 30549 12952 30583
rect 12900 30540 12952 30549
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 7472 30379 7524 30388
rect 7472 30345 7481 30379
rect 7481 30345 7515 30379
rect 7515 30345 7524 30379
rect 7472 30336 7524 30345
rect 10600 30336 10652 30388
rect 12256 30336 12308 30388
rect 8392 30268 8444 30320
rect 11244 30268 11296 30320
rect 11796 30268 11848 30320
rect 6368 30200 6420 30252
rect 11152 30200 11204 30252
rect 12716 30200 12768 30252
rect 13728 30200 13780 30252
rect 11060 30132 11112 30184
rect 12440 30175 12492 30184
rect 12440 30141 12449 30175
rect 12449 30141 12483 30175
rect 12483 30141 12492 30175
rect 12440 30132 12492 30141
rect 7380 29996 7432 30048
rect 12348 29996 12400 30048
rect 15568 30132 15620 30184
rect 17592 30200 17644 30252
rect 14096 29996 14148 30048
rect 15752 29996 15804 30048
rect 18144 29996 18196 30048
rect 19984 29996 20036 30048
rect 21548 30039 21600 30048
rect 21548 30005 21557 30039
rect 21557 30005 21591 30039
rect 21591 30005 21600 30039
rect 21548 29996 21600 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12440 29792 12492 29844
rect 12716 29792 12768 29844
rect 7840 29767 7892 29776
rect 7840 29733 7849 29767
rect 7849 29733 7883 29767
rect 7883 29733 7892 29767
rect 7840 29724 7892 29733
rect 12900 29656 12952 29708
rect 5816 29631 5868 29640
rect 5816 29597 5825 29631
rect 5825 29597 5859 29631
rect 5859 29597 5868 29631
rect 5816 29588 5868 29597
rect 6276 29588 6328 29640
rect 7380 29631 7432 29640
rect 7380 29597 7398 29631
rect 7398 29597 7432 29631
rect 7380 29588 7432 29597
rect 6092 29520 6144 29572
rect 7196 29520 7248 29572
rect 5356 29452 5408 29504
rect 6000 29495 6052 29504
rect 6000 29461 6009 29495
rect 6009 29461 6043 29495
rect 6043 29461 6052 29495
rect 6000 29452 6052 29461
rect 7104 29452 7156 29504
rect 8300 29588 8352 29640
rect 8484 29563 8536 29572
rect 8484 29529 8493 29563
rect 8493 29529 8527 29563
rect 8527 29529 8536 29563
rect 9680 29588 9732 29640
rect 17592 29792 17644 29844
rect 13728 29656 13780 29708
rect 14096 29656 14148 29708
rect 8484 29520 8536 29529
rect 9588 29520 9640 29572
rect 8668 29452 8720 29504
rect 10784 29520 10836 29572
rect 13268 29631 13320 29640
rect 13268 29597 13277 29631
rect 13277 29597 13311 29631
rect 13311 29597 13320 29631
rect 13268 29588 13320 29597
rect 15752 29588 15804 29640
rect 19984 29588 20036 29640
rect 21548 29588 21600 29640
rect 14740 29563 14792 29572
rect 14740 29529 14749 29563
rect 14749 29529 14783 29563
rect 14783 29529 14792 29563
rect 14740 29520 14792 29529
rect 16488 29563 16540 29572
rect 16488 29529 16497 29563
rect 16497 29529 16531 29563
rect 16531 29529 16540 29563
rect 16488 29520 16540 29529
rect 16856 29563 16908 29572
rect 16856 29529 16865 29563
rect 16865 29529 16899 29563
rect 16899 29529 16908 29563
rect 16856 29520 16908 29529
rect 17592 29520 17644 29572
rect 11060 29452 11112 29504
rect 13360 29495 13412 29504
rect 13360 29461 13369 29495
rect 13369 29461 13403 29495
rect 13403 29461 13412 29495
rect 13360 29452 13412 29461
rect 17040 29452 17092 29504
rect 20444 29452 20496 29504
rect 22192 29495 22244 29504
rect 22192 29461 22201 29495
rect 22201 29461 22235 29495
rect 22235 29461 22244 29495
rect 22192 29452 22244 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 5816 29248 5868 29300
rect 6000 29248 6052 29300
rect 9680 29291 9732 29300
rect 9680 29257 9689 29291
rect 9689 29257 9723 29291
rect 9723 29257 9732 29291
rect 9680 29248 9732 29257
rect 11152 29291 11204 29300
rect 11152 29257 11161 29291
rect 11161 29257 11195 29291
rect 11195 29257 11204 29291
rect 11152 29248 11204 29257
rect 14740 29248 14792 29300
rect 15200 29248 15252 29300
rect 6368 29180 6420 29232
rect 6276 29112 6328 29164
rect 6644 29112 6696 29164
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 8944 29112 8996 29164
rect 10048 29155 10100 29164
rect 10048 29121 10082 29155
rect 10082 29121 10100 29155
rect 10048 29112 10100 29121
rect 13360 29180 13412 29232
rect 15108 29180 15160 29232
rect 15200 29155 15252 29164
rect 15200 29121 15209 29155
rect 15209 29121 15243 29155
rect 15243 29121 15252 29155
rect 15200 29112 15252 29121
rect 16488 29180 16540 29232
rect 16856 29248 16908 29300
rect 17500 29248 17552 29300
rect 17592 29248 17644 29300
rect 6552 29044 6604 29096
rect 6460 28976 6512 29028
rect 8024 29087 8076 29096
rect 8024 29053 8033 29087
rect 8033 29053 8067 29087
rect 8067 29053 8076 29087
rect 8024 29044 8076 29053
rect 11060 29044 11112 29096
rect 12348 29087 12400 29096
rect 12348 29053 12357 29087
rect 12357 29053 12391 29087
rect 12391 29053 12400 29087
rect 12348 29044 12400 29053
rect 12624 29087 12676 29096
rect 12624 29053 12633 29087
rect 12633 29053 12667 29087
rect 12667 29053 12676 29087
rect 12624 29044 12676 29053
rect 14556 29044 14608 29096
rect 17040 29155 17092 29164
rect 17040 29121 17049 29155
rect 17049 29121 17083 29155
rect 17083 29121 17092 29155
rect 17040 29112 17092 29121
rect 17132 29155 17184 29164
rect 17132 29121 17141 29155
rect 17141 29121 17175 29155
rect 17175 29121 17184 29155
rect 17132 29112 17184 29121
rect 18052 29180 18104 29232
rect 19984 29248 20036 29300
rect 19524 29180 19576 29232
rect 14188 28976 14240 29028
rect 17500 29044 17552 29096
rect 5540 28908 5592 28960
rect 6644 28908 6696 28960
rect 7288 28951 7340 28960
rect 7288 28917 7297 28951
rect 7297 28917 7331 28951
rect 7331 28917 7340 28951
rect 7288 28908 7340 28917
rect 7472 28951 7524 28960
rect 7472 28917 7481 28951
rect 7481 28917 7515 28951
rect 7515 28917 7524 28951
rect 7472 28908 7524 28917
rect 14280 28951 14332 28960
rect 14280 28917 14289 28951
rect 14289 28917 14323 28951
rect 14323 28917 14332 28951
rect 14280 28908 14332 28917
rect 18144 29044 18196 29096
rect 18512 29044 18564 29096
rect 17960 28908 18012 28960
rect 18236 28908 18288 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 6552 28704 6604 28756
rect 5540 28568 5592 28620
rect 5356 28500 5408 28552
rect 6092 28611 6144 28620
rect 6092 28577 6101 28611
rect 6101 28577 6135 28611
rect 6135 28577 6144 28611
rect 6092 28568 6144 28577
rect 6368 28611 6420 28620
rect 6368 28577 6377 28611
rect 6377 28577 6411 28611
rect 6411 28577 6420 28611
rect 6368 28568 6420 28577
rect 8024 28704 8076 28756
rect 8944 28747 8996 28756
rect 8944 28713 8953 28747
rect 8953 28713 8987 28747
rect 8987 28713 8996 28747
rect 8944 28704 8996 28713
rect 12624 28704 12676 28756
rect 18236 28747 18288 28756
rect 18236 28713 18245 28747
rect 18245 28713 18279 28747
rect 18279 28713 18288 28747
rect 18236 28704 18288 28713
rect 18328 28704 18380 28756
rect 9588 28568 9640 28620
rect 5816 28432 5868 28484
rect 8668 28500 8720 28552
rect 6644 28475 6696 28484
rect 6644 28441 6678 28475
rect 6678 28441 6696 28475
rect 6644 28432 6696 28441
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 12348 28611 12400 28620
rect 12348 28577 12357 28611
rect 12357 28577 12391 28611
rect 12391 28577 12400 28611
rect 12348 28568 12400 28577
rect 13268 28636 13320 28688
rect 18512 28636 18564 28688
rect 16396 28611 16448 28620
rect 16396 28577 16405 28611
rect 16405 28577 16439 28611
rect 16439 28577 16448 28611
rect 16396 28568 16448 28577
rect 16764 28568 16816 28620
rect 18052 28568 18104 28620
rect 10692 28432 10744 28484
rect 9588 28364 9640 28416
rect 12072 28475 12124 28484
rect 12072 28441 12081 28475
rect 12081 28441 12115 28475
rect 12115 28441 12124 28475
rect 12072 28432 12124 28441
rect 13820 28500 13872 28552
rect 14188 28500 14240 28552
rect 14280 28500 14332 28552
rect 16304 28543 16356 28552
rect 16304 28509 16313 28543
rect 16313 28509 16347 28543
rect 16347 28509 16356 28543
rect 16304 28500 16356 28509
rect 17040 28500 17092 28552
rect 17408 28500 17460 28552
rect 17960 28500 18012 28552
rect 19524 28704 19576 28756
rect 13176 28475 13228 28484
rect 13176 28441 13185 28475
rect 13185 28441 13219 28475
rect 13219 28441 13228 28475
rect 13176 28432 13228 28441
rect 14004 28364 14056 28416
rect 18512 28475 18564 28484
rect 18512 28441 18521 28475
rect 18521 28441 18555 28475
rect 18555 28441 18564 28475
rect 18512 28432 18564 28441
rect 18604 28475 18656 28484
rect 18604 28441 18613 28475
rect 18613 28441 18647 28475
rect 18647 28441 18656 28475
rect 18604 28432 18656 28441
rect 19984 28500 20036 28552
rect 20444 28500 20496 28552
rect 21088 28432 21140 28484
rect 19156 28364 19208 28416
rect 19248 28364 19300 28416
rect 20996 28364 21048 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 5816 28160 5868 28212
rect 6460 28160 6512 28212
rect 6644 28160 6696 28212
rect 7288 28160 7340 28212
rect 5540 27820 5592 27872
rect 6920 28092 6972 28144
rect 10784 28160 10836 28212
rect 12072 28160 12124 28212
rect 9588 28092 9640 28144
rect 13728 28160 13780 28212
rect 9220 28067 9272 28076
rect 9220 28033 9229 28067
rect 9229 28033 9263 28067
rect 9263 28033 9272 28067
rect 9220 28024 9272 28033
rect 9404 28067 9456 28076
rect 9404 28033 9413 28067
rect 9413 28033 9447 28067
rect 9447 28033 9456 28067
rect 9404 28024 9456 28033
rect 14004 28160 14056 28212
rect 15200 28160 15252 28212
rect 10232 28067 10284 28076
rect 10232 28033 10241 28067
rect 10241 28033 10275 28067
rect 10275 28033 10284 28067
rect 10232 28024 10284 28033
rect 13084 28067 13136 28076
rect 13084 28033 13093 28067
rect 13093 28033 13127 28067
rect 13127 28033 13136 28067
rect 13084 28024 13136 28033
rect 13360 28024 13412 28076
rect 9680 27956 9732 28008
rect 9772 27999 9824 28008
rect 9772 27965 9781 27999
rect 9781 27965 9815 27999
rect 9815 27965 9824 27999
rect 9772 27956 9824 27965
rect 13268 27956 13320 28008
rect 7472 27820 7524 27872
rect 8484 27863 8536 27872
rect 8484 27829 8493 27863
rect 8493 27829 8527 27863
rect 8527 27829 8536 27863
rect 8484 27820 8536 27829
rect 10140 27863 10192 27872
rect 10140 27829 10149 27863
rect 10149 27829 10183 27863
rect 10183 27829 10192 27863
rect 10140 27820 10192 27829
rect 10416 27863 10468 27872
rect 10416 27829 10425 27863
rect 10425 27829 10459 27863
rect 10459 27829 10468 27863
rect 10416 27820 10468 27829
rect 14372 27820 14424 27872
rect 18604 28160 18656 28212
rect 19156 28203 19208 28212
rect 19156 28169 19165 28203
rect 19165 28169 19199 28203
rect 19199 28169 19208 28203
rect 19156 28160 19208 28169
rect 19248 28160 19300 28212
rect 15752 28067 15804 28076
rect 15752 28033 15761 28067
rect 15761 28033 15795 28067
rect 15795 28033 15804 28067
rect 15752 28024 15804 28033
rect 16396 28092 16448 28144
rect 16488 28135 16540 28144
rect 16488 28101 16497 28135
rect 16497 28101 16531 28135
rect 16531 28101 16540 28135
rect 16488 28092 16540 28101
rect 18512 28135 18564 28144
rect 18512 28101 18521 28135
rect 18521 28101 18555 28135
rect 18555 28101 18564 28135
rect 18512 28092 18564 28101
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 18696 28067 18748 28076
rect 18696 28033 18705 28067
rect 18705 28033 18739 28067
rect 18739 28033 18748 28067
rect 18696 28024 18748 28033
rect 19156 28024 19208 28076
rect 20996 28092 21048 28144
rect 22008 28092 22060 28144
rect 22376 28092 22428 28144
rect 20904 28067 20956 28076
rect 20904 28033 20913 28067
rect 20913 28033 20947 28067
rect 20947 28033 20956 28067
rect 22652 28092 22704 28144
rect 20904 28024 20956 28033
rect 14740 27931 14792 27940
rect 14740 27897 14749 27931
rect 14749 27897 14783 27931
rect 14783 27897 14792 27931
rect 14740 27888 14792 27897
rect 19340 27999 19392 28008
rect 19340 27965 19349 27999
rect 19349 27965 19383 27999
rect 19383 27965 19392 27999
rect 19340 27956 19392 27965
rect 22008 27999 22060 28008
rect 22008 27965 22017 27999
rect 22017 27965 22051 27999
rect 22051 27965 22060 27999
rect 22008 27956 22060 27965
rect 22836 28067 22888 28076
rect 22836 28033 22845 28067
rect 22845 28033 22879 28067
rect 22879 28033 22888 28067
rect 22836 28024 22888 28033
rect 22192 27888 22244 27940
rect 23480 27888 23532 27940
rect 14648 27820 14700 27872
rect 15384 27820 15436 27872
rect 16304 27863 16356 27872
rect 16304 27829 16313 27863
rect 16313 27829 16347 27863
rect 16347 27829 16356 27863
rect 16304 27820 16356 27829
rect 19708 27820 19760 27872
rect 22468 27863 22520 27872
rect 22468 27829 22477 27863
rect 22477 27829 22511 27863
rect 22511 27829 22520 27863
rect 22468 27820 22520 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4068 27616 4120 27668
rect 5540 27616 5592 27668
rect 6460 27616 6512 27668
rect 9404 27616 9456 27668
rect 13176 27616 13228 27668
rect 14740 27616 14792 27668
rect 3792 27455 3844 27464
rect 3792 27421 3801 27455
rect 3801 27421 3835 27455
rect 3835 27421 3844 27455
rect 3792 27412 3844 27421
rect 8484 27480 8536 27532
rect 4160 27344 4212 27396
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 5264 27319 5316 27328
rect 5264 27285 5273 27319
rect 5273 27285 5307 27319
rect 5307 27285 5316 27319
rect 5264 27276 5316 27285
rect 6092 27276 6144 27328
rect 7380 27319 7432 27328
rect 7380 27285 7389 27319
rect 7389 27285 7423 27319
rect 7423 27285 7432 27319
rect 7380 27276 7432 27285
rect 9772 27412 9824 27464
rect 10416 27412 10468 27464
rect 11060 27455 11112 27464
rect 11060 27421 11069 27455
rect 11069 27421 11103 27455
rect 11103 27421 11112 27455
rect 11060 27412 11112 27421
rect 11980 27455 12032 27464
rect 11980 27421 11989 27455
rect 11989 27421 12023 27455
rect 12023 27421 12032 27455
rect 11980 27412 12032 27421
rect 15108 27548 15160 27600
rect 13268 27523 13320 27532
rect 13268 27489 13277 27523
rect 13277 27489 13311 27523
rect 13311 27489 13320 27523
rect 13268 27480 13320 27489
rect 13636 27523 13688 27532
rect 13636 27489 13645 27523
rect 13645 27489 13679 27523
rect 13679 27489 13688 27523
rect 13636 27480 13688 27489
rect 12624 27455 12676 27464
rect 12624 27421 12633 27455
rect 12633 27421 12667 27455
rect 12667 27421 12676 27455
rect 12624 27412 12676 27421
rect 10324 27276 10376 27328
rect 12440 27276 12492 27328
rect 13544 27344 13596 27396
rect 13360 27319 13412 27328
rect 13360 27285 13369 27319
rect 13369 27285 13403 27319
rect 13403 27285 13412 27319
rect 14648 27480 14700 27532
rect 14280 27455 14332 27464
rect 14280 27421 14289 27455
rect 14289 27421 14323 27455
rect 14323 27421 14332 27455
rect 14280 27412 14332 27421
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 14556 27455 14608 27464
rect 14556 27421 14565 27455
rect 14565 27421 14599 27455
rect 14599 27421 14608 27455
rect 14556 27412 14608 27421
rect 15016 27412 15068 27464
rect 13360 27276 13412 27285
rect 13820 27319 13872 27328
rect 13820 27285 13829 27319
rect 13829 27285 13863 27319
rect 13863 27285 13872 27319
rect 13820 27276 13872 27285
rect 15292 27455 15344 27464
rect 15292 27421 15301 27455
rect 15301 27421 15335 27455
rect 15335 27421 15344 27455
rect 15292 27412 15344 27421
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 15660 27455 15712 27464
rect 15660 27421 15669 27455
rect 15669 27421 15703 27455
rect 15703 27421 15712 27455
rect 15660 27412 15712 27421
rect 16580 27455 16632 27464
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 17132 27548 17184 27600
rect 18696 27659 18748 27668
rect 18696 27625 18705 27659
rect 18705 27625 18739 27659
rect 18739 27625 18748 27659
rect 18696 27616 18748 27625
rect 20904 27616 20956 27668
rect 22836 27616 22888 27668
rect 16948 27480 17000 27532
rect 16764 27412 16816 27464
rect 17132 27344 17184 27396
rect 18236 27412 18288 27464
rect 18052 27344 18104 27396
rect 18328 27387 18380 27396
rect 18328 27353 18337 27387
rect 18337 27353 18371 27387
rect 18371 27353 18380 27387
rect 18328 27344 18380 27353
rect 19524 27412 19576 27464
rect 22560 27480 22612 27532
rect 19064 27344 19116 27396
rect 19984 27412 20036 27464
rect 20536 27387 20588 27396
rect 20536 27353 20545 27387
rect 20545 27353 20579 27387
rect 20579 27353 20588 27387
rect 20536 27344 20588 27353
rect 21272 27344 21324 27396
rect 19156 27276 19208 27328
rect 19800 27276 19852 27328
rect 22008 27319 22060 27328
rect 22008 27285 22017 27319
rect 22017 27285 22051 27319
rect 22051 27285 22060 27319
rect 22008 27276 22060 27285
rect 23480 27412 23532 27464
rect 23940 27412 23992 27464
rect 22744 27276 22796 27328
rect 22836 27276 22888 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 4160 27115 4212 27124
rect 4160 27081 4169 27115
rect 4169 27081 4203 27115
rect 4203 27081 4212 27115
rect 4160 27072 4212 27081
rect 5264 27072 5316 27124
rect 5540 27072 5592 27124
rect 7380 27072 7432 27124
rect 10232 27072 10284 27124
rect 12624 27072 12676 27124
rect 13084 27072 13136 27124
rect 13544 27072 13596 27124
rect 13728 27072 13780 27124
rect 13820 27072 13872 27124
rect 14280 27072 14332 27124
rect 15660 27072 15712 27124
rect 17040 27115 17092 27124
rect 6092 26936 6144 26988
rect 3332 26911 3384 26920
rect 3332 26877 3341 26911
rect 3341 26877 3375 26911
rect 3375 26877 3384 26911
rect 3332 26868 3384 26877
rect 8208 26979 8260 26988
rect 8208 26945 8217 26979
rect 8217 26945 8251 26979
rect 8251 26945 8260 26979
rect 8208 26936 8260 26945
rect 11060 27004 11112 27056
rect 7840 26911 7892 26920
rect 7840 26877 7849 26911
rect 7849 26877 7883 26911
rect 7883 26877 7892 26911
rect 7840 26868 7892 26877
rect 10140 26936 10192 26988
rect 10784 26979 10836 26988
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 5632 26800 5684 26852
rect 9772 26843 9824 26852
rect 9772 26809 9781 26843
rect 9781 26809 9815 26843
rect 9815 26809 9824 26843
rect 9772 26800 9824 26809
rect 4620 26732 4672 26784
rect 5540 26775 5592 26784
rect 5540 26741 5549 26775
rect 5549 26741 5583 26775
rect 5583 26741 5592 26775
rect 5540 26732 5592 26741
rect 7196 26775 7248 26784
rect 7196 26741 7205 26775
rect 7205 26741 7239 26775
rect 7239 26741 7248 26775
rect 7196 26732 7248 26741
rect 9496 26732 9548 26784
rect 10324 26868 10376 26920
rect 10968 26868 11020 26920
rect 10508 26800 10560 26852
rect 11888 26936 11940 26988
rect 12532 26936 12584 26988
rect 13268 26936 13320 26988
rect 12440 26800 12492 26852
rect 13176 26868 13228 26920
rect 13912 26911 13964 26920
rect 13912 26877 13921 26911
rect 13921 26877 13955 26911
rect 13955 26877 13964 26911
rect 13912 26868 13964 26877
rect 12532 26732 12584 26784
rect 17040 27081 17049 27115
rect 17049 27081 17083 27115
rect 17083 27081 17092 27115
rect 17040 27072 17092 27081
rect 16304 27004 16356 27056
rect 14464 26936 14516 26988
rect 14740 26868 14792 26920
rect 15200 26979 15252 26988
rect 15200 26945 15209 26979
rect 15209 26945 15243 26979
rect 15243 26945 15252 26979
rect 15200 26936 15252 26945
rect 15384 26979 15436 26988
rect 15384 26945 15393 26979
rect 15393 26945 15427 26979
rect 15427 26945 15436 26979
rect 15384 26936 15436 26945
rect 15568 26936 15620 26988
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 17316 27004 17368 27056
rect 18328 27115 18380 27124
rect 18328 27081 18337 27115
rect 18337 27081 18371 27115
rect 18371 27081 18380 27115
rect 18328 27072 18380 27081
rect 18420 27115 18472 27124
rect 18420 27081 18429 27115
rect 18429 27081 18463 27115
rect 18463 27081 18472 27115
rect 18420 27072 18472 27081
rect 19524 27072 19576 27124
rect 20536 27072 20588 27124
rect 21272 27072 21324 27124
rect 22468 27072 22520 27124
rect 22652 27115 22704 27124
rect 22652 27081 22661 27115
rect 22661 27081 22695 27115
rect 22695 27081 22704 27115
rect 22652 27072 22704 27081
rect 23940 27072 23992 27124
rect 18696 27047 18748 27056
rect 18696 27013 18705 27047
rect 18705 27013 18739 27047
rect 18739 27013 18748 27047
rect 18696 27004 18748 27013
rect 18788 27047 18840 27056
rect 18788 27013 18797 27047
rect 18797 27013 18831 27047
rect 18831 27013 18840 27047
rect 18788 27004 18840 27013
rect 16948 26936 17000 26988
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 17408 26936 17460 26945
rect 17684 26979 17736 26988
rect 17684 26945 17693 26979
rect 17693 26945 17727 26979
rect 17727 26945 17736 26979
rect 17684 26936 17736 26945
rect 17776 26936 17828 26988
rect 18052 26936 18104 26988
rect 16948 26800 17000 26852
rect 18420 26868 18472 26920
rect 17500 26843 17552 26852
rect 17500 26809 17509 26843
rect 17509 26809 17543 26843
rect 17543 26809 17552 26843
rect 17500 26800 17552 26809
rect 20720 27004 20772 27056
rect 21088 27004 21140 27056
rect 19800 26800 19852 26852
rect 20352 26800 20404 26852
rect 20996 26868 21048 26920
rect 21180 26868 21232 26920
rect 22008 26936 22060 26988
rect 21732 26868 21784 26920
rect 22836 26979 22888 26988
rect 22836 26945 22845 26979
rect 22845 26945 22879 26979
rect 22879 26945 22888 26979
rect 22836 26936 22888 26945
rect 17316 26732 17368 26784
rect 19156 26732 19208 26784
rect 19708 26732 19760 26784
rect 22744 26732 22796 26784
rect 23388 26732 23440 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3332 26528 3384 26580
rect 6092 26528 6144 26580
rect 8208 26528 8260 26580
rect 9220 26528 9272 26580
rect 9496 26528 9548 26580
rect 9772 26528 9824 26580
rect 11060 26528 11112 26580
rect 15200 26571 15252 26580
rect 15200 26537 15209 26571
rect 15209 26537 15243 26571
rect 15243 26537 15252 26571
rect 15200 26528 15252 26537
rect 16580 26528 16632 26580
rect 18052 26528 18104 26580
rect 19708 26528 19760 26580
rect 3792 26392 3844 26444
rect 4436 26367 4488 26376
rect 4436 26333 4445 26367
rect 4445 26333 4479 26367
rect 4479 26333 4488 26367
rect 4436 26324 4488 26333
rect 6368 26392 6420 26444
rect 7196 26324 7248 26376
rect 8484 26324 8536 26376
rect 9680 26392 9732 26444
rect 10416 26392 10468 26444
rect 18696 26460 18748 26512
rect 3608 26256 3660 26308
rect 3884 26231 3936 26240
rect 3884 26197 3893 26231
rect 3893 26197 3927 26231
rect 3927 26197 3936 26231
rect 3884 26188 3936 26197
rect 4804 26188 4856 26240
rect 8392 26256 8444 26308
rect 9864 26324 9916 26376
rect 10968 26324 11020 26376
rect 11980 26324 12032 26376
rect 13728 26324 13780 26376
rect 15016 26324 15068 26376
rect 15660 26324 15712 26376
rect 15752 26324 15804 26376
rect 16856 26392 16908 26444
rect 22284 26460 22336 26512
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 17500 26324 17552 26376
rect 22744 26392 22796 26444
rect 11152 26256 11204 26308
rect 16580 26299 16632 26308
rect 16580 26265 16589 26299
rect 16589 26265 16623 26299
rect 16623 26265 16632 26299
rect 16580 26256 16632 26265
rect 20168 26299 20220 26308
rect 15568 26188 15620 26240
rect 20168 26265 20177 26299
rect 20177 26265 20211 26299
rect 20211 26265 20220 26299
rect 20168 26256 20220 26265
rect 20352 26299 20404 26308
rect 20352 26265 20361 26299
rect 20361 26265 20395 26299
rect 20395 26265 20404 26299
rect 20352 26256 20404 26265
rect 22100 26256 22152 26308
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23296 26324 23348 26333
rect 17776 26188 17828 26240
rect 20996 26188 21048 26240
rect 22008 26188 22060 26240
rect 22376 26231 22428 26240
rect 22376 26197 22385 26231
rect 22385 26197 22419 26231
rect 22419 26197 22428 26231
rect 22376 26188 22428 26197
rect 22928 26188 22980 26240
rect 23388 26188 23440 26240
rect 28908 26256 28960 26308
rect 23572 26231 23624 26240
rect 23572 26197 23581 26231
rect 23581 26197 23615 26231
rect 23615 26197 23624 26231
rect 23572 26188 23624 26197
rect 26976 26188 27028 26240
rect 28264 26188 28316 26240
rect 29184 26231 29236 26240
rect 29184 26197 29193 26231
rect 29193 26197 29227 26231
rect 29227 26197 29236 26231
rect 29184 26188 29236 26197
rect 30564 26188 30616 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 4436 25984 4488 26036
rect 4620 25984 4672 26036
rect 4804 25984 4856 26036
rect 5540 25984 5592 26036
rect 9680 25984 9732 26036
rect 9864 25984 9916 26036
rect 10692 25984 10744 26036
rect 11244 26027 11296 26036
rect 11244 25993 11253 26027
rect 11253 25993 11287 26027
rect 11287 25993 11296 26027
rect 11244 25984 11296 25993
rect 13636 25984 13688 26036
rect 13728 25984 13780 26036
rect 13912 25984 13964 26036
rect 16856 26027 16908 26036
rect 16856 25993 16865 26027
rect 16865 25993 16899 26027
rect 16899 25993 16908 26027
rect 16856 25984 16908 25993
rect 2780 25891 2832 25900
rect 2780 25857 2798 25891
rect 2798 25857 2832 25891
rect 2780 25848 2832 25857
rect 3516 25891 3568 25900
rect 3516 25857 3525 25891
rect 3525 25857 3559 25891
rect 3559 25857 3568 25891
rect 3516 25848 3568 25857
rect 3792 25848 3844 25900
rect 4068 25823 4120 25832
rect 4068 25789 4077 25823
rect 4077 25789 4111 25823
rect 4111 25789 4120 25823
rect 4068 25780 4120 25789
rect 1676 25687 1728 25696
rect 1676 25653 1685 25687
rect 1685 25653 1719 25687
rect 1719 25653 1728 25687
rect 5632 25848 5684 25900
rect 7840 25848 7892 25900
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 6920 25712 6972 25764
rect 8208 25712 8260 25764
rect 11612 25848 11664 25900
rect 12440 25848 12492 25900
rect 12532 25848 12584 25900
rect 13452 25891 13504 25900
rect 13452 25857 13461 25891
rect 13461 25857 13495 25891
rect 13495 25857 13504 25891
rect 13452 25848 13504 25857
rect 18420 26027 18472 26036
rect 18420 25993 18429 26027
rect 18429 25993 18463 26027
rect 18463 25993 18472 26027
rect 18420 25984 18472 25993
rect 19340 25984 19392 26036
rect 20076 25984 20128 26036
rect 12256 25780 12308 25832
rect 13360 25780 13412 25832
rect 1676 25644 1728 25653
rect 3148 25644 3200 25696
rect 3700 25644 3752 25696
rect 5264 25644 5316 25696
rect 9404 25687 9456 25696
rect 9404 25653 9413 25687
rect 9413 25653 9447 25687
rect 9447 25653 9456 25687
rect 9404 25644 9456 25653
rect 10048 25644 10100 25696
rect 11520 25644 11572 25696
rect 11888 25644 11940 25696
rect 12624 25644 12676 25696
rect 15016 25644 15068 25696
rect 16764 25848 16816 25900
rect 20812 25916 20864 25968
rect 21180 25916 21232 25968
rect 22376 25984 22428 26036
rect 23296 25984 23348 26036
rect 18236 25848 18288 25900
rect 18420 25848 18472 25900
rect 19248 25848 19300 25900
rect 20168 25848 20220 25900
rect 20720 25891 20772 25900
rect 20720 25857 20729 25891
rect 20729 25857 20763 25891
rect 20763 25857 20772 25891
rect 20720 25848 20772 25857
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 21272 25891 21324 25900
rect 21272 25857 21281 25891
rect 21281 25857 21315 25891
rect 21315 25857 21324 25891
rect 21272 25848 21324 25857
rect 21456 25891 21508 25900
rect 21456 25857 21465 25891
rect 21465 25857 21499 25891
rect 21499 25857 21508 25891
rect 21456 25848 21508 25857
rect 22284 25848 22336 25900
rect 19156 25780 19208 25832
rect 23388 25916 23440 25968
rect 23572 25916 23624 25968
rect 30380 25984 30432 26036
rect 30564 25984 30616 26036
rect 35440 25984 35492 26036
rect 22560 25848 22612 25900
rect 23940 25848 23992 25900
rect 28356 25848 28408 25900
rect 29184 25848 29236 25900
rect 30472 25916 30524 25968
rect 25136 25780 25188 25832
rect 17316 25712 17368 25764
rect 16580 25644 16632 25696
rect 17500 25644 17552 25696
rect 17592 25687 17644 25696
rect 17592 25653 17601 25687
rect 17601 25653 17635 25687
rect 17635 25653 17644 25687
rect 17592 25644 17644 25653
rect 19432 25644 19484 25696
rect 19984 25687 20036 25696
rect 19984 25653 19993 25687
rect 19993 25653 20027 25687
rect 20027 25653 20036 25687
rect 19984 25644 20036 25653
rect 21916 25644 21968 25696
rect 22100 25644 22152 25696
rect 22376 25687 22428 25696
rect 22376 25653 22385 25687
rect 22385 25653 22419 25687
rect 22419 25653 22428 25687
rect 22376 25644 22428 25653
rect 28264 25644 28316 25696
rect 29736 25823 29788 25832
rect 29736 25789 29745 25823
rect 29745 25789 29779 25823
rect 29779 25789 29788 25823
rect 29736 25780 29788 25789
rect 33324 25780 33376 25832
rect 31208 25687 31260 25696
rect 31208 25653 31217 25687
rect 31217 25653 31251 25687
rect 31251 25653 31260 25687
rect 31208 25644 31260 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2780 25440 2832 25492
rect 3332 25440 3384 25492
rect 3516 25483 3568 25492
rect 3516 25449 3525 25483
rect 3525 25449 3559 25483
rect 3559 25449 3568 25483
rect 3516 25440 3568 25449
rect 3608 25440 3660 25492
rect 8668 25440 8720 25492
rect 3148 25415 3200 25424
rect 3148 25381 3157 25415
rect 3157 25381 3191 25415
rect 3191 25381 3200 25415
rect 3148 25372 3200 25381
rect 9864 25440 9916 25492
rect 10968 25440 11020 25492
rect 12624 25440 12676 25492
rect 13452 25440 13504 25492
rect 15016 25440 15068 25492
rect 15384 25440 15436 25492
rect 3240 25347 3292 25356
rect 3240 25313 3249 25347
rect 3249 25313 3283 25347
rect 3283 25313 3292 25347
rect 3240 25304 3292 25313
rect 940 25100 992 25152
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 4068 25304 4120 25356
rect 3884 25236 3936 25288
rect 5264 25279 5316 25288
rect 5264 25245 5273 25279
rect 5273 25245 5307 25279
rect 5307 25245 5316 25279
rect 5264 25236 5316 25245
rect 5448 25279 5500 25288
rect 5448 25245 5457 25279
rect 5457 25245 5491 25279
rect 5491 25245 5500 25279
rect 5448 25236 5500 25245
rect 5540 25279 5592 25288
rect 5540 25245 5549 25279
rect 5549 25245 5583 25279
rect 5583 25245 5592 25279
rect 5540 25236 5592 25245
rect 11612 25372 11664 25424
rect 8024 25304 8076 25356
rect 12716 25304 12768 25356
rect 9956 25236 10008 25288
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 11244 25236 11296 25288
rect 12256 25236 12308 25288
rect 2872 25211 2924 25220
rect 2872 25177 2881 25211
rect 2881 25177 2915 25211
rect 2915 25177 2924 25211
rect 2872 25168 2924 25177
rect 4804 25100 4856 25152
rect 7840 25168 7892 25220
rect 9404 25211 9456 25220
rect 9404 25177 9438 25211
rect 9438 25177 9456 25211
rect 9404 25168 9456 25177
rect 12440 25168 12492 25220
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 11336 25143 11388 25152
rect 11336 25109 11345 25143
rect 11345 25109 11379 25143
rect 11379 25109 11388 25143
rect 11336 25100 11388 25109
rect 11428 25100 11480 25152
rect 12716 25100 12768 25152
rect 14832 25168 14884 25220
rect 15292 25236 15344 25288
rect 15752 25236 15804 25288
rect 16764 25483 16816 25492
rect 16764 25449 16773 25483
rect 16773 25449 16807 25483
rect 16807 25449 16816 25483
rect 16764 25440 16816 25449
rect 17316 25483 17368 25492
rect 17316 25449 17325 25483
rect 17325 25449 17359 25483
rect 17359 25449 17368 25483
rect 17316 25440 17368 25449
rect 17500 25483 17552 25492
rect 17500 25449 17509 25483
rect 17509 25449 17543 25483
rect 17543 25449 17552 25483
rect 17500 25440 17552 25449
rect 17592 25440 17644 25492
rect 20720 25440 20772 25492
rect 20904 25483 20956 25492
rect 20904 25449 20913 25483
rect 20913 25449 20947 25483
rect 20947 25449 20956 25483
rect 20904 25440 20956 25449
rect 22100 25440 22152 25492
rect 15384 25211 15436 25220
rect 15384 25177 15393 25211
rect 15393 25177 15427 25211
rect 15427 25177 15436 25211
rect 15384 25168 15436 25177
rect 16304 25236 16356 25288
rect 17040 25304 17092 25356
rect 20628 25372 20680 25424
rect 20076 25236 20128 25288
rect 20260 25279 20312 25288
rect 20260 25245 20269 25279
rect 20269 25245 20303 25279
rect 20303 25245 20312 25279
rect 20260 25236 20312 25245
rect 21180 25279 21232 25288
rect 21180 25245 21189 25279
rect 21189 25245 21223 25279
rect 21223 25245 21232 25279
rect 21180 25236 21232 25245
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 22376 25440 22428 25492
rect 22560 25483 22612 25492
rect 22560 25449 22569 25483
rect 22569 25449 22603 25483
rect 22603 25449 22612 25483
rect 22560 25440 22612 25449
rect 23388 25483 23440 25492
rect 23388 25449 23397 25483
rect 23397 25449 23431 25483
rect 23431 25449 23440 25483
rect 23388 25440 23440 25449
rect 29736 25483 29788 25492
rect 29736 25449 29745 25483
rect 29745 25449 29779 25483
rect 29779 25449 29788 25483
rect 29736 25440 29788 25449
rect 30472 25440 30524 25492
rect 28080 25372 28132 25424
rect 35440 25372 35492 25424
rect 22744 25279 22796 25288
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 22928 25279 22980 25288
rect 22928 25245 22937 25279
rect 22937 25245 22971 25279
rect 22971 25245 22980 25279
rect 22928 25236 22980 25245
rect 23296 25236 23348 25288
rect 25136 25236 25188 25288
rect 26976 25236 27028 25288
rect 17132 25100 17184 25152
rect 19064 25100 19116 25152
rect 25688 25211 25740 25220
rect 25688 25177 25697 25211
rect 25697 25177 25731 25211
rect 25731 25177 25740 25211
rect 25688 25168 25740 25177
rect 26424 25168 26476 25220
rect 29552 25279 29604 25288
rect 29552 25245 29561 25279
rect 29561 25245 29595 25279
rect 29595 25245 29604 25279
rect 29552 25236 29604 25245
rect 20168 25100 20220 25152
rect 20352 25100 20404 25152
rect 27160 25143 27212 25152
rect 27160 25109 27169 25143
rect 27169 25109 27203 25143
rect 27203 25109 27212 25143
rect 27160 25100 27212 25109
rect 30656 25100 30708 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 1952 24939 2004 24948
rect 1952 24905 1961 24939
rect 1961 24905 1995 24939
rect 1995 24905 2004 24939
rect 1952 24896 2004 24905
rect 2136 24828 2188 24880
rect 3700 24896 3752 24948
rect 5540 24896 5592 24948
rect 1676 24760 1728 24812
rect 3240 24828 3292 24880
rect 4804 24828 4856 24880
rect 10784 24939 10836 24948
rect 10784 24905 10793 24939
rect 10793 24905 10827 24939
rect 10827 24905 10836 24939
rect 10784 24896 10836 24905
rect 11336 24896 11388 24948
rect 11428 24896 11480 24948
rect 13820 24896 13872 24948
rect 2872 24760 2924 24812
rect 3332 24760 3384 24812
rect 3792 24760 3844 24812
rect 3884 24692 3936 24744
rect 5540 24692 5592 24744
rect 6184 24760 6236 24812
rect 11152 24828 11204 24880
rect 8208 24760 8260 24812
rect 8300 24803 8352 24812
rect 8300 24769 8309 24803
rect 8309 24769 8343 24803
rect 8343 24769 8352 24803
rect 8300 24760 8352 24769
rect 10692 24760 10744 24812
rect 10876 24760 10928 24812
rect 11520 24803 11572 24812
rect 11520 24769 11529 24803
rect 11529 24769 11563 24803
rect 11563 24769 11572 24803
rect 11520 24760 11572 24769
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 13636 24871 13688 24880
rect 13636 24837 13645 24871
rect 13645 24837 13679 24871
rect 13679 24837 13688 24871
rect 13636 24828 13688 24837
rect 13360 24760 13412 24812
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 13820 24760 13872 24812
rect 13912 24803 13964 24812
rect 13912 24769 13921 24803
rect 13921 24769 13955 24803
rect 13955 24769 13964 24803
rect 13912 24760 13964 24769
rect 1124 24556 1176 24608
rect 3700 24599 3752 24608
rect 3700 24565 3709 24599
rect 3709 24565 3743 24599
rect 3743 24565 3752 24599
rect 3700 24556 3752 24565
rect 5540 24556 5592 24608
rect 6828 24624 6880 24676
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 14464 24896 14516 24948
rect 15384 24896 15436 24948
rect 15752 24896 15804 24948
rect 19064 24896 19116 24948
rect 20168 24939 20220 24948
rect 20168 24905 20177 24939
rect 20177 24905 20211 24939
rect 20211 24905 20220 24939
rect 20168 24896 20220 24905
rect 22560 24896 22612 24948
rect 25688 24896 25740 24948
rect 26424 24939 26476 24948
rect 26424 24905 26433 24939
rect 26433 24905 26467 24939
rect 26467 24905 26476 24939
rect 26424 24896 26476 24905
rect 27528 24896 27580 24948
rect 28448 24896 28500 24948
rect 29552 24896 29604 24948
rect 31208 24896 31260 24948
rect 14556 24803 14608 24812
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 15108 24760 15160 24812
rect 17040 24871 17092 24880
rect 17040 24837 17049 24871
rect 17049 24837 17083 24871
rect 17083 24837 17092 24871
rect 17040 24828 17092 24837
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 16764 24803 16816 24812
rect 16764 24769 16773 24803
rect 16773 24769 16807 24803
rect 16807 24769 16816 24803
rect 16764 24760 16816 24769
rect 18880 24803 18932 24812
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 20260 24803 20312 24812
rect 20260 24769 20269 24803
rect 20269 24769 20303 24803
rect 20303 24769 20312 24803
rect 20260 24760 20312 24769
rect 20720 24760 20772 24812
rect 21180 24760 21232 24812
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 21456 24828 21508 24880
rect 22284 24828 22336 24880
rect 22100 24692 22152 24744
rect 23388 24760 23440 24812
rect 26148 24803 26200 24812
rect 26148 24769 26157 24803
rect 26157 24769 26191 24803
rect 26191 24769 26200 24803
rect 26148 24760 26200 24769
rect 28080 24760 28132 24812
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 30564 24828 30616 24880
rect 7380 24556 7432 24608
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 10968 24556 11020 24565
rect 11060 24556 11112 24608
rect 11244 24556 11296 24608
rect 13544 24556 13596 24608
rect 19248 24624 19300 24676
rect 15476 24556 15528 24608
rect 17224 24556 17276 24608
rect 19616 24556 19668 24608
rect 21456 24556 21508 24608
rect 21548 24599 21600 24608
rect 21548 24565 21557 24599
rect 21557 24565 21591 24599
rect 21591 24565 21600 24599
rect 21548 24556 21600 24565
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 22008 24556 22060 24608
rect 27160 24624 27212 24676
rect 24308 24556 24360 24608
rect 25136 24556 25188 24608
rect 25228 24599 25280 24608
rect 25228 24565 25237 24599
rect 25237 24565 25271 24599
rect 25271 24565 25280 24599
rect 25228 24556 25280 24565
rect 25412 24556 25464 24608
rect 28908 24760 28960 24812
rect 30472 24760 30524 24812
rect 28448 24599 28500 24608
rect 28448 24565 28457 24599
rect 28457 24565 28491 24599
rect 28491 24565 28500 24599
rect 28448 24556 28500 24565
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 29000 24624 29052 24676
rect 30656 24692 30708 24744
rect 32220 24828 32272 24880
rect 30656 24556 30708 24608
rect 31116 24556 31168 24608
rect 31668 24599 31720 24608
rect 31668 24565 31677 24599
rect 31677 24565 31711 24599
rect 31711 24565 31720 24599
rect 31668 24556 31720 24565
rect 33140 24692 33192 24744
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3240 24352 3292 24404
rect 5448 24352 5500 24404
rect 4804 24284 4856 24336
rect 6184 24352 6236 24404
rect 3792 24259 3844 24268
rect 3792 24225 3801 24259
rect 3801 24225 3835 24259
rect 3835 24225 3844 24259
rect 3792 24216 3844 24225
rect 7380 24352 7432 24404
rect 10048 24352 10100 24404
rect 18880 24352 18932 24404
rect 13912 24284 13964 24336
rect 3240 24148 3292 24200
rect 3332 24191 3384 24200
rect 3332 24157 3341 24191
rect 3341 24157 3375 24191
rect 3375 24157 3384 24191
rect 3332 24148 3384 24157
rect 2044 24080 2096 24132
rect 3240 24055 3292 24064
rect 3240 24021 3249 24055
rect 3249 24021 3283 24055
rect 3283 24021 3292 24055
rect 3240 24012 3292 24021
rect 3700 24148 3752 24200
rect 5356 24148 5408 24200
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 4160 24012 4212 24064
rect 4712 24012 4764 24064
rect 5448 24012 5500 24064
rect 8300 24216 8352 24268
rect 9956 24216 10008 24268
rect 13544 24259 13596 24268
rect 13544 24225 13553 24259
rect 13553 24225 13587 24259
rect 13587 24225 13596 24259
rect 13544 24216 13596 24225
rect 11060 24191 11112 24200
rect 11060 24157 11069 24191
rect 11069 24157 11103 24191
rect 11103 24157 11112 24191
rect 11060 24148 11112 24157
rect 7656 24080 7708 24132
rect 11244 24080 11296 24132
rect 11612 24080 11664 24132
rect 12348 24080 12400 24132
rect 17960 24216 18012 24268
rect 21824 24352 21876 24404
rect 17316 24191 17368 24200
rect 17316 24157 17325 24191
rect 17325 24157 17359 24191
rect 17359 24157 17368 24191
rect 17316 24148 17368 24157
rect 21916 24148 21968 24200
rect 23388 24352 23440 24404
rect 26148 24352 26200 24404
rect 25136 24216 25188 24268
rect 26976 24216 27028 24268
rect 27160 24352 27212 24404
rect 29000 24352 29052 24404
rect 33600 24395 33652 24404
rect 33600 24361 33609 24395
rect 33609 24361 33643 24395
rect 33643 24361 33652 24395
rect 33600 24352 33652 24361
rect 35348 24352 35400 24404
rect 27252 24259 27304 24268
rect 27252 24225 27261 24259
rect 27261 24225 27295 24259
rect 27295 24225 27304 24259
rect 27252 24216 27304 24225
rect 28816 24216 28868 24268
rect 24308 24148 24360 24200
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 28080 24191 28132 24200
rect 28080 24157 28089 24191
rect 28089 24157 28123 24191
rect 28123 24157 28132 24191
rect 28080 24148 28132 24157
rect 28908 24148 28960 24200
rect 29460 24216 29512 24268
rect 30380 24216 30432 24268
rect 31116 24216 31168 24268
rect 18880 24080 18932 24132
rect 23020 24080 23072 24132
rect 24676 24123 24728 24132
rect 24676 24089 24685 24123
rect 24685 24089 24719 24123
rect 24719 24089 24728 24123
rect 24676 24080 24728 24089
rect 25412 24080 25464 24132
rect 28172 24080 28224 24132
rect 6828 24012 6880 24064
rect 8576 24055 8628 24064
rect 8576 24021 8585 24055
rect 8585 24021 8619 24055
rect 8619 24021 8628 24055
rect 8576 24012 8628 24021
rect 9680 24012 9732 24064
rect 10968 24012 11020 24064
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 13176 24012 13228 24064
rect 13268 24055 13320 24064
rect 13268 24021 13277 24055
rect 13277 24021 13311 24055
rect 13311 24021 13320 24055
rect 13268 24012 13320 24021
rect 14832 24012 14884 24064
rect 19156 24012 19208 24064
rect 20076 24012 20128 24064
rect 22376 24012 22428 24064
rect 26056 24012 26108 24064
rect 27988 24055 28040 24064
rect 27988 24021 27997 24055
rect 27997 24021 28031 24055
rect 28031 24021 28040 24055
rect 30472 24148 30524 24200
rect 32588 24191 32640 24200
rect 32588 24157 32597 24191
rect 32597 24157 32631 24191
rect 32631 24157 32640 24191
rect 32588 24148 32640 24157
rect 27988 24012 28040 24021
rect 28356 24055 28408 24064
rect 28356 24021 28365 24055
rect 28365 24021 28399 24055
rect 28399 24021 28408 24055
rect 31668 24080 31720 24132
rect 28356 24012 28408 24021
rect 28632 24012 28684 24064
rect 28908 24055 28960 24064
rect 28908 24021 28917 24055
rect 28917 24021 28951 24055
rect 28951 24021 28960 24055
rect 28908 24012 28960 24021
rect 30288 24055 30340 24064
rect 30288 24021 30297 24055
rect 30297 24021 30331 24055
rect 30331 24021 30340 24055
rect 30288 24012 30340 24021
rect 30472 24012 30524 24064
rect 30656 24012 30708 24064
rect 33140 24012 33192 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 2044 23851 2096 23860
rect 2044 23817 2053 23851
rect 2053 23817 2087 23851
rect 2087 23817 2096 23851
rect 2044 23808 2096 23817
rect 2136 23808 2188 23860
rect 3240 23808 3292 23860
rect 3884 23851 3936 23860
rect 3884 23817 3893 23851
rect 3893 23817 3927 23851
rect 3927 23817 3936 23851
rect 3884 23808 3936 23817
rect 4068 23808 4120 23860
rect 5356 23808 5408 23860
rect 5448 23808 5500 23860
rect 7656 23851 7708 23860
rect 7656 23817 7665 23851
rect 7665 23817 7699 23851
rect 7699 23817 7708 23851
rect 7656 23808 7708 23817
rect 6828 23740 6880 23792
rect 4712 23647 4764 23656
rect 4712 23613 4721 23647
rect 4721 23613 4755 23647
rect 4755 23613 4764 23647
rect 4712 23604 4764 23613
rect 4804 23579 4856 23588
rect 4804 23545 4813 23579
rect 4813 23545 4847 23579
rect 4847 23545 4856 23579
rect 4804 23536 4856 23545
rect 7840 23715 7892 23724
rect 7840 23681 7849 23715
rect 7849 23681 7883 23715
rect 7883 23681 7892 23715
rect 7840 23672 7892 23681
rect 8024 23672 8076 23724
rect 9220 23672 9272 23724
rect 8576 23604 8628 23656
rect 9036 23604 9088 23656
rect 10692 23740 10744 23792
rect 11612 23851 11664 23860
rect 11612 23817 11621 23851
rect 11621 23817 11655 23851
rect 11655 23817 11664 23851
rect 11612 23808 11664 23817
rect 11704 23808 11756 23860
rect 12348 23851 12400 23860
rect 12348 23817 12357 23851
rect 12357 23817 12391 23851
rect 12391 23817 12400 23851
rect 12348 23808 12400 23817
rect 12900 23808 12952 23860
rect 13268 23808 13320 23860
rect 13912 23808 13964 23860
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 9680 23672 9732 23724
rect 10876 23672 10928 23724
rect 12532 23672 12584 23724
rect 15200 23672 15252 23724
rect 17132 23851 17184 23860
rect 17132 23817 17141 23851
rect 17141 23817 17175 23851
rect 17175 23817 17184 23851
rect 17132 23808 17184 23817
rect 19156 23808 19208 23860
rect 21548 23808 21600 23860
rect 23756 23808 23808 23860
rect 24676 23851 24728 23860
rect 24676 23817 24685 23851
rect 24685 23817 24719 23851
rect 24719 23817 24728 23851
rect 24676 23808 24728 23817
rect 18880 23740 18932 23792
rect 18972 23740 19024 23792
rect 9496 23536 9548 23588
rect 9588 23579 9640 23588
rect 9588 23545 9597 23579
rect 9597 23545 9631 23579
rect 9631 23545 9640 23579
rect 9588 23536 9640 23545
rect 9864 23536 9916 23588
rect 14832 23647 14884 23656
rect 14832 23613 14841 23647
rect 14841 23613 14875 23647
rect 14875 23613 14884 23647
rect 14832 23604 14884 23613
rect 14740 23536 14792 23588
rect 15016 23536 15068 23588
rect 16764 23536 16816 23588
rect 18420 23604 18472 23656
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 20076 23604 20128 23656
rect 22376 23604 22428 23656
rect 22652 23672 22704 23724
rect 28816 23808 28868 23860
rect 28908 23808 28960 23860
rect 30288 23808 30340 23860
rect 32588 23808 32640 23860
rect 25136 23672 25188 23724
rect 26424 23715 26476 23724
rect 26424 23681 26433 23715
rect 26433 23681 26467 23715
rect 26467 23681 26476 23715
rect 26424 23672 26476 23681
rect 28080 23672 28132 23724
rect 26056 23604 26108 23656
rect 27252 23604 27304 23656
rect 25872 23536 25924 23588
rect 13912 23511 13964 23520
rect 13912 23477 13921 23511
rect 13921 23477 13955 23511
rect 13955 23477 13964 23511
rect 13912 23468 13964 23477
rect 15752 23468 15804 23520
rect 18236 23511 18288 23520
rect 18236 23477 18245 23511
rect 18245 23477 18279 23511
rect 18279 23477 18288 23511
rect 18236 23468 18288 23477
rect 19064 23468 19116 23520
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 20628 23468 20680 23520
rect 24584 23511 24636 23520
rect 24584 23477 24593 23511
rect 24593 23477 24627 23511
rect 24627 23477 24636 23511
rect 24584 23468 24636 23477
rect 26148 23468 26200 23520
rect 27988 23536 28040 23588
rect 33140 23740 33192 23792
rect 32588 23536 32640 23588
rect 33600 23715 33652 23724
rect 33600 23681 33609 23715
rect 33609 23681 33643 23715
rect 33643 23681 33652 23715
rect 33600 23672 33652 23681
rect 33692 23672 33744 23724
rect 28816 23511 28868 23520
rect 28816 23477 28825 23511
rect 28825 23477 28859 23511
rect 28859 23477 28868 23511
rect 28816 23468 28868 23477
rect 30656 23511 30708 23520
rect 30656 23477 30665 23511
rect 30665 23477 30699 23511
rect 30699 23477 30708 23511
rect 30656 23468 30708 23477
rect 30840 23511 30892 23520
rect 30840 23477 30849 23511
rect 30849 23477 30883 23511
rect 30883 23477 30892 23511
rect 30840 23468 30892 23477
rect 32864 23511 32916 23520
rect 32864 23477 32873 23511
rect 32873 23477 32907 23511
rect 32907 23477 32916 23511
rect 32864 23468 32916 23477
rect 33876 23468 33928 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8024 23264 8076 23316
rect 9588 23264 9640 23316
rect 9680 23264 9732 23316
rect 16764 23264 16816 23316
rect 17960 23264 18012 23316
rect 21180 23307 21232 23316
rect 21180 23273 21189 23307
rect 21189 23273 21223 23307
rect 21223 23273 21232 23307
rect 21180 23264 21232 23273
rect 2872 23103 2924 23112
rect 2872 23069 2881 23103
rect 2881 23069 2915 23103
rect 2915 23069 2924 23103
rect 2872 23060 2924 23069
rect 4528 23103 4580 23112
rect 4528 23069 4537 23103
rect 4537 23069 4571 23103
rect 4571 23069 4580 23103
rect 4528 23060 4580 23069
rect 6368 23103 6420 23112
rect 6368 23069 6377 23103
rect 6377 23069 6411 23103
rect 6411 23069 6420 23103
rect 6368 23060 6420 23069
rect 9036 23103 9088 23112
rect 9036 23069 9045 23103
rect 9045 23069 9079 23103
rect 9079 23069 9088 23103
rect 9036 23060 9088 23069
rect 12532 23128 12584 23180
rect 13544 23128 13596 23180
rect 13820 23128 13872 23180
rect 14556 23128 14608 23180
rect 17316 23128 17368 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 19800 23128 19852 23180
rect 24308 23128 24360 23180
rect 3608 22924 3660 22976
rect 7196 22924 7248 22976
rect 9864 22967 9916 22976
rect 9864 22933 9873 22967
rect 9873 22933 9907 22967
rect 9907 22933 9916 22967
rect 9864 22924 9916 22933
rect 11796 22924 11848 22976
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 15752 22992 15804 23044
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18236 23060 18288 23112
rect 18972 23060 19024 23112
rect 17960 22967 18012 22976
rect 17960 22933 17969 22967
rect 17969 22933 18003 22967
rect 18003 22933 18012 22967
rect 17960 22924 18012 22933
rect 18604 22967 18656 22976
rect 18604 22933 18613 22967
rect 18613 22933 18647 22967
rect 18647 22933 18656 22967
rect 18604 22924 18656 22933
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 25228 23264 25280 23316
rect 25872 23264 25924 23316
rect 27528 23264 27580 23316
rect 28172 23264 28224 23316
rect 26148 23196 26200 23248
rect 35440 23264 35492 23316
rect 33140 23239 33192 23248
rect 33140 23205 33149 23239
rect 33149 23205 33183 23239
rect 33183 23205 33192 23239
rect 33140 23196 33192 23205
rect 33692 23196 33744 23248
rect 22100 22992 22152 23044
rect 22284 22992 22336 23044
rect 23388 22992 23440 23044
rect 27528 23060 27580 23112
rect 21456 22924 21508 22976
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 26516 22967 26568 22976
rect 26516 22933 26525 22967
rect 26525 22933 26559 22967
rect 26559 22933 26568 22967
rect 26516 22924 26568 22933
rect 27436 22967 27488 22976
rect 27436 22933 27451 22967
rect 27451 22933 27485 22967
rect 27485 22933 27488 22967
rect 27436 22924 27488 22933
rect 27620 22924 27672 22976
rect 28172 23171 28224 23180
rect 28172 23137 28181 23171
rect 28181 23137 28215 23171
rect 28215 23137 28224 23171
rect 28172 23128 28224 23137
rect 28908 23171 28960 23180
rect 28908 23137 28917 23171
rect 28917 23137 28951 23171
rect 28951 23137 28960 23171
rect 28908 23128 28960 23137
rect 29736 23128 29788 23180
rect 32864 23171 32916 23180
rect 32864 23137 32873 23171
rect 32873 23137 32907 23171
rect 32907 23137 32916 23171
rect 32864 23128 32916 23137
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 28816 23060 28868 23112
rect 30656 23103 30708 23112
rect 30656 23069 30665 23103
rect 30665 23069 30699 23103
rect 30699 23069 30708 23103
rect 30656 23060 30708 23069
rect 28264 22992 28316 23044
rect 28632 22992 28684 23044
rect 29092 22967 29144 22976
rect 29092 22933 29101 22967
rect 29101 22933 29135 22967
rect 29135 22933 29144 22967
rect 29092 22924 29144 22933
rect 29368 22924 29420 22976
rect 29552 22924 29604 22976
rect 30748 22967 30800 22976
rect 30748 22933 30757 22967
rect 30757 22933 30791 22967
rect 30791 22933 30800 22967
rect 30748 22924 30800 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 2872 22720 2924 22772
rect 3792 22720 3844 22772
rect 4528 22720 4580 22772
rect 6368 22763 6420 22772
rect 6368 22729 6377 22763
rect 6377 22729 6411 22763
rect 6411 22729 6420 22763
rect 6368 22720 6420 22729
rect 9680 22720 9732 22772
rect 9864 22720 9916 22772
rect 13636 22720 13688 22772
rect 3608 22627 3660 22636
rect 3608 22593 3642 22627
rect 3642 22593 3660 22627
rect 3608 22584 3660 22593
rect 5264 22584 5316 22636
rect 5816 22584 5868 22636
rect 5448 22559 5500 22568
rect 5448 22525 5457 22559
rect 5457 22525 5491 22559
rect 5491 22525 5500 22559
rect 5448 22516 5500 22525
rect 4068 22380 4120 22432
rect 5540 22448 5592 22500
rect 7288 22559 7340 22568
rect 7288 22525 7297 22559
rect 7297 22525 7331 22559
rect 7331 22525 7340 22559
rect 7288 22516 7340 22525
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 11060 22584 11112 22636
rect 11888 22652 11940 22704
rect 12440 22652 12492 22704
rect 13912 22720 13964 22772
rect 15200 22763 15252 22772
rect 15200 22729 15209 22763
rect 15209 22729 15243 22763
rect 15243 22729 15252 22763
rect 15200 22720 15252 22729
rect 14464 22652 14516 22704
rect 17960 22720 18012 22772
rect 19616 22720 19668 22772
rect 20536 22720 20588 22772
rect 21180 22720 21232 22772
rect 21456 22720 21508 22772
rect 22284 22720 22336 22772
rect 22652 22720 22704 22772
rect 18604 22652 18656 22704
rect 20352 22627 20404 22636
rect 8116 22516 8168 22568
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 8760 22516 8812 22568
rect 10140 22559 10192 22568
rect 10140 22525 10149 22559
rect 10149 22525 10183 22559
rect 10183 22525 10192 22559
rect 10140 22516 10192 22525
rect 11796 22559 11848 22568
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 11888 22516 11940 22568
rect 16856 22516 16908 22568
rect 17316 22516 17368 22568
rect 20352 22593 20361 22627
rect 20361 22593 20395 22627
rect 20395 22593 20404 22627
rect 20352 22584 20404 22593
rect 20812 22652 20864 22704
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 20076 22559 20128 22568
rect 20076 22525 20085 22559
rect 20085 22525 20119 22559
rect 20119 22525 20128 22559
rect 20076 22516 20128 22525
rect 20720 22516 20772 22568
rect 20904 22559 20956 22568
rect 20904 22525 20913 22559
rect 20913 22525 20947 22559
rect 20947 22525 20956 22559
rect 20904 22516 20956 22525
rect 21732 22584 21784 22636
rect 22836 22627 22888 22636
rect 22836 22593 22845 22627
rect 22845 22593 22879 22627
rect 22879 22593 22888 22627
rect 22836 22584 22888 22593
rect 24584 22720 24636 22772
rect 26424 22720 26476 22772
rect 27436 22720 27488 22772
rect 23388 22584 23440 22636
rect 22652 22516 22704 22568
rect 25320 22627 25372 22636
rect 25320 22593 25329 22627
rect 25329 22593 25363 22627
rect 25363 22593 25372 22627
rect 25320 22584 25372 22593
rect 22192 22448 22244 22500
rect 25780 22516 25832 22568
rect 25964 22559 26016 22568
rect 25964 22525 25973 22559
rect 25973 22525 26007 22559
rect 26007 22525 26016 22559
rect 25964 22516 26016 22525
rect 26516 22584 26568 22636
rect 27068 22584 27120 22636
rect 27528 22584 27580 22636
rect 28172 22720 28224 22772
rect 28356 22720 28408 22772
rect 28448 22720 28500 22772
rect 28908 22627 28960 22636
rect 28908 22593 28917 22627
rect 28917 22593 28951 22627
rect 28951 22593 28960 22627
rect 28908 22584 28960 22593
rect 29184 22627 29236 22636
rect 29184 22593 29193 22627
rect 29193 22593 29227 22627
rect 29227 22593 29236 22627
rect 29184 22584 29236 22593
rect 4528 22380 4580 22432
rect 6092 22423 6144 22432
rect 6092 22389 6101 22423
rect 6101 22389 6135 22423
rect 6135 22389 6144 22423
rect 6092 22380 6144 22389
rect 6920 22380 6972 22432
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 8668 22423 8720 22432
rect 8668 22389 8692 22423
rect 8692 22389 8720 22423
rect 8668 22380 8720 22389
rect 9036 22380 9088 22432
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 10784 22423 10836 22432
rect 10784 22389 10793 22423
rect 10793 22389 10827 22423
rect 10827 22389 10836 22423
rect 10784 22380 10836 22389
rect 13544 22380 13596 22432
rect 15568 22380 15620 22432
rect 19064 22380 19116 22432
rect 19340 22423 19392 22432
rect 19340 22389 19349 22423
rect 19349 22389 19383 22423
rect 19383 22389 19392 22423
rect 19340 22380 19392 22389
rect 22468 22423 22520 22432
rect 22468 22389 22477 22423
rect 22477 22389 22511 22423
rect 22511 22389 22520 22423
rect 22468 22380 22520 22389
rect 23296 22380 23348 22432
rect 23756 22423 23808 22432
rect 23756 22389 23765 22423
rect 23765 22389 23799 22423
rect 23799 22389 23808 22423
rect 23756 22380 23808 22389
rect 24032 22423 24084 22432
rect 24032 22389 24041 22423
rect 24041 22389 24075 22423
rect 24075 22389 24084 22423
rect 24032 22380 24084 22389
rect 28724 22559 28776 22568
rect 28724 22525 28733 22559
rect 28733 22525 28767 22559
rect 28767 22525 28776 22559
rect 28724 22516 28776 22525
rect 28908 22448 28960 22500
rect 29552 22720 29604 22772
rect 30564 22763 30616 22772
rect 30564 22729 30573 22763
rect 30573 22729 30607 22763
rect 30607 22729 30616 22763
rect 30564 22720 30616 22729
rect 30840 22720 30892 22772
rect 30748 22652 30800 22704
rect 29460 22627 29512 22636
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 30288 22627 30340 22636
rect 30288 22593 30297 22627
rect 30297 22593 30331 22627
rect 30331 22593 30340 22627
rect 30288 22584 30340 22593
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 32956 22720 33008 22772
rect 29368 22559 29420 22568
rect 29368 22525 29377 22559
rect 29377 22525 29411 22559
rect 29411 22525 29420 22559
rect 29368 22516 29420 22525
rect 29920 22559 29972 22568
rect 29920 22525 29929 22559
rect 29929 22525 29963 22559
rect 29963 22525 29972 22559
rect 29920 22516 29972 22525
rect 31300 22516 31352 22568
rect 32956 22516 33008 22568
rect 33692 22584 33744 22636
rect 29920 22380 29972 22432
rect 30748 22423 30800 22432
rect 30748 22389 30757 22423
rect 30757 22389 30791 22423
rect 30791 22389 30800 22423
rect 30748 22380 30800 22389
rect 32588 22423 32640 22432
rect 32588 22389 32597 22423
rect 32597 22389 32631 22423
rect 32631 22389 32640 22423
rect 32588 22380 32640 22389
rect 32864 22380 32916 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3792 22176 3844 22228
rect 3976 22176 4028 22228
rect 5816 22219 5868 22228
rect 5816 22185 5825 22219
rect 5825 22185 5859 22219
rect 5859 22185 5868 22219
rect 5816 22176 5868 22185
rect 8484 22108 8536 22160
rect 8760 22108 8812 22160
rect 12440 22219 12492 22228
rect 12440 22185 12449 22219
rect 12449 22185 12483 22219
rect 12483 22185 12492 22219
rect 12440 22176 12492 22185
rect 6920 22015 6972 22024
rect 6920 21981 6938 22015
rect 6938 21981 6972 22015
rect 6920 21972 6972 21981
rect 8300 21972 8352 22024
rect 4804 21904 4856 21956
rect 7564 21947 7616 21956
rect 7564 21913 7598 21947
rect 7598 21913 7616 21947
rect 7564 21904 7616 21913
rect 8484 21904 8536 21956
rect 10784 22015 10836 22024
rect 10784 21981 10802 22015
rect 10802 21981 10836 22015
rect 10784 21972 10836 21981
rect 10968 21972 11020 22024
rect 11520 21972 11572 22024
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 3240 21836 3292 21888
rect 3976 21836 4028 21888
rect 5724 21879 5776 21888
rect 5724 21845 5733 21879
rect 5733 21845 5767 21879
rect 5767 21845 5776 21879
rect 5724 21836 5776 21845
rect 8944 21879 8996 21888
rect 8944 21845 8953 21879
rect 8953 21845 8987 21879
rect 8987 21845 8996 21879
rect 8944 21836 8996 21845
rect 9036 21836 9088 21888
rect 13268 21904 13320 21956
rect 14004 22040 14056 22092
rect 17500 22176 17552 22228
rect 18144 22176 18196 22228
rect 20812 22176 20864 22228
rect 22100 22219 22152 22228
rect 22100 22185 22109 22219
rect 22109 22185 22143 22219
rect 22143 22185 22152 22219
rect 22100 22176 22152 22185
rect 25964 22176 26016 22228
rect 29184 22176 29236 22228
rect 30288 22176 30340 22228
rect 30380 22176 30432 22228
rect 32588 22176 32640 22228
rect 17132 22108 17184 22160
rect 20536 22151 20588 22160
rect 20536 22117 20545 22151
rect 20545 22117 20579 22151
rect 20579 22117 20588 22151
rect 20536 22108 20588 22117
rect 20628 22108 20680 22160
rect 24400 22108 24452 22160
rect 29920 22108 29972 22160
rect 31300 22108 31352 22160
rect 20076 22040 20128 22092
rect 14004 21836 14056 21888
rect 16580 21972 16632 22024
rect 14648 21904 14700 21956
rect 19340 21972 19392 22024
rect 15108 21879 15160 21888
rect 15108 21845 15117 21879
rect 15117 21845 15151 21879
rect 15151 21845 15160 21879
rect 15108 21836 15160 21845
rect 15568 21879 15620 21888
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 15752 21879 15804 21888
rect 15752 21845 15761 21879
rect 15761 21845 15795 21879
rect 15795 21845 15804 21879
rect 15752 21836 15804 21845
rect 18696 21904 18748 21956
rect 23020 22040 23072 22092
rect 23756 22040 23808 22092
rect 22468 21972 22520 22024
rect 23572 22015 23624 22024
rect 23572 21981 23581 22015
rect 23581 21981 23615 22015
rect 23615 21981 23624 22015
rect 23572 21972 23624 21981
rect 27068 22040 27120 22092
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 26516 21972 26568 22024
rect 28724 22015 28776 22024
rect 28724 21981 28733 22015
rect 28733 21981 28767 22015
rect 28767 21981 28776 22015
rect 28724 21972 28776 21981
rect 29276 22015 29328 22024
rect 29276 21981 29285 22015
rect 29285 21981 29319 22015
rect 29319 21981 29328 22015
rect 29276 21972 29328 21981
rect 29736 22015 29788 22024
rect 29736 21981 29745 22015
rect 29745 21981 29779 22015
rect 29779 21981 29788 22015
rect 29736 21972 29788 21981
rect 30748 22040 30800 22092
rect 31760 22015 31812 22024
rect 31760 21981 31769 22015
rect 31769 21981 31803 22015
rect 31803 21981 31812 22015
rect 31760 21972 31812 21981
rect 32128 21972 32180 22024
rect 18880 21836 18932 21888
rect 20720 21836 20772 21888
rect 21916 21836 21968 21888
rect 23940 21879 23992 21888
rect 23940 21845 23949 21879
rect 23949 21845 23983 21879
rect 23983 21845 23992 21879
rect 23940 21836 23992 21845
rect 24492 21836 24544 21888
rect 28540 21879 28592 21888
rect 28540 21845 28549 21879
rect 28549 21845 28583 21879
rect 28583 21845 28592 21879
rect 28540 21836 28592 21845
rect 29276 21836 29328 21888
rect 30380 21879 30432 21888
rect 30380 21845 30389 21879
rect 30389 21845 30423 21879
rect 30423 21845 30432 21879
rect 30380 21836 30432 21845
rect 30656 21947 30708 21956
rect 30656 21913 30684 21947
rect 30684 21913 30708 21947
rect 30656 21904 30708 21913
rect 32588 21972 32640 22024
rect 32864 21972 32916 22024
rect 33600 22176 33652 22228
rect 33692 21972 33744 22024
rect 32220 21836 32272 21888
rect 33048 21836 33100 21888
rect 33140 21836 33192 21888
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 33784 21836 33836 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 4804 21675 4856 21684
rect 4804 21641 4813 21675
rect 4813 21641 4847 21675
rect 4847 21641 4856 21675
rect 4804 21632 4856 21641
rect 5264 21632 5316 21684
rect 5724 21632 5776 21684
rect 7288 21675 7340 21684
rect 7288 21641 7297 21675
rect 7297 21641 7331 21675
rect 7331 21641 7340 21675
rect 7288 21632 7340 21641
rect 8392 21632 8444 21684
rect 8852 21675 8904 21684
rect 8852 21641 8861 21675
rect 8861 21641 8895 21675
rect 8895 21641 8904 21675
rect 8852 21632 8904 21641
rect 8944 21632 8996 21684
rect 11520 21632 11572 21684
rect 13636 21632 13688 21684
rect 15292 21632 15344 21684
rect 15568 21632 15620 21684
rect 15752 21632 15804 21684
rect 16580 21632 16632 21684
rect 3240 21539 3292 21548
rect 3240 21505 3249 21539
rect 3249 21505 3283 21539
rect 3283 21505 3292 21539
rect 3240 21496 3292 21505
rect 4068 21496 4120 21548
rect 5816 21564 5868 21616
rect 4712 21428 4764 21480
rect 5540 21428 5592 21480
rect 7196 21539 7248 21548
rect 7196 21505 7205 21539
rect 7205 21505 7239 21539
rect 7239 21505 7248 21539
rect 7196 21496 7248 21505
rect 9036 21564 9088 21616
rect 10048 21607 10100 21616
rect 10048 21573 10066 21607
rect 10066 21573 10100 21607
rect 10048 21564 10100 21573
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 8392 21496 8444 21548
rect 12072 21564 12124 21616
rect 14188 21496 14240 21548
rect 15016 21564 15068 21616
rect 8668 21428 8720 21480
rect 8576 21360 8628 21412
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 15108 21539 15160 21548
rect 15108 21505 15117 21539
rect 15117 21505 15151 21539
rect 15151 21505 15160 21539
rect 15108 21496 15160 21505
rect 15568 21496 15620 21548
rect 15660 21428 15712 21480
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 17500 21496 17552 21548
rect 17776 21496 17828 21548
rect 18788 21496 18840 21548
rect 20720 21496 20772 21548
rect 22008 21632 22060 21684
rect 22836 21632 22888 21684
rect 21916 21607 21968 21616
rect 21916 21573 21925 21607
rect 21925 21573 21959 21607
rect 21959 21573 21968 21607
rect 21916 21564 21968 21573
rect 20904 21496 20956 21548
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 15200 21360 15252 21412
rect 15292 21403 15344 21412
rect 15292 21369 15301 21403
rect 15301 21369 15335 21403
rect 15335 21369 15344 21403
rect 15292 21360 15344 21369
rect 3976 21292 4028 21344
rect 5080 21292 5132 21344
rect 8116 21292 8168 21344
rect 12808 21292 12860 21344
rect 13268 21335 13320 21344
rect 13268 21301 13277 21335
rect 13277 21301 13311 21335
rect 13311 21301 13320 21335
rect 13268 21292 13320 21301
rect 14464 21292 14516 21344
rect 14924 21292 14976 21344
rect 20076 21360 20128 21412
rect 20996 21428 21048 21480
rect 23664 21564 23716 21616
rect 30380 21632 30432 21684
rect 30656 21632 30708 21684
rect 31760 21675 31812 21684
rect 31760 21641 31775 21675
rect 31775 21641 31809 21675
rect 31809 21641 31812 21675
rect 31760 21632 31812 21641
rect 32128 21675 32180 21684
rect 32128 21641 32137 21675
rect 32137 21641 32171 21675
rect 32171 21641 32180 21675
rect 32128 21632 32180 21641
rect 32864 21632 32916 21684
rect 33508 21632 33560 21684
rect 23940 21496 23992 21548
rect 21180 21360 21232 21412
rect 15476 21335 15528 21344
rect 15476 21301 15485 21335
rect 15485 21301 15519 21335
rect 15519 21301 15528 21335
rect 15476 21292 15528 21301
rect 16764 21292 16816 21344
rect 17040 21292 17092 21344
rect 17960 21292 18012 21344
rect 19708 21335 19760 21344
rect 19708 21301 19717 21335
rect 19717 21301 19751 21335
rect 19751 21301 19760 21335
rect 19708 21292 19760 21301
rect 24492 21496 24544 21548
rect 24400 21471 24452 21480
rect 24400 21437 24409 21471
rect 24409 21437 24443 21471
rect 24443 21437 24452 21471
rect 28632 21564 28684 21616
rect 24768 21539 24820 21548
rect 24768 21505 24777 21539
rect 24777 21505 24811 21539
rect 24811 21505 24820 21539
rect 24768 21496 24820 21505
rect 24400 21428 24452 21437
rect 23388 21292 23440 21344
rect 24124 21292 24176 21344
rect 26056 21496 26108 21548
rect 26516 21428 26568 21480
rect 31944 21539 31996 21548
rect 31944 21505 31953 21539
rect 31953 21505 31987 21539
rect 31987 21505 31996 21539
rect 31944 21496 31996 21505
rect 32404 21471 32456 21480
rect 32404 21437 32413 21471
rect 32413 21437 32447 21471
rect 32447 21437 32456 21471
rect 32404 21428 32456 21437
rect 33048 21496 33100 21548
rect 25872 21335 25924 21344
rect 25872 21301 25881 21335
rect 25881 21301 25915 21335
rect 25915 21301 25924 21335
rect 25872 21292 25924 21301
rect 27620 21292 27672 21344
rect 31484 21292 31536 21344
rect 31576 21292 31628 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4712 21088 4764 21140
rect 5356 21088 5408 21140
rect 5540 21131 5592 21140
rect 5540 21097 5549 21131
rect 5549 21097 5583 21131
rect 5583 21097 5592 21131
rect 5540 21088 5592 21097
rect 9036 21088 9088 21140
rect 10140 21088 10192 21140
rect 11796 21131 11848 21140
rect 11796 21097 11805 21131
rect 11805 21097 11839 21131
rect 11839 21097 11848 21131
rect 11796 21088 11848 21097
rect 12072 21131 12124 21140
rect 12072 21097 12081 21131
rect 12081 21097 12115 21131
rect 12115 21097 12124 21131
rect 12072 21088 12124 21097
rect 17684 21088 17736 21140
rect 19708 21088 19760 21140
rect 5264 20952 5316 21004
rect 8116 20952 8168 21004
rect 5080 20927 5132 20936
rect 5080 20893 5089 20927
rect 5089 20893 5123 20927
rect 5123 20893 5132 20927
rect 5080 20884 5132 20893
rect 5448 20927 5500 20936
rect 5448 20893 5457 20927
rect 5457 20893 5491 20927
rect 5491 20893 5500 20927
rect 5448 20884 5500 20893
rect 6092 20884 6144 20936
rect 15108 21063 15160 21072
rect 15108 21029 15117 21063
rect 15117 21029 15151 21063
rect 15151 21029 15160 21063
rect 15108 21020 15160 21029
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 14096 20884 14148 20936
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 14924 20927 14976 20936
rect 14924 20893 14934 20927
rect 14934 20893 14968 20927
rect 14968 20893 14976 20927
rect 14924 20884 14976 20893
rect 15292 20884 15344 20936
rect 16580 20884 16632 20936
rect 11060 20748 11112 20800
rect 15384 20859 15436 20868
rect 15384 20825 15393 20859
rect 15393 20825 15427 20859
rect 15427 20825 15436 20859
rect 15384 20816 15436 20825
rect 17960 20884 18012 20936
rect 16856 20816 16908 20868
rect 15660 20748 15712 20800
rect 15844 20748 15896 20800
rect 18696 20859 18748 20868
rect 18696 20825 18705 20859
rect 18705 20825 18739 20859
rect 18739 20825 18748 20859
rect 18696 20816 18748 20825
rect 21548 20952 21600 21004
rect 25320 21088 25372 21140
rect 25504 21088 25556 21140
rect 25872 21088 25924 21140
rect 28448 21088 28500 21140
rect 27620 21020 27672 21072
rect 28540 21020 28592 21072
rect 30380 21088 30432 21140
rect 33140 21131 33192 21140
rect 33140 21097 33149 21131
rect 33149 21097 33183 21131
rect 33183 21097 33192 21131
rect 33140 21088 33192 21097
rect 28816 21020 28868 21072
rect 31576 21020 31628 21072
rect 26056 20995 26108 21004
rect 26056 20961 26065 20995
rect 26065 20961 26099 20995
rect 26099 20961 26108 20995
rect 26056 20952 26108 20961
rect 22560 20884 22612 20936
rect 22652 20927 22704 20936
rect 22652 20893 22661 20927
rect 22661 20893 22695 20927
rect 22695 20893 22704 20927
rect 22652 20884 22704 20893
rect 25320 20884 25372 20936
rect 25688 20884 25740 20936
rect 27988 20884 28040 20936
rect 28448 20927 28500 20936
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 20812 20816 20864 20868
rect 21088 20859 21140 20868
rect 21088 20825 21097 20859
rect 21097 20825 21131 20859
rect 21131 20825 21140 20859
rect 21088 20816 21140 20825
rect 23388 20816 23440 20868
rect 17316 20748 17368 20800
rect 19524 20791 19576 20800
rect 19524 20757 19533 20791
rect 19533 20757 19567 20791
rect 19567 20757 19576 20791
rect 19524 20748 19576 20757
rect 19984 20748 20036 20800
rect 20168 20748 20220 20800
rect 23756 20748 23808 20800
rect 25412 20791 25464 20800
rect 25412 20757 25421 20791
rect 25421 20757 25455 20791
rect 25455 20757 25464 20791
rect 25412 20748 25464 20757
rect 25596 20859 25648 20868
rect 25596 20825 25605 20859
rect 25605 20825 25639 20859
rect 25639 20825 25648 20859
rect 25596 20816 25648 20825
rect 25780 20859 25832 20868
rect 25780 20825 25789 20859
rect 25789 20825 25823 20859
rect 25823 20825 25832 20859
rect 25780 20816 25832 20825
rect 26056 20748 26108 20800
rect 26332 20791 26384 20800
rect 26332 20757 26341 20791
rect 26341 20757 26375 20791
rect 26375 20757 26384 20791
rect 26332 20748 26384 20757
rect 27712 20748 27764 20800
rect 28356 20816 28408 20868
rect 28724 20884 28776 20936
rect 30104 20927 30156 20936
rect 30104 20893 30113 20927
rect 30113 20893 30147 20927
rect 30147 20893 30156 20927
rect 30104 20884 30156 20893
rect 31484 20927 31536 20936
rect 31484 20893 31493 20927
rect 31493 20893 31527 20927
rect 31527 20893 31536 20927
rect 31484 20884 31536 20893
rect 30288 20859 30340 20868
rect 30288 20825 30297 20859
rect 30297 20825 30331 20859
rect 30331 20825 30340 20859
rect 30288 20816 30340 20825
rect 31392 20816 31444 20868
rect 28632 20748 28684 20800
rect 33048 20748 33100 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 4068 20544 4120 20596
rect 15200 20544 15252 20596
rect 16580 20544 16632 20596
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 11060 20408 11112 20460
rect 11704 20408 11756 20460
rect 11980 20340 12032 20392
rect 13084 20476 13136 20528
rect 13544 20451 13596 20460
rect 12716 20340 12768 20392
rect 11612 20272 11664 20324
rect 12532 20272 12584 20324
rect 13268 20340 13320 20392
rect 13544 20417 13554 20451
rect 13554 20417 13596 20451
rect 13544 20408 13596 20417
rect 15016 20408 15068 20460
rect 20628 20544 20680 20596
rect 20720 20587 20772 20596
rect 20720 20553 20729 20587
rect 20729 20553 20763 20587
rect 20763 20553 20772 20587
rect 20720 20544 20772 20553
rect 21088 20544 21140 20596
rect 14004 20340 14056 20392
rect 15108 20340 15160 20392
rect 16856 20340 16908 20392
rect 17960 20408 18012 20460
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 19524 20476 19576 20528
rect 19984 20476 20036 20528
rect 17408 20383 17460 20392
rect 17408 20349 17417 20383
rect 17417 20349 17451 20383
rect 17451 20349 17460 20383
rect 17408 20340 17460 20349
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 17776 20383 17828 20392
rect 17776 20349 17785 20383
rect 17785 20349 17819 20383
rect 17819 20349 17828 20383
rect 17776 20340 17828 20349
rect 20812 20408 20864 20460
rect 23296 20476 23348 20528
rect 14740 20272 14792 20324
rect 22100 20340 22152 20392
rect 22560 20408 22612 20460
rect 23480 20451 23532 20460
rect 23480 20417 23489 20451
rect 23489 20417 23523 20451
rect 23523 20417 23532 20451
rect 23480 20408 23532 20417
rect 23572 20408 23624 20460
rect 24124 20519 24176 20528
rect 24124 20485 24133 20519
rect 24133 20485 24167 20519
rect 24167 20485 24176 20519
rect 24124 20476 24176 20485
rect 25412 20544 25464 20596
rect 25780 20544 25832 20596
rect 27712 20544 27764 20596
rect 28356 20587 28408 20596
rect 28356 20553 28365 20587
rect 28365 20553 28399 20587
rect 28399 20553 28408 20587
rect 28356 20544 28408 20553
rect 28724 20544 28776 20596
rect 31944 20544 31996 20596
rect 23848 20408 23900 20460
rect 22468 20383 22520 20392
rect 22468 20349 22477 20383
rect 22477 20349 22511 20383
rect 22511 20349 22520 20383
rect 22468 20340 22520 20349
rect 24860 20451 24912 20460
rect 24860 20417 24869 20451
rect 24869 20417 24903 20451
rect 24903 20417 24912 20451
rect 24860 20408 24912 20417
rect 25320 20451 25372 20460
rect 25320 20417 25329 20451
rect 25329 20417 25363 20451
rect 25363 20417 25372 20451
rect 25320 20408 25372 20417
rect 25504 20408 25556 20460
rect 25688 20408 25740 20460
rect 26332 20451 26384 20460
rect 26332 20417 26341 20451
rect 26341 20417 26375 20451
rect 26375 20417 26384 20451
rect 26332 20408 26384 20417
rect 22192 20272 22244 20324
rect 22836 20272 22888 20324
rect 23388 20272 23440 20324
rect 9312 20204 9364 20256
rect 9864 20247 9916 20256
rect 9864 20213 9873 20247
rect 9873 20213 9907 20247
rect 9907 20213 9916 20247
rect 9864 20204 9916 20213
rect 11888 20247 11940 20256
rect 11888 20213 11897 20247
rect 11897 20213 11931 20247
rect 11931 20213 11940 20247
rect 11888 20204 11940 20213
rect 12716 20204 12768 20256
rect 13728 20204 13780 20256
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 17868 20204 17920 20256
rect 18052 20204 18104 20256
rect 19064 20204 19116 20256
rect 23572 20204 23624 20256
rect 25412 20272 25464 20324
rect 26148 20315 26200 20324
rect 26148 20281 26157 20315
rect 26157 20281 26191 20315
rect 26191 20281 26200 20315
rect 26148 20272 26200 20281
rect 27620 20408 27672 20460
rect 24768 20204 24820 20256
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 27988 20340 28040 20392
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29092 20408 29144 20460
rect 29276 20451 29328 20460
rect 29276 20417 29285 20451
rect 29285 20417 29319 20451
rect 29319 20417 29328 20451
rect 29276 20408 29328 20417
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 30012 20408 30064 20460
rect 30104 20408 30156 20460
rect 30840 20451 30892 20460
rect 30840 20417 30849 20451
rect 30849 20417 30883 20451
rect 30883 20417 30892 20451
rect 30840 20408 30892 20417
rect 31300 20451 31352 20460
rect 31300 20417 31309 20451
rect 31309 20417 31343 20451
rect 31343 20417 31352 20451
rect 31300 20408 31352 20417
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 30288 20272 30340 20324
rect 33140 20408 33192 20460
rect 33692 20408 33744 20460
rect 34336 20408 34388 20460
rect 32956 20272 33008 20324
rect 26792 20204 26844 20256
rect 26976 20247 27028 20256
rect 26976 20213 26985 20247
rect 26985 20213 27019 20247
rect 27019 20213 27028 20247
rect 26976 20204 27028 20213
rect 27436 20204 27488 20256
rect 29644 20204 29696 20256
rect 29736 20247 29788 20256
rect 29736 20213 29745 20247
rect 29745 20213 29779 20247
rect 29779 20213 29788 20247
rect 29736 20204 29788 20213
rect 30472 20204 30524 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 14004 20000 14056 20052
rect 14648 20000 14700 20052
rect 15200 20000 15252 20052
rect 17868 20000 17920 20052
rect 11980 19975 12032 19984
rect 11980 19941 11989 19975
rect 11989 19941 12023 19975
rect 12023 19941 12032 19975
rect 11980 19932 12032 19941
rect 9312 19864 9364 19916
rect 8300 19796 8352 19848
rect 10968 19796 11020 19848
rect 9864 19728 9916 19780
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 12624 19932 12676 19984
rect 13912 19932 13964 19984
rect 17592 19932 17644 19984
rect 20996 20000 21048 20052
rect 23480 20000 23532 20052
rect 25044 20000 25096 20052
rect 29644 20000 29696 20052
rect 22100 19932 22152 19984
rect 23388 19932 23440 19984
rect 24860 19932 24912 19984
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 13360 19864 13412 19916
rect 14188 19864 14240 19916
rect 11888 19796 11940 19805
rect 12716 19796 12768 19848
rect 13728 19796 13780 19848
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 14924 19839 14976 19848
rect 14924 19805 14933 19839
rect 14933 19805 14967 19839
rect 14967 19805 14976 19839
rect 14924 19796 14976 19805
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 18972 19907 19024 19916
rect 18972 19873 18981 19907
rect 18981 19873 19015 19907
rect 19015 19873 19024 19907
rect 18972 19864 19024 19873
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 24768 19907 24820 19916
rect 24768 19873 24777 19907
rect 24777 19873 24811 19907
rect 24811 19873 24820 19907
rect 24768 19864 24820 19873
rect 15844 19839 15896 19848
rect 15844 19805 15879 19839
rect 15879 19805 15896 19839
rect 15844 19796 15896 19805
rect 16120 19796 16172 19848
rect 17776 19796 17828 19848
rect 18420 19796 18472 19848
rect 9956 19660 10008 19712
rect 15384 19728 15436 19780
rect 10692 19703 10744 19712
rect 10692 19669 10701 19703
rect 10701 19669 10735 19703
rect 10735 19669 10744 19703
rect 10692 19660 10744 19669
rect 11704 19660 11756 19712
rect 13728 19660 13780 19712
rect 27528 19932 27580 19984
rect 29920 20000 29972 20052
rect 30748 20000 30800 20052
rect 30840 20000 30892 20052
rect 25596 19796 25648 19848
rect 26148 19796 26200 19848
rect 26332 19839 26384 19848
rect 26332 19805 26341 19839
rect 26341 19805 26375 19839
rect 26375 19805 26384 19839
rect 26332 19796 26384 19805
rect 26792 19839 26844 19848
rect 26792 19805 26801 19839
rect 26801 19805 26835 19839
rect 26835 19805 26844 19839
rect 26792 19796 26844 19805
rect 27712 19864 27764 19916
rect 33140 20000 33192 20052
rect 32772 19907 32824 19916
rect 32772 19873 32781 19907
rect 32781 19873 32815 19907
rect 32815 19873 32824 19907
rect 32772 19864 32824 19873
rect 33416 19864 33468 19916
rect 27436 19839 27488 19848
rect 27436 19805 27445 19839
rect 27445 19805 27479 19839
rect 27479 19805 27488 19839
rect 27436 19796 27488 19805
rect 24124 19728 24176 19780
rect 28448 19796 28500 19848
rect 30472 19839 30524 19848
rect 30472 19805 30481 19839
rect 30481 19805 30515 19839
rect 30515 19805 30524 19839
rect 30472 19796 30524 19805
rect 29000 19728 29052 19780
rect 29644 19728 29696 19780
rect 16304 19660 16356 19712
rect 18604 19660 18656 19712
rect 19616 19660 19668 19712
rect 27068 19660 27120 19712
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 29092 19660 29144 19712
rect 30288 19728 30340 19780
rect 31392 19796 31444 19848
rect 31024 19660 31076 19712
rect 32036 19839 32088 19848
rect 32036 19805 32045 19839
rect 32045 19805 32079 19839
rect 32079 19805 32088 19839
rect 32036 19796 32088 19805
rect 32220 19796 32272 19848
rect 33048 19839 33100 19848
rect 33048 19805 33057 19839
rect 33057 19805 33091 19839
rect 33091 19805 33100 19839
rect 33048 19796 33100 19805
rect 32404 19728 32456 19780
rect 32588 19728 32640 19780
rect 35532 19728 35584 19780
rect 33784 19703 33836 19712
rect 33784 19669 33793 19703
rect 33793 19669 33827 19703
rect 33827 19669 33836 19703
rect 33784 19660 33836 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 4068 19456 4120 19508
rect 9956 19456 10008 19508
rect 14280 19456 14332 19508
rect 15108 19499 15160 19508
rect 15108 19465 15117 19499
rect 15117 19465 15151 19499
rect 15151 19465 15160 19499
rect 15108 19456 15160 19465
rect 3424 19388 3476 19440
rect 12992 19388 13044 19440
rect 15568 19456 15620 19508
rect 16212 19456 16264 19508
rect 16304 19499 16356 19508
rect 16304 19465 16313 19499
rect 16313 19465 16347 19499
rect 16347 19465 16356 19499
rect 16304 19456 16356 19465
rect 18972 19456 19024 19508
rect 10692 19320 10744 19372
rect 10968 19320 11020 19372
rect 11152 19320 11204 19372
rect 13544 19320 13596 19372
rect 13728 19320 13780 19372
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14464 19320 14516 19372
rect 16672 19431 16724 19440
rect 16672 19397 16681 19431
rect 16681 19397 16715 19431
rect 16715 19397 16724 19431
rect 16672 19388 16724 19397
rect 17684 19388 17736 19440
rect 15476 19252 15528 19304
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 18512 19363 18564 19372
rect 16396 19320 16448 19329
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20628 19320 20680 19372
rect 20904 19388 20956 19440
rect 22376 19456 22428 19508
rect 24032 19456 24084 19508
rect 25688 19499 25740 19508
rect 25688 19465 25697 19499
rect 25697 19465 25731 19499
rect 25731 19465 25740 19499
rect 25688 19456 25740 19465
rect 21824 19363 21876 19372
rect 21824 19329 21833 19363
rect 21833 19329 21867 19363
rect 21867 19329 21876 19363
rect 21824 19320 21876 19329
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 22836 19320 22888 19372
rect 23940 19320 23992 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 21180 19252 21232 19304
rect 19248 19184 19300 19236
rect 24032 19252 24084 19304
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 25412 19320 25464 19372
rect 26976 19320 27028 19372
rect 29460 19388 29512 19440
rect 29736 19456 29788 19508
rect 31024 19499 31076 19508
rect 31024 19465 31033 19499
rect 31033 19465 31067 19499
rect 31067 19465 31076 19499
rect 31024 19456 31076 19465
rect 30564 19388 30616 19440
rect 32036 19456 32088 19508
rect 32588 19456 32640 19508
rect 33416 19456 33468 19508
rect 33784 19456 33836 19508
rect 34336 19499 34388 19508
rect 34336 19465 34345 19499
rect 34345 19465 34379 19499
rect 34379 19465 34388 19499
rect 34336 19456 34388 19465
rect 32220 19388 32272 19440
rect 32956 19363 33008 19372
rect 32956 19329 32965 19363
rect 32965 19329 32999 19363
rect 32999 19329 33008 19363
rect 32956 19320 33008 19329
rect 25872 19252 25924 19304
rect 27712 19252 27764 19304
rect 33324 19295 33376 19304
rect 33324 19261 33333 19295
rect 33333 19261 33367 19295
rect 33367 19261 33376 19295
rect 33324 19252 33376 19261
rect 13636 19116 13688 19168
rect 18144 19116 18196 19168
rect 20536 19116 20588 19168
rect 20812 19116 20864 19168
rect 23204 19116 23256 19168
rect 23296 19159 23348 19168
rect 23296 19125 23305 19159
rect 23305 19125 23339 19159
rect 23339 19125 23348 19159
rect 23296 19116 23348 19125
rect 23572 19116 23624 19168
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 27528 19159 27580 19168
rect 27528 19125 27537 19159
rect 27537 19125 27571 19159
rect 27571 19125 27580 19159
rect 27528 19116 27580 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10876 18912 10928 18964
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 13176 18912 13228 18964
rect 13268 18912 13320 18964
rect 17960 18955 18012 18964
rect 17960 18921 17969 18955
rect 17969 18921 18003 18955
rect 18003 18921 18012 18955
rect 17960 18912 18012 18921
rect 18512 18912 18564 18964
rect 20628 18912 20680 18964
rect 22468 18912 22520 18964
rect 22836 18912 22888 18964
rect 14556 18844 14608 18896
rect 12716 18819 12768 18828
rect 12716 18785 12725 18819
rect 12725 18785 12759 18819
rect 12759 18785 12768 18819
rect 12716 18776 12768 18785
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 13360 18776 13412 18828
rect 13544 18708 13596 18760
rect 14740 18776 14792 18828
rect 15476 18776 15528 18828
rect 19156 18844 19208 18896
rect 14464 18708 14516 18760
rect 15108 18708 15160 18760
rect 15384 18708 15436 18760
rect 16120 18708 16172 18760
rect 16304 18751 16356 18760
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 16764 18708 16816 18760
rect 12992 18683 13044 18692
rect 12992 18649 13001 18683
rect 13001 18649 13035 18683
rect 13035 18649 13044 18683
rect 12992 18640 13044 18649
rect 17592 18751 17644 18760
rect 17592 18717 17601 18751
rect 17601 18717 17635 18751
rect 17635 18717 17644 18751
rect 17592 18708 17644 18717
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 18144 18708 18196 18760
rect 9864 18572 9916 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 14924 18572 14976 18624
rect 18144 18572 18196 18624
rect 19708 18776 19760 18828
rect 20720 18776 20772 18828
rect 21824 18776 21876 18828
rect 23848 18912 23900 18964
rect 24032 18912 24084 18964
rect 25412 18912 25464 18964
rect 28724 18955 28776 18964
rect 28724 18921 28733 18955
rect 28733 18921 28767 18955
rect 28767 18921 28776 18955
rect 28724 18912 28776 18921
rect 30012 18912 30064 18964
rect 30564 18912 30616 18964
rect 18788 18708 18840 18760
rect 20444 18640 20496 18692
rect 23204 18708 23256 18760
rect 24860 18844 24912 18896
rect 26056 18844 26108 18896
rect 24124 18776 24176 18828
rect 27528 18776 27580 18828
rect 26976 18751 27028 18760
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 21548 18640 21600 18692
rect 26976 18717 26985 18751
rect 26985 18717 27019 18751
rect 27019 18717 27028 18751
rect 26976 18708 27028 18717
rect 27068 18708 27120 18760
rect 29184 18708 29236 18760
rect 30380 18776 30432 18828
rect 18328 18572 18380 18624
rect 18604 18572 18656 18624
rect 19432 18572 19484 18624
rect 20904 18572 20956 18624
rect 21088 18572 21140 18624
rect 21732 18615 21784 18624
rect 21732 18581 21741 18615
rect 21741 18581 21775 18615
rect 21775 18581 21784 18615
rect 21732 18572 21784 18581
rect 25412 18683 25464 18692
rect 25412 18649 25421 18683
rect 25421 18649 25455 18683
rect 25455 18649 25464 18683
rect 25412 18640 25464 18649
rect 26148 18640 26200 18692
rect 35440 18844 35492 18896
rect 23204 18572 23256 18624
rect 27528 18615 27580 18624
rect 27528 18581 27537 18615
rect 27537 18581 27571 18615
rect 27571 18581 27580 18615
rect 27528 18572 27580 18581
rect 30840 18615 30892 18624
rect 30840 18581 30849 18615
rect 30849 18581 30883 18615
rect 30883 18581 30892 18615
rect 30840 18572 30892 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 11520 18368 11572 18420
rect 12164 18368 12216 18420
rect 14372 18368 14424 18420
rect 14464 18368 14516 18420
rect 16304 18368 16356 18420
rect 9772 18300 9824 18352
rect 16764 18300 16816 18352
rect 12992 18232 13044 18284
rect 15384 18275 15436 18284
rect 15384 18241 15393 18275
rect 15393 18241 15427 18275
rect 15427 18241 15436 18275
rect 15384 18232 15436 18241
rect 4068 18164 4120 18216
rect 8300 18164 8352 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 12532 18207 12584 18216
rect 12532 18173 12541 18207
rect 12541 18173 12575 18207
rect 12575 18173 12584 18207
rect 12532 18164 12584 18173
rect 14280 18164 14332 18216
rect 17776 18368 17828 18420
rect 18328 18343 18380 18352
rect 18328 18309 18337 18343
rect 18337 18309 18371 18343
rect 18371 18309 18380 18343
rect 18328 18300 18380 18309
rect 19708 18368 19760 18420
rect 20536 18368 20588 18420
rect 23296 18368 23348 18420
rect 23664 18368 23716 18420
rect 23940 18368 23992 18420
rect 25320 18368 25372 18420
rect 26148 18411 26200 18420
rect 26148 18377 26157 18411
rect 26157 18377 26191 18411
rect 26191 18377 26200 18411
rect 26148 18368 26200 18377
rect 19156 18275 19208 18284
rect 19156 18241 19165 18275
rect 19165 18241 19199 18275
rect 19199 18241 19208 18275
rect 19156 18232 19208 18241
rect 20260 18232 20312 18284
rect 20904 18343 20956 18352
rect 20904 18309 20913 18343
rect 20913 18309 20947 18343
rect 20947 18309 20956 18343
rect 20904 18300 20956 18309
rect 16764 18139 16816 18148
rect 16764 18105 16773 18139
rect 16773 18105 16807 18139
rect 16807 18105 16816 18139
rect 16764 18096 16816 18105
rect 17408 18096 17460 18148
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 19524 18207 19576 18216
rect 19524 18173 19533 18207
rect 19533 18173 19567 18207
rect 19567 18173 19576 18207
rect 19524 18164 19576 18173
rect 19984 18164 20036 18216
rect 21088 18139 21140 18148
rect 9864 18028 9916 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 16120 18028 16172 18080
rect 21088 18105 21097 18139
rect 21097 18105 21131 18139
rect 21131 18105 21140 18139
rect 21088 18096 21140 18105
rect 21732 18164 21784 18216
rect 23480 18096 23532 18148
rect 24860 18300 24912 18352
rect 27528 18368 27580 18420
rect 30840 18300 30892 18352
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 32496 18275 32548 18284
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 18604 18028 18656 18080
rect 20444 18028 20496 18080
rect 25320 18139 25372 18148
rect 25320 18105 25329 18139
rect 25329 18105 25363 18139
rect 25363 18105 25372 18139
rect 27620 18207 27672 18216
rect 27620 18173 27629 18207
rect 27629 18173 27663 18207
rect 27663 18173 27672 18207
rect 27620 18164 27672 18173
rect 29460 18164 29512 18216
rect 25320 18096 25372 18105
rect 26608 18071 26660 18080
rect 26608 18037 26617 18071
rect 26617 18037 26651 18071
rect 26651 18037 26660 18071
rect 26608 18028 26660 18037
rect 27344 18028 27396 18080
rect 30748 18028 30800 18080
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 35348 18232 35400 18284
rect 33324 18207 33376 18216
rect 33324 18173 33333 18207
rect 33333 18173 33367 18207
rect 33367 18173 33376 18207
rect 33324 18164 33376 18173
rect 32312 18028 32364 18080
rect 32680 18028 32732 18080
rect 34336 18071 34388 18080
rect 34336 18037 34345 18071
rect 34345 18037 34379 18071
rect 34379 18037 34388 18071
rect 34336 18028 34388 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8760 17824 8812 17876
rect 9772 17824 9824 17876
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 12900 17824 12952 17876
rect 14832 17824 14884 17876
rect 21364 17824 21416 17876
rect 22284 17824 22336 17876
rect 14280 17756 14332 17808
rect 10876 17731 10928 17740
rect 10876 17697 10885 17731
rect 10885 17697 10919 17731
rect 10919 17697 10928 17731
rect 10876 17688 10928 17697
rect 11612 17688 11664 17740
rect 20260 17756 20312 17808
rect 21640 17756 21692 17808
rect 21824 17756 21876 17808
rect 9220 17663 9272 17672
rect 9220 17629 9229 17663
rect 9229 17629 9263 17663
rect 9263 17629 9272 17663
rect 9220 17620 9272 17629
rect 9680 17620 9732 17672
rect 10232 17620 10284 17672
rect 12532 17620 12584 17672
rect 12992 17620 13044 17672
rect 14556 17620 14608 17672
rect 14832 17620 14884 17672
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 14740 17552 14792 17604
rect 19984 17688 20036 17740
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 25228 17824 25280 17876
rect 25780 17824 25832 17876
rect 27344 17824 27396 17876
rect 29552 17824 29604 17876
rect 32496 17824 32548 17876
rect 32956 17824 33008 17876
rect 33508 17867 33560 17876
rect 33508 17833 33517 17867
rect 33517 17833 33551 17867
rect 33551 17833 33560 17867
rect 33508 17824 33560 17833
rect 34336 17824 34388 17876
rect 25688 17688 25740 17740
rect 34060 17756 34112 17808
rect 17684 17620 17736 17672
rect 9128 17484 9180 17536
rect 12716 17527 12768 17536
rect 12716 17493 12725 17527
rect 12725 17493 12759 17527
rect 12759 17493 12768 17527
rect 12716 17484 12768 17493
rect 14096 17527 14148 17536
rect 14096 17493 14105 17527
rect 14105 17493 14139 17527
rect 14139 17493 14148 17527
rect 14096 17484 14148 17493
rect 17040 17484 17092 17536
rect 18788 17620 18840 17672
rect 19524 17620 19576 17672
rect 21732 17620 21784 17672
rect 20628 17552 20680 17604
rect 20904 17552 20956 17604
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 22008 17552 22060 17604
rect 24032 17663 24084 17672
rect 24032 17629 24041 17663
rect 24041 17629 24075 17663
rect 24075 17629 24084 17663
rect 24032 17620 24084 17629
rect 25320 17620 25372 17672
rect 29184 17688 29236 17740
rect 29552 17688 29604 17740
rect 30196 17688 30248 17740
rect 32496 17688 32548 17740
rect 21732 17484 21784 17536
rect 22192 17484 22244 17536
rect 22744 17484 22796 17536
rect 23020 17527 23072 17536
rect 23020 17493 23029 17527
rect 23029 17493 23063 17527
rect 23063 17493 23072 17527
rect 23020 17484 23072 17493
rect 23204 17527 23256 17536
rect 23204 17493 23213 17527
rect 23213 17493 23247 17527
rect 23247 17493 23256 17527
rect 23204 17484 23256 17493
rect 23296 17484 23348 17536
rect 26608 17595 26660 17604
rect 26608 17561 26617 17595
rect 26617 17561 26651 17595
rect 26651 17561 26660 17595
rect 26608 17552 26660 17561
rect 29368 17620 29420 17672
rect 30564 17620 30616 17672
rect 31300 17620 31352 17672
rect 32404 17552 32456 17604
rect 33508 17620 33560 17672
rect 32864 17552 32916 17604
rect 27528 17484 27580 17536
rect 28356 17484 28408 17536
rect 28632 17484 28684 17536
rect 30104 17527 30156 17536
rect 30104 17493 30113 17527
rect 30113 17493 30147 17527
rect 30147 17493 30156 17527
rect 30104 17484 30156 17493
rect 30656 17527 30708 17536
rect 30656 17493 30665 17527
rect 30665 17493 30699 17527
rect 30699 17493 30708 17527
rect 30656 17484 30708 17493
rect 30748 17527 30800 17536
rect 30748 17493 30757 17527
rect 30757 17493 30791 17527
rect 30791 17493 30800 17527
rect 30748 17484 30800 17493
rect 32220 17484 32272 17536
rect 33048 17484 33100 17536
rect 33692 17527 33744 17536
rect 33692 17493 33701 17527
rect 33701 17493 33735 17527
rect 33735 17493 33744 17527
rect 33692 17484 33744 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 11612 17280 11664 17332
rect 12716 17280 12768 17332
rect 11336 17212 11388 17264
rect 15108 17280 15160 17332
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 14648 17144 14700 17196
rect 14924 17144 14976 17196
rect 18880 17280 18932 17332
rect 17408 17212 17460 17264
rect 22744 17280 22796 17332
rect 23756 17280 23808 17332
rect 24032 17280 24084 17332
rect 18420 17144 18472 17196
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 10968 17076 11020 17128
rect 17868 17076 17920 17128
rect 16948 17051 17000 17060
rect 16948 17017 16957 17051
rect 16957 17017 16991 17051
rect 16991 17017 17000 17051
rect 16948 17008 17000 17017
rect 17040 17008 17092 17060
rect 8300 16940 8352 16992
rect 11980 16940 12032 16992
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 17776 16940 17828 16992
rect 18972 16940 19024 16992
rect 21456 17187 21508 17196
rect 21456 17153 21465 17187
rect 21465 17153 21499 17187
rect 21499 17153 21508 17187
rect 21456 17144 21508 17153
rect 23204 17144 23256 17196
rect 28632 17212 28684 17264
rect 30656 17280 30708 17332
rect 32220 17280 32272 17332
rect 33048 17280 33100 17332
rect 25688 17187 25740 17196
rect 25688 17153 25699 17187
rect 25699 17153 25733 17187
rect 25733 17153 25740 17187
rect 25688 17144 25740 17153
rect 25780 17144 25832 17196
rect 29552 17144 29604 17196
rect 29828 17187 29880 17196
rect 29828 17153 29837 17187
rect 29837 17153 29871 17187
rect 29871 17153 29880 17187
rect 29828 17144 29880 17153
rect 32404 17255 32456 17264
rect 32404 17221 32413 17255
rect 32413 17221 32447 17255
rect 32447 17221 32456 17255
rect 32404 17212 32456 17221
rect 32588 17255 32640 17264
rect 32588 17221 32597 17255
rect 32597 17221 32631 17255
rect 32631 17221 32640 17255
rect 32588 17212 32640 17221
rect 32772 17212 32824 17264
rect 33232 17144 33284 17196
rect 20720 17076 20772 17128
rect 21824 17119 21876 17128
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 23296 17076 23348 17128
rect 24860 17008 24912 17060
rect 23204 16940 23256 16992
rect 27528 17076 27580 17128
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 29920 17119 29972 17128
rect 29920 17085 29929 17119
rect 29929 17085 29963 17119
rect 29963 17085 29972 17119
rect 29920 17076 29972 17085
rect 30196 17076 30248 17128
rect 29276 17008 29328 17060
rect 31668 17076 31720 17128
rect 32404 17008 32456 17060
rect 28356 16940 28408 16992
rect 31024 16983 31076 16992
rect 31024 16949 31033 16983
rect 31033 16949 31067 16983
rect 31067 16949 31076 16983
rect 31024 16940 31076 16949
rect 31300 16940 31352 16992
rect 32864 16983 32916 16992
rect 32864 16949 32873 16983
rect 32873 16949 32907 16983
rect 32907 16949 32916 16983
rect 32864 16940 32916 16949
rect 33048 16983 33100 16992
rect 33048 16949 33057 16983
rect 33057 16949 33091 16983
rect 33091 16949 33100 16983
rect 38844 17076 38896 17128
rect 33048 16940 33100 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 9220 16736 9272 16788
rect 10232 16736 10284 16788
rect 12716 16736 12768 16788
rect 13820 16736 13872 16788
rect 14280 16736 14332 16788
rect 14464 16736 14516 16788
rect 10324 16600 10376 16652
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11152 16600 11204 16652
rect 9956 16532 10008 16584
rect 10692 16532 10744 16584
rect 13728 16668 13780 16720
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 9404 16507 9456 16516
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 12164 16464 12216 16516
rect 13544 16532 13596 16584
rect 20720 16736 20772 16788
rect 21456 16736 21508 16788
rect 21732 16736 21784 16788
rect 18880 16668 18932 16720
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 19248 16600 19300 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 17684 16532 17736 16584
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 13360 16464 13412 16516
rect 16028 16507 16080 16516
rect 16028 16473 16037 16507
rect 16037 16473 16071 16507
rect 16071 16473 16080 16507
rect 16028 16464 16080 16473
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 17868 16396 17920 16448
rect 18972 16396 19024 16448
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 22008 16600 22060 16652
rect 22192 16643 22244 16652
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 27896 16736 27948 16788
rect 29828 16736 29880 16788
rect 31024 16736 31076 16788
rect 31668 16779 31720 16788
rect 31668 16745 31677 16779
rect 31677 16745 31711 16779
rect 31711 16745 31720 16779
rect 31668 16736 31720 16745
rect 32956 16736 33008 16788
rect 29276 16600 29328 16652
rect 19892 16532 19944 16584
rect 22560 16575 22612 16584
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 23020 16532 23072 16584
rect 23296 16464 23348 16516
rect 24676 16575 24728 16584
rect 24676 16541 24685 16575
rect 24685 16541 24719 16575
rect 24719 16541 24728 16575
rect 24676 16532 24728 16541
rect 26056 16507 26108 16516
rect 26056 16473 26065 16507
rect 26065 16473 26099 16507
rect 26099 16473 26108 16507
rect 26056 16464 26108 16473
rect 29276 16464 29328 16516
rect 20720 16439 20772 16448
rect 20720 16405 20729 16439
rect 20729 16405 20763 16439
rect 20763 16405 20772 16439
rect 20720 16396 20772 16405
rect 22468 16396 22520 16448
rect 25412 16396 25464 16448
rect 26148 16439 26200 16448
rect 26148 16405 26157 16439
rect 26157 16405 26191 16439
rect 26191 16405 26200 16439
rect 26148 16396 26200 16405
rect 27068 16396 27120 16448
rect 30104 16575 30156 16584
rect 30104 16541 30139 16575
rect 30139 16541 30156 16575
rect 30104 16532 30156 16541
rect 30564 16532 30616 16584
rect 31024 16643 31076 16652
rect 31024 16609 31034 16643
rect 31034 16609 31068 16643
rect 31068 16609 31076 16643
rect 31024 16600 31076 16609
rect 31576 16600 31628 16652
rect 33232 16711 33284 16720
rect 33232 16677 33241 16711
rect 33241 16677 33275 16711
rect 33275 16677 33284 16711
rect 33232 16668 33284 16677
rect 30012 16507 30064 16516
rect 30012 16473 30021 16507
rect 30021 16473 30055 16507
rect 30055 16473 30064 16507
rect 30012 16464 30064 16473
rect 30472 16464 30524 16516
rect 32128 16464 32180 16516
rect 33692 16532 33744 16584
rect 31024 16396 31076 16448
rect 31116 16396 31168 16448
rect 31392 16396 31444 16448
rect 32404 16439 32456 16448
rect 32404 16405 32413 16439
rect 32413 16405 32447 16439
rect 32447 16405 32456 16439
rect 32404 16396 32456 16405
rect 32956 16507 33008 16516
rect 32956 16473 32965 16507
rect 32965 16473 32999 16507
rect 32999 16473 33008 16507
rect 32956 16464 33008 16473
rect 33508 16439 33560 16448
rect 33508 16405 33517 16439
rect 33517 16405 33551 16439
rect 33551 16405 33560 16439
rect 33508 16396 33560 16405
rect 33692 16439 33744 16448
rect 33692 16405 33719 16439
rect 33719 16405 33744 16439
rect 33692 16396 33744 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 10784 16192 10836 16244
rect 8300 16124 8352 16176
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 10048 16056 10100 16108
rect 11152 16124 11204 16176
rect 11520 16056 11572 16108
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 12072 16124 12124 16176
rect 14280 16192 14332 16244
rect 14648 16192 14700 16244
rect 16028 16192 16080 16244
rect 18972 16235 19024 16244
rect 18972 16201 18981 16235
rect 18981 16201 19015 16235
rect 19015 16201 19024 16235
rect 18972 16192 19024 16201
rect 19616 16192 19668 16244
rect 9128 15920 9180 15972
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 17868 16124 17920 16176
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15108 16056 15160 16108
rect 16120 16056 16172 16108
rect 18420 16056 18472 16108
rect 20720 16124 20772 16176
rect 22008 16124 22060 16176
rect 23664 16167 23716 16176
rect 23664 16133 23673 16167
rect 23673 16133 23707 16167
rect 23707 16133 23716 16167
rect 23664 16124 23716 16133
rect 25412 16124 25464 16176
rect 23756 16056 23808 16108
rect 26424 16056 26476 16108
rect 17040 15988 17092 16040
rect 18788 15963 18840 15972
rect 18788 15929 18797 15963
rect 18797 15929 18831 15963
rect 18831 15929 18840 15963
rect 18788 15920 18840 15929
rect 19800 15920 19852 15972
rect 19892 15920 19944 15972
rect 22560 15920 22612 15972
rect 9864 15852 9916 15904
rect 9956 15852 10008 15904
rect 11980 15895 12032 15904
rect 11980 15861 11989 15895
rect 11989 15861 12023 15895
rect 12023 15861 12032 15895
rect 11980 15852 12032 15861
rect 12164 15852 12216 15904
rect 14096 15852 14148 15904
rect 20076 15895 20128 15904
rect 20076 15861 20085 15895
rect 20085 15861 20119 15895
rect 20119 15861 20128 15895
rect 20076 15852 20128 15861
rect 21548 15852 21600 15904
rect 23940 15852 23992 15904
rect 24860 15895 24912 15904
rect 24860 15861 24869 15895
rect 24869 15861 24903 15895
rect 24903 15861 24912 15895
rect 24860 15852 24912 15861
rect 25872 15988 25924 16040
rect 29920 16192 29972 16244
rect 32128 16235 32180 16244
rect 32128 16201 32137 16235
rect 32137 16201 32171 16235
rect 32171 16201 32180 16235
rect 32128 16192 32180 16201
rect 27252 16099 27304 16108
rect 27252 16065 27261 16099
rect 27261 16065 27295 16099
rect 27295 16065 27304 16099
rect 27252 16056 27304 16065
rect 30840 16124 30892 16176
rect 30656 16056 30708 16108
rect 31116 16056 31168 16108
rect 31300 16056 31352 16108
rect 32956 16192 33008 16244
rect 33232 16192 33284 16244
rect 32404 16056 32456 16108
rect 29368 15988 29420 16040
rect 29920 15988 29972 16040
rect 31392 16031 31444 16040
rect 31392 15997 31401 16031
rect 31401 15997 31435 16031
rect 31435 15997 31444 16031
rect 31392 15988 31444 15997
rect 31484 16031 31536 16040
rect 31484 15997 31493 16031
rect 31493 15997 31527 16031
rect 31527 15997 31536 16031
rect 31484 15988 31536 15997
rect 32312 15988 32364 16040
rect 25504 15852 25556 15904
rect 27988 15963 28040 15972
rect 27988 15929 27997 15963
rect 27997 15929 28031 15963
rect 28031 15929 28040 15963
rect 37280 16056 37332 16108
rect 27988 15920 28040 15929
rect 28172 15852 28224 15904
rect 29184 15895 29236 15904
rect 29184 15861 29193 15895
rect 29193 15861 29227 15895
rect 29227 15861 29236 15895
rect 29184 15852 29236 15861
rect 29276 15852 29328 15904
rect 31300 15852 31352 15904
rect 33508 15852 33560 15904
rect 33784 15852 33836 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8024 15648 8076 15700
rect 10416 15648 10468 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 11152 15580 11204 15632
rect 14924 15648 14976 15700
rect 29184 15648 29236 15700
rect 29276 15648 29328 15700
rect 35440 15648 35492 15700
rect 10692 15555 10744 15564
rect 10692 15521 10701 15555
rect 10701 15521 10735 15555
rect 10735 15521 10744 15555
rect 10692 15512 10744 15521
rect 11980 15512 12032 15564
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 9956 15444 10008 15496
rect 2780 15376 2832 15428
rect 11520 15444 11572 15496
rect 12164 15444 12216 15496
rect 28172 15580 28224 15632
rect 28540 15623 28592 15632
rect 28540 15589 28549 15623
rect 28549 15589 28583 15623
rect 28583 15589 28592 15623
rect 28540 15580 28592 15589
rect 13728 15512 13780 15564
rect 11980 15376 12032 15428
rect 13820 15444 13872 15496
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 17132 15512 17184 15564
rect 20076 15512 20128 15564
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 16948 15444 17000 15496
rect 20628 15512 20680 15564
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 22100 15512 22152 15564
rect 23756 15555 23808 15564
rect 23756 15521 23765 15555
rect 23765 15521 23799 15555
rect 23799 15521 23808 15555
rect 23756 15512 23808 15521
rect 10048 15308 10100 15360
rect 11152 15351 11204 15360
rect 11152 15317 11161 15351
rect 11161 15317 11195 15351
rect 11195 15317 11204 15351
rect 11152 15308 11204 15317
rect 12072 15308 12124 15360
rect 13912 15351 13964 15360
rect 13912 15317 13921 15351
rect 13921 15317 13955 15351
rect 13955 15317 13964 15351
rect 13912 15308 13964 15317
rect 14924 15351 14976 15360
rect 14924 15317 14933 15351
rect 14933 15317 14967 15351
rect 14967 15317 14976 15351
rect 14924 15308 14976 15317
rect 17776 15308 17828 15360
rect 21272 15376 21324 15428
rect 23572 15444 23624 15496
rect 23848 15444 23900 15496
rect 24400 15444 24452 15496
rect 27988 15444 28040 15496
rect 30472 15623 30524 15632
rect 30472 15589 30481 15623
rect 30481 15589 30515 15623
rect 30515 15589 30524 15623
rect 30472 15580 30524 15589
rect 31024 15623 31076 15632
rect 31024 15589 31033 15623
rect 31033 15589 31067 15623
rect 31067 15589 31076 15623
rect 31024 15580 31076 15589
rect 32312 15580 32364 15632
rect 33784 15580 33836 15632
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 21548 15308 21600 15360
rect 25596 15308 25648 15360
rect 27252 15376 27304 15428
rect 28264 15419 28316 15428
rect 28264 15385 28273 15419
rect 28273 15385 28307 15419
rect 28307 15385 28316 15419
rect 28264 15376 28316 15385
rect 27528 15308 27580 15360
rect 29460 15376 29512 15428
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 29000 15308 29052 15360
rect 29920 15351 29972 15360
rect 29920 15317 29929 15351
rect 29929 15317 29963 15351
rect 29963 15317 29972 15351
rect 29920 15308 29972 15317
rect 30104 15351 30156 15360
rect 30104 15317 30113 15351
rect 30113 15317 30147 15351
rect 30147 15317 30156 15351
rect 30104 15308 30156 15317
rect 31576 15376 31628 15428
rect 31484 15308 31536 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 18420 15104 18472 15156
rect 21824 15104 21876 15156
rect 25872 15147 25924 15156
rect 25872 15113 25881 15147
rect 25881 15113 25915 15147
rect 25915 15113 25924 15147
rect 25872 15104 25924 15113
rect 26424 15147 26476 15156
rect 26424 15113 26433 15147
rect 26433 15113 26467 15147
rect 26467 15113 26476 15147
rect 26424 15104 26476 15113
rect 11152 15036 11204 15088
rect 18604 15036 18656 15088
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 13912 14900 13964 14952
rect 13728 14875 13780 14884
rect 13728 14841 13737 14875
rect 13737 14841 13771 14875
rect 13771 14841 13780 14875
rect 13728 14832 13780 14841
rect 14464 14968 14516 15020
rect 16948 14968 17000 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 22100 15036 22152 15088
rect 23572 15036 23624 15088
rect 27252 15104 27304 15156
rect 15016 14900 15068 14952
rect 16672 14943 16724 14952
rect 16672 14909 16681 14943
rect 16681 14909 16715 14943
rect 16715 14909 16724 14943
rect 16672 14900 16724 14909
rect 17132 14943 17184 14952
rect 17132 14909 17141 14943
rect 17141 14909 17175 14943
rect 17175 14909 17184 14943
rect 17132 14900 17184 14909
rect 17592 14900 17644 14952
rect 17776 14943 17828 14952
rect 17776 14909 17785 14943
rect 17785 14909 17819 14943
rect 17819 14909 17828 14943
rect 17776 14900 17828 14909
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 17960 14943 18012 14952
rect 17960 14909 17969 14943
rect 17969 14909 18003 14943
rect 18003 14909 18012 14943
rect 17960 14900 18012 14909
rect 19708 14900 19760 14952
rect 19156 14832 19208 14884
rect 12992 14764 13044 14816
rect 14096 14764 14148 14816
rect 19616 14764 19668 14816
rect 20536 14968 20588 15020
rect 21548 15011 21600 15020
rect 21548 14977 21557 15011
rect 21557 14977 21591 15011
rect 21591 14977 21600 15011
rect 21548 14968 21600 14977
rect 25596 14968 25648 15020
rect 23572 14900 23624 14952
rect 23204 14832 23256 14884
rect 20720 14764 20772 14816
rect 21088 14807 21140 14816
rect 21088 14773 21097 14807
rect 21097 14773 21131 14807
rect 21131 14773 21140 14807
rect 21088 14764 21140 14773
rect 21364 14764 21416 14816
rect 22284 14764 22336 14816
rect 23756 14807 23808 14816
rect 23756 14773 23765 14807
rect 23765 14773 23799 14807
rect 23799 14773 23808 14807
rect 23756 14764 23808 14773
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 30104 15104 30156 15156
rect 27712 15036 27764 15088
rect 28540 15036 28592 15088
rect 30012 15036 30064 15088
rect 27528 14943 27580 14952
rect 27528 14909 27537 14943
rect 27537 14909 27571 14943
rect 27571 14909 27580 14943
rect 27528 14900 27580 14909
rect 29000 15011 29052 15020
rect 29000 14977 29009 15011
rect 29009 14977 29043 15011
rect 29043 14977 29052 15011
rect 29000 14968 29052 14977
rect 29920 15011 29972 15020
rect 29920 14977 29929 15011
rect 29929 14977 29963 15011
rect 29963 14977 29972 15011
rect 29920 14968 29972 14977
rect 28724 14900 28776 14952
rect 29644 14900 29696 14952
rect 30656 14900 30708 14952
rect 28264 14875 28316 14884
rect 28264 14841 28273 14875
rect 28273 14841 28307 14875
rect 28307 14841 28316 14875
rect 28264 14832 28316 14841
rect 28356 14832 28408 14884
rect 28908 14832 28960 14884
rect 28816 14807 28868 14816
rect 28816 14773 28825 14807
rect 28825 14773 28859 14807
rect 28859 14773 28868 14807
rect 28816 14764 28868 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 10048 14424 10100 14476
rect 10324 14424 10376 14476
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 14096 14560 14148 14612
rect 16672 14560 16724 14612
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 17960 14560 18012 14612
rect 19984 14560 20036 14612
rect 20076 14603 20128 14612
rect 20076 14569 20085 14603
rect 20085 14569 20119 14603
rect 20119 14569 20128 14603
rect 20076 14560 20128 14569
rect 21088 14560 21140 14612
rect 13728 14492 13780 14544
rect 14924 14492 14976 14544
rect 15200 14492 15252 14544
rect 8300 14220 8352 14272
rect 11152 14356 11204 14408
rect 12624 14356 12676 14408
rect 13176 14399 13228 14408
rect 13176 14365 13185 14399
rect 13185 14365 13219 14399
rect 13219 14365 13228 14399
rect 13176 14356 13228 14365
rect 13912 14356 13964 14408
rect 15200 14399 15252 14408
rect 15200 14365 15209 14399
rect 15209 14365 15243 14399
rect 15243 14365 15252 14399
rect 15200 14356 15252 14365
rect 15752 14356 15804 14408
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 19340 14492 19392 14544
rect 16948 14467 17000 14476
rect 16948 14433 16957 14467
rect 16957 14433 16991 14467
rect 16991 14433 17000 14467
rect 16948 14424 17000 14433
rect 17960 14424 18012 14476
rect 17132 14356 17184 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 9680 14220 9732 14272
rect 12900 14331 12952 14340
rect 12900 14297 12909 14331
rect 12909 14297 12943 14331
rect 12943 14297 12952 14331
rect 12900 14288 12952 14297
rect 14832 14288 14884 14340
rect 12992 14220 13044 14272
rect 14556 14263 14608 14272
rect 14556 14229 14565 14263
rect 14565 14229 14599 14263
rect 14599 14229 14608 14263
rect 14556 14220 14608 14229
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 17316 14331 17368 14340
rect 17316 14297 17325 14331
rect 17325 14297 17359 14331
rect 17359 14297 17368 14331
rect 17316 14288 17368 14297
rect 17592 14331 17644 14340
rect 17592 14297 17601 14331
rect 17601 14297 17635 14331
rect 17635 14297 17644 14331
rect 17592 14288 17644 14297
rect 17684 14288 17736 14340
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 19064 14399 19116 14408
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 19156 14356 19208 14408
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 18788 14220 18840 14272
rect 20628 14220 20680 14272
rect 22468 14603 22520 14612
rect 22468 14569 22477 14603
rect 22477 14569 22511 14603
rect 22511 14569 22520 14603
rect 22468 14560 22520 14569
rect 21548 14424 21600 14476
rect 22284 14356 22336 14408
rect 22376 14356 22428 14408
rect 26148 14560 26200 14612
rect 26884 14560 26936 14612
rect 27344 14560 27396 14612
rect 28816 14560 28868 14612
rect 29092 14560 29144 14612
rect 29184 14560 29236 14612
rect 29736 14560 29788 14612
rect 31116 14603 31168 14612
rect 31116 14569 31125 14603
rect 31125 14569 31159 14603
rect 31159 14569 31168 14603
rect 31116 14560 31168 14569
rect 31576 14603 31628 14612
rect 31576 14569 31585 14603
rect 31585 14569 31619 14603
rect 31619 14569 31628 14603
rect 31576 14560 31628 14569
rect 28724 14492 28776 14544
rect 23296 14424 23348 14476
rect 23480 14424 23532 14476
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 24860 14356 24912 14408
rect 22100 14288 22152 14340
rect 22744 14331 22796 14340
rect 22744 14297 22753 14331
rect 22753 14297 22787 14331
rect 22787 14297 22796 14331
rect 22744 14288 22796 14297
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 28632 14424 28684 14476
rect 26884 14399 26936 14408
rect 26884 14365 26893 14399
rect 26893 14365 26927 14399
rect 26927 14365 26936 14399
rect 26884 14356 26936 14365
rect 27068 14399 27120 14408
rect 27068 14365 27077 14399
rect 27077 14365 27111 14399
rect 27111 14365 27120 14399
rect 27068 14356 27120 14365
rect 22192 14220 22244 14272
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 23756 14263 23808 14272
rect 23756 14229 23765 14263
rect 23765 14229 23799 14263
rect 23799 14229 23808 14263
rect 23756 14220 23808 14229
rect 27252 14220 27304 14272
rect 27528 14220 27580 14272
rect 27620 14220 27672 14272
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 28724 14288 28776 14340
rect 28908 14220 28960 14272
rect 30840 14356 30892 14408
rect 32128 14492 32180 14544
rect 32496 14467 32548 14476
rect 32496 14433 32505 14467
rect 32505 14433 32539 14467
rect 32539 14433 32548 14467
rect 32496 14424 32548 14433
rect 31852 14356 31904 14408
rect 32036 14356 32088 14408
rect 31576 14288 31628 14340
rect 30380 14220 30432 14272
rect 31392 14220 31444 14272
rect 35624 14356 35676 14408
rect 33048 14263 33100 14272
rect 33048 14229 33057 14263
rect 33057 14229 33091 14263
rect 33091 14229 33100 14263
rect 33048 14220 33100 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 7748 14016 7800 14068
rect 8944 14016 8996 14068
rect 9680 14016 9732 14068
rect 11520 14016 11572 14068
rect 12624 14016 12676 14068
rect 13820 14016 13872 14068
rect 14096 14016 14148 14068
rect 8300 13948 8352 14000
rect 8668 13948 8720 14000
rect 9864 13880 9916 13932
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 11888 13880 11940 13932
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 14924 14016 14976 14068
rect 15660 14016 15712 14068
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 18420 14016 18472 14068
rect 19064 14016 19116 14068
rect 19616 14016 19668 14068
rect 19708 14016 19760 14068
rect 23296 14016 23348 14068
rect 23572 14059 23624 14068
rect 23572 14025 23581 14059
rect 23581 14025 23615 14059
rect 23615 14025 23624 14059
rect 23572 14016 23624 14025
rect 23664 14016 23716 14068
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 27252 14016 27304 14068
rect 14464 13948 14516 14000
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 13268 13676 13320 13728
rect 14556 13812 14608 13864
rect 14832 13855 14884 13864
rect 14832 13821 14841 13855
rect 14841 13821 14875 13855
rect 14875 13821 14884 13855
rect 14832 13812 14884 13821
rect 17316 13948 17368 14000
rect 17776 13923 17828 13932
rect 17776 13889 17785 13923
rect 17785 13889 17819 13923
rect 17819 13889 17828 13923
rect 17776 13880 17828 13889
rect 18052 13880 18104 13932
rect 18788 13923 18840 13932
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 20812 13855 20864 13864
rect 20812 13821 20821 13855
rect 20821 13821 20855 13855
rect 20855 13821 20864 13855
rect 20812 13812 20864 13821
rect 21272 13812 21324 13864
rect 23020 13880 23072 13932
rect 23112 13923 23164 13932
rect 23112 13889 23121 13923
rect 23121 13889 23155 13923
rect 23155 13889 23164 13923
rect 23112 13880 23164 13889
rect 14556 13719 14608 13728
rect 14556 13685 14565 13719
rect 14565 13685 14599 13719
rect 14599 13685 14608 13719
rect 14556 13676 14608 13685
rect 14832 13676 14884 13728
rect 20996 13719 21048 13728
rect 20996 13685 21005 13719
rect 21005 13685 21039 13719
rect 21039 13685 21048 13719
rect 20996 13676 21048 13685
rect 27528 13948 27580 14000
rect 23756 13880 23808 13932
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 27252 13923 27304 13932
rect 27252 13889 27261 13923
rect 27261 13889 27295 13923
rect 27295 13889 27304 13923
rect 27252 13880 27304 13889
rect 27620 13923 27672 13932
rect 27620 13889 27629 13923
rect 27629 13889 27663 13923
rect 27663 13889 27672 13923
rect 27620 13880 27672 13889
rect 27436 13812 27488 13864
rect 29552 13948 29604 14000
rect 29736 13948 29788 14000
rect 31484 14059 31536 14068
rect 31484 14025 31493 14059
rect 31493 14025 31527 14059
rect 31527 14025 31536 14059
rect 31484 14016 31536 14025
rect 31576 14016 31628 14068
rect 32036 14016 32088 14068
rect 33048 14016 33100 14068
rect 25596 13744 25648 13796
rect 26976 13744 27028 13796
rect 28448 13880 28500 13932
rect 28632 13812 28684 13864
rect 29276 13880 29328 13932
rect 30564 13880 30616 13932
rect 31208 13923 31260 13932
rect 31208 13889 31217 13923
rect 31217 13889 31251 13923
rect 31251 13889 31260 13923
rect 31208 13880 31260 13889
rect 31392 13923 31444 13932
rect 31392 13889 31401 13923
rect 31401 13889 31435 13923
rect 31435 13889 31444 13923
rect 31392 13880 31444 13889
rect 32036 13880 32088 13932
rect 32220 13880 32272 13932
rect 32496 13923 32548 13932
rect 32496 13889 32505 13923
rect 32505 13889 32539 13923
rect 32539 13889 32548 13923
rect 32496 13880 32548 13889
rect 24952 13719 25004 13728
rect 24952 13685 24961 13719
rect 24961 13685 24995 13719
rect 24995 13685 25004 13719
rect 24952 13676 25004 13685
rect 25504 13719 25556 13728
rect 25504 13685 25513 13719
rect 25513 13685 25547 13719
rect 25547 13685 25556 13719
rect 25504 13676 25556 13685
rect 27620 13676 27672 13728
rect 27896 13676 27948 13728
rect 30472 13676 30524 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4068 13472 4120 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9956 13472 10008 13524
rect 13728 13472 13780 13524
rect 13820 13472 13872 13524
rect 14004 13472 14056 13524
rect 14464 13472 14516 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 11888 13404 11940 13456
rect 12992 13404 13044 13456
rect 13360 13447 13412 13456
rect 13360 13413 13369 13447
rect 13369 13413 13403 13447
rect 13403 13413 13412 13447
rect 13360 13404 13412 13413
rect 22376 13472 22428 13524
rect 23112 13472 23164 13524
rect 9680 13268 9732 13320
rect 9128 13200 9180 13252
rect 9864 13268 9916 13320
rect 10324 13268 10376 13320
rect 12992 13268 13044 13320
rect 13268 13268 13320 13320
rect 12256 13243 12308 13252
rect 12256 13209 12265 13243
rect 12265 13209 12299 13243
rect 12299 13209 12308 13243
rect 12256 13200 12308 13209
rect 12900 13200 12952 13252
rect 13728 13311 13780 13320
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 13452 13200 13504 13252
rect 18052 13379 18104 13388
rect 18052 13345 18061 13379
rect 18061 13345 18095 13379
rect 18095 13345 18104 13379
rect 18052 13336 18104 13345
rect 21088 13336 21140 13388
rect 27252 13472 27304 13524
rect 27620 13472 27672 13524
rect 27988 13472 28040 13524
rect 30840 13472 30892 13524
rect 31208 13472 31260 13524
rect 31852 13515 31904 13524
rect 31852 13481 31861 13515
rect 31861 13481 31895 13515
rect 31895 13481 31904 13515
rect 31852 13472 31904 13481
rect 24308 13404 24360 13456
rect 17224 13268 17276 13320
rect 17776 13268 17828 13320
rect 24400 13336 24452 13388
rect 21272 13268 21324 13320
rect 22100 13268 22152 13320
rect 22560 13268 22612 13320
rect 22744 13268 22796 13320
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 23112 13311 23164 13320
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 19708 13200 19760 13252
rect 24952 13336 25004 13388
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 27712 13268 27764 13320
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 27896 13268 27948 13320
rect 28724 13268 28776 13320
rect 29552 13311 29604 13320
rect 29552 13277 29561 13311
rect 29561 13277 29595 13311
rect 29595 13277 29604 13311
rect 29552 13268 29604 13277
rect 32220 13379 32272 13388
rect 32220 13345 32229 13379
rect 32229 13345 32263 13379
rect 32263 13345 32272 13379
rect 32220 13336 32272 13345
rect 31944 13268 31996 13320
rect 28080 13200 28132 13252
rect 29828 13243 29880 13252
rect 29828 13209 29837 13243
rect 29837 13209 29871 13243
rect 29871 13209 29880 13243
rect 29828 13200 29880 13209
rect 30380 13200 30432 13252
rect 14464 13132 14516 13184
rect 25136 13175 25188 13184
rect 25136 13141 25145 13175
rect 25145 13141 25179 13175
rect 25179 13141 25188 13175
rect 25136 13132 25188 13141
rect 25688 13175 25740 13184
rect 25688 13141 25697 13175
rect 25697 13141 25731 13175
rect 25731 13141 25740 13175
rect 25688 13132 25740 13141
rect 27620 13132 27672 13184
rect 27896 13132 27948 13184
rect 30104 13132 30156 13184
rect 31760 13132 31812 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 11980 12928 12032 12980
rect 12348 12928 12400 12980
rect 12532 12928 12584 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13360 12928 13412 12980
rect 14556 12928 14608 12980
rect 17132 12928 17184 12980
rect 20996 12928 21048 12980
rect 22560 12928 22612 12980
rect 22928 12928 22980 12980
rect 24768 12971 24820 12980
rect 24768 12937 24777 12971
rect 24777 12937 24811 12971
rect 24811 12937 24820 12971
rect 24768 12928 24820 12937
rect 24952 12928 25004 12980
rect 25596 12928 25648 12980
rect 27712 12971 27764 12980
rect 27712 12937 27721 12971
rect 27721 12937 27755 12971
rect 27755 12937 27764 12971
rect 27712 12928 27764 12937
rect 27988 12928 28040 12980
rect 29276 12971 29328 12980
rect 29276 12937 29285 12971
rect 29285 12937 29319 12971
rect 29319 12937 29328 12971
rect 29276 12928 29328 12937
rect 29828 12928 29880 12980
rect 30472 12928 30524 12980
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12164 12724 12216 12776
rect 12808 12792 12860 12844
rect 16672 12792 16724 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18236 12792 18288 12844
rect 19800 12792 19852 12844
rect 20536 12792 20588 12844
rect 20812 12835 20864 12844
rect 20812 12801 20821 12835
rect 20821 12801 20855 12835
rect 20855 12801 20864 12835
rect 20812 12792 20864 12801
rect 24308 12860 24360 12912
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 17224 12699 17276 12708
rect 17224 12665 17233 12699
rect 17233 12665 17267 12699
rect 17267 12665 17276 12699
rect 17224 12656 17276 12665
rect 19064 12724 19116 12776
rect 18420 12656 18472 12708
rect 19800 12656 19852 12708
rect 20812 12656 20864 12708
rect 21364 12835 21416 12844
rect 21364 12801 21373 12835
rect 21373 12801 21407 12835
rect 21407 12801 21416 12835
rect 21364 12792 21416 12801
rect 8852 12588 8904 12640
rect 12440 12588 12492 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 20996 12631 21048 12640
rect 20996 12597 21005 12631
rect 21005 12597 21039 12631
rect 21039 12597 21048 12631
rect 20996 12588 21048 12597
rect 21088 12588 21140 12640
rect 22744 12792 22796 12844
rect 24768 12835 24820 12844
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 25228 12860 25280 12912
rect 25688 12903 25740 12912
rect 25688 12869 25697 12903
rect 25697 12869 25731 12903
rect 25731 12869 25740 12903
rect 25688 12860 25740 12869
rect 27436 12860 27488 12912
rect 30104 12903 30156 12912
rect 30104 12869 30113 12903
rect 30113 12869 30147 12903
rect 30147 12869 30156 12903
rect 30104 12860 30156 12869
rect 31944 12860 31996 12912
rect 32036 12860 32088 12912
rect 25136 12792 25188 12844
rect 25504 12792 25556 12844
rect 25964 12724 26016 12776
rect 27528 12835 27580 12844
rect 27528 12801 27537 12835
rect 27537 12801 27571 12835
rect 27571 12801 27580 12835
rect 27528 12792 27580 12801
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 28172 12835 28224 12844
rect 28172 12801 28181 12835
rect 28181 12801 28215 12835
rect 28215 12801 28224 12835
rect 28172 12792 28224 12801
rect 27620 12724 27672 12776
rect 27804 12724 27856 12776
rect 28264 12724 28316 12776
rect 25872 12699 25924 12708
rect 25872 12665 25881 12699
rect 25881 12665 25915 12699
rect 25915 12665 25924 12699
rect 25872 12656 25924 12665
rect 27896 12699 27948 12708
rect 27896 12665 27905 12699
rect 27905 12665 27939 12699
rect 27939 12665 27948 12699
rect 29460 12724 29512 12776
rect 30840 12835 30892 12844
rect 30840 12801 30849 12835
rect 30849 12801 30883 12835
rect 30883 12801 30892 12835
rect 30840 12792 30892 12801
rect 32128 12835 32180 12844
rect 32128 12801 32137 12835
rect 32137 12801 32171 12835
rect 32171 12801 32180 12835
rect 32128 12792 32180 12801
rect 32588 12792 32640 12844
rect 30196 12767 30248 12776
rect 30196 12733 30205 12767
rect 30205 12733 30239 12767
rect 30239 12733 30248 12767
rect 30196 12724 30248 12733
rect 30564 12724 30616 12776
rect 27896 12656 27948 12665
rect 25044 12631 25096 12640
rect 25044 12597 25053 12631
rect 25053 12597 25087 12631
rect 25087 12597 25096 12631
rect 25044 12588 25096 12597
rect 31852 12588 31904 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12256 12384 12308 12436
rect 13728 12384 13780 12436
rect 16856 12384 16908 12436
rect 13452 12316 13504 12368
rect 11796 12248 11848 12300
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 8852 12180 8904 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9680 12112 9732 12164
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 13636 12180 13688 12232
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 16304 12112 16356 12164
rect 18328 12384 18380 12436
rect 18420 12384 18472 12436
rect 17132 12112 17184 12164
rect 20720 12384 20772 12436
rect 21364 12384 21416 12436
rect 22744 12384 22796 12436
rect 22928 12384 22980 12436
rect 25504 12384 25556 12436
rect 26056 12384 26108 12436
rect 27160 12384 27212 12436
rect 28816 12384 28868 12436
rect 31392 12384 31444 12436
rect 32128 12384 32180 12436
rect 20996 12248 21048 12300
rect 20536 12223 20588 12232
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 20720 12223 20772 12232
rect 20720 12189 20729 12223
rect 20729 12189 20763 12223
rect 20763 12189 20772 12223
rect 20720 12180 20772 12189
rect 20812 12180 20864 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 22008 12316 22060 12368
rect 22836 12223 22888 12232
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 9864 12044 9916 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 12256 12044 12308 12096
rect 17868 12044 17920 12096
rect 18696 12044 18748 12096
rect 19616 12044 19668 12096
rect 20812 12044 20864 12096
rect 21456 12044 21508 12096
rect 23112 12180 23164 12232
rect 31760 12359 31812 12368
rect 31760 12325 31769 12359
rect 31769 12325 31803 12359
rect 31803 12325 31812 12359
rect 31760 12316 31812 12325
rect 25044 12291 25096 12300
rect 25044 12257 25053 12291
rect 25053 12257 25087 12291
rect 25087 12257 25096 12291
rect 25044 12248 25096 12257
rect 25320 12291 25372 12300
rect 25320 12257 25329 12291
rect 25329 12257 25363 12291
rect 25363 12257 25372 12291
rect 25320 12248 25372 12257
rect 23756 12180 23808 12232
rect 29460 12248 29512 12300
rect 25964 12223 26016 12232
rect 25964 12189 25973 12223
rect 25973 12189 26007 12223
rect 26007 12189 26016 12223
rect 25964 12180 26016 12189
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 28080 12180 28132 12232
rect 25872 12112 25924 12164
rect 27804 12155 27856 12164
rect 27804 12121 27813 12155
rect 27813 12121 27847 12155
rect 27847 12121 27856 12155
rect 27804 12112 27856 12121
rect 23296 12087 23348 12096
rect 23296 12053 23305 12087
rect 23305 12053 23339 12087
rect 23339 12053 23348 12087
rect 23296 12044 23348 12053
rect 25412 12044 25464 12096
rect 25596 12044 25648 12096
rect 27436 12087 27488 12096
rect 27436 12053 27445 12087
rect 27445 12053 27479 12087
rect 27479 12053 27488 12087
rect 27436 12044 27488 12053
rect 31208 12044 31260 12096
rect 31852 12248 31904 12300
rect 32220 12180 32272 12232
rect 32128 12112 32180 12164
rect 34152 12223 34204 12232
rect 34152 12189 34161 12223
rect 34161 12189 34195 12223
rect 34195 12189 34204 12223
rect 34152 12180 34204 12189
rect 34520 12180 34572 12232
rect 31668 12044 31720 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 9680 11840 9732 11892
rect 11796 11840 11848 11892
rect 16304 11883 16356 11892
rect 16304 11849 16313 11883
rect 16313 11849 16347 11883
rect 16347 11849 16356 11883
rect 16304 11840 16356 11849
rect 16672 11883 16724 11892
rect 16672 11849 16681 11883
rect 16681 11849 16715 11883
rect 16715 11849 16724 11883
rect 16672 11840 16724 11849
rect 9128 11636 9180 11688
rect 4068 11568 4120 11620
rect 9864 11704 9916 11756
rect 17132 11815 17184 11824
rect 17132 11781 17141 11815
rect 17141 11781 17175 11815
rect 17175 11781 17184 11815
rect 17132 11772 17184 11781
rect 17868 11772 17920 11824
rect 19708 11815 19760 11824
rect 19708 11781 19717 11815
rect 19717 11781 19751 11815
rect 19751 11781 19760 11815
rect 19708 11772 19760 11781
rect 19800 11815 19852 11824
rect 19800 11781 19809 11815
rect 19809 11781 19843 11815
rect 19843 11781 19852 11815
rect 19800 11772 19852 11781
rect 20720 11840 20772 11892
rect 20904 11840 20956 11892
rect 20996 11883 21048 11892
rect 20996 11849 21021 11883
rect 21021 11849 21048 11883
rect 20996 11840 21048 11849
rect 21180 11883 21232 11892
rect 21180 11849 21189 11883
rect 21189 11849 21223 11883
rect 21223 11849 21232 11883
rect 21180 11840 21232 11849
rect 26056 11840 26108 11892
rect 26148 11840 26200 11892
rect 26608 11840 26660 11892
rect 20812 11815 20864 11824
rect 17408 11704 17460 11756
rect 19616 11747 19668 11756
rect 19616 11713 19625 11747
rect 19625 11713 19659 11747
rect 19659 11713 19668 11747
rect 19616 11704 19668 11713
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20812 11781 20821 11815
rect 20821 11781 20855 11815
rect 20855 11781 20864 11815
rect 20812 11772 20864 11781
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 24860 11704 24912 11756
rect 18972 11500 19024 11552
rect 25688 11704 25740 11756
rect 26148 11704 26200 11756
rect 31668 11840 31720 11892
rect 32128 11815 32180 11824
rect 32128 11781 32137 11815
rect 32137 11781 32171 11815
rect 32171 11781 32180 11815
rect 32128 11772 32180 11781
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 31852 11704 31904 11756
rect 25412 11568 25464 11620
rect 27528 11611 27580 11620
rect 27528 11577 27537 11611
rect 27537 11577 27571 11611
rect 27571 11577 27580 11611
rect 27528 11568 27580 11577
rect 31392 11679 31444 11688
rect 31392 11645 31401 11679
rect 31401 11645 31435 11679
rect 31435 11645 31444 11679
rect 31392 11636 31444 11645
rect 21456 11500 21508 11552
rect 31944 11568 31996 11620
rect 32588 11883 32640 11892
rect 32588 11849 32597 11883
rect 32597 11849 32631 11883
rect 32631 11849 32640 11883
rect 32588 11840 32640 11849
rect 28264 11500 28316 11552
rect 28632 11500 28684 11552
rect 28908 11543 28960 11552
rect 28908 11509 28917 11543
rect 28917 11509 28951 11543
rect 28951 11509 28960 11543
rect 28908 11500 28960 11509
rect 30472 11500 30524 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12348 11228 12400 11280
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 10692 11092 10744 11144
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 11980 11092 12032 11144
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 9128 11024 9180 11076
rect 10784 11024 10836 11076
rect 14372 11203 14424 11212
rect 14372 11169 14381 11203
rect 14381 11169 14415 11203
rect 14415 11169 14424 11203
rect 14372 11160 14424 11169
rect 14832 11160 14884 11212
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 16120 11160 16172 11212
rect 17408 11160 17460 11212
rect 13544 11092 13596 11101
rect 14004 10956 14056 11008
rect 14280 10956 14332 11008
rect 14832 10956 14884 11008
rect 15568 11092 15620 11144
rect 17224 11092 17276 11144
rect 17868 11024 17920 11076
rect 18420 11092 18472 11144
rect 23296 11296 23348 11348
rect 23388 11296 23440 11348
rect 24308 11296 24360 11348
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 23388 11160 23440 11212
rect 22836 11024 22888 11076
rect 23388 11067 23440 11076
rect 23388 11033 23397 11067
rect 23397 11033 23431 11067
rect 23431 11033 23440 11067
rect 23388 11024 23440 11033
rect 15384 10999 15436 11008
rect 15384 10965 15393 10999
rect 15393 10965 15427 10999
rect 15427 10965 15436 10999
rect 15384 10956 15436 10965
rect 18052 10956 18104 11008
rect 18512 10956 18564 11008
rect 22284 10999 22336 11008
rect 22284 10965 22293 10999
rect 22293 10965 22327 10999
rect 22327 10965 22336 10999
rect 22284 10956 22336 10965
rect 22744 10999 22796 11008
rect 22744 10965 22753 10999
rect 22753 10965 22787 10999
rect 22787 10965 22796 10999
rect 25688 11296 25740 11348
rect 25872 11339 25924 11348
rect 25872 11305 25881 11339
rect 25881 11305 25915 11339
rect 25915 11305 25924 11339
rect 25872 11296 25924 11305
rect 28724 11339 28776 11348
rect 28724 11305 28733 11339
rect 28733 11305 28767 11339
rect 28767 11305 28776 11339
rect 28724 11296 28776 11305
rect 28908 11296 28960 11348
rect 32220 11296 32272 11348
rect 38200 11296 38252 11348
rect 24768 11203 24820 11212
rect 24768 11169 24777 11203
rect 24777 11169 24811 11203
rect 24811 11169 24820 11203
rect 24768 11160 24820 11169
rect 25228 11203 25280 11212
rect 25228 11169 25237 11203
rect 25237 11169 25271 11203
rect 25271 11169 25280 11203
rect 25228 11160 25280 11169
rect 26976 11160 27028 11212
rect 24676 11092 24728 11144
rect 25228 11024 25280 11076
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 28080 11024 28132 11076
rect 28632 11092 28684 11144
rect 30472 11135 30524 11144
rect 30472 11101 30481 11135
rect 30481 11101 30515 11135
rect 30515 11101 30524 11135
rect 30472 11092 30524 11101
rect 22744 10956 22796 10965
rect 28264 10956 28316 11008
rect 28356 10956 28408 11008
rect 32128 11024 32180 11076
rect 28816 10956 28868 11008
rect 28908 10999 28960 11008
rect 28908 10965 28917 10999
rect 28917 10965 28951 10999
rect 28951 10965 28960 10999
rect 28908 10956 28960 10965
rect 30932 10956 30984 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 10508 10616 10560 10668
rect 12440 10684 12492 10736
rect 10232 10591 10284 10600
rect 10232 10557 10241 10591
rect 10241 10557 10275 10591
rect 10275 10557 10284 10591
rect 10232 10548 10284 10557
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 10784 10548 10836 10600
rect 12348 10591 12400 10600
rect 12348 10557 12357 10591
rect 12357 10557 12391 10591
rect 12391 10557 12400 10591
rect 12348 10548 12400 10557
rect 13544 10548 13596 10600
rect 14280 10616 14332 10668
rect 14372 10616 14424 10668
rect 12532 10480 12584 10532
rect 9772 10412 9824 10464
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 13912 10480 13964 10532
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 15384 10752 15436 10804
rect 16120 10616 16172 10668
rect 17224 10659 17276 10668
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 24676 10752 24728 10804
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 27436 10752 27488 10804
rect 28172 10752 28224 10804
rect 18052 10684 18104 10736
rect 17868 10616 17920 10668
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 18512 10616 18564 10668
rect 22284 10616 22336 10668
rect 25228 10616 25280 10668
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 25504 10659 25556 10668
rect 25504 10625 25513 10659
rect 25513 10625 25547 10659
rect 25547 10625 25556 10659
rect 25504 10616 25556 10625
rect 26056 10684 26108 10736
rect 26976 10684 27028 10736
rect 28908 10752 28960 10804
rect 15568 10412 15620 10464
rect 22744 10548 22796 10600
rect 17868 10523 17920 10532
rect 17868 10489 17877 10523
rect 17877 10489 17911 10523
rect 17911 10489 17920 10523
rect 17868 10480 17920 10489
rect 18788 10480 18840 10532
rect 23388 10480 23440 10532
rect 24032 10480 24084 10532
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 19892 10412 19944 10464
rect 21640 10412 21692 10464
rect 25412 10412 25464 10464
rect 31392 10752 31444 10804
rect 32128 10795 32180 10804
rect 32128 10761 32137 10795
rect 32137 10761 32171 10795
rect 32171 10761 32180 10795
rect 32128 10752 32180 10761
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 27988 10659 28040 10668
rect 27988 10625 27997 10659
rect 27997 10625 28031 10659
rect 28031 10625 28040 10659
rect 27988 10616 28040 10625
rect 28356 10616 28408 10668
rect 28448 10659 28500 10668
rect 28448 10625 28457 10659
rect 28457 10625 28491 10659
rect 28491 10625 28500 10659
rect 28448 10616 28500 10625
rect 28724 10659 28776 10668
rect 28724 10625 28733 10659
rect 28733 10625 28767 10659
rect 28767 10625 28776 10659
rect 28724 10616 28776 10625
rect 28908 10659 28960 10668
rect 28908 10625 28917 10659
rect 28917 10625 28951 10659
rect 28951 10625 28960 10659
rect 28908 10616 28960 10625
rect 27528 10480 27580 10532
rect 29736 10659 29788 10668
rect 29736 10625 29745 10659
rect 29745 10625 29779 10659
rect 29779 10625 29788 10659
rect 29736 10616 29788 10625
rect 30932 10727 30984 10736
rect 30932 10693 30941 10727
rect 30941 10693 30975 10727
rect 30975 10693 30984 10727
rect 30932 10684 30984 10693
rect 31300 10616 31352 10668
rect 32864 10659 32916 10668
rect 32864 10625 32873 10659
rect 32873 10625 32907 10659
rect 32907 10625 32916 10659
rect 32864 10616 32916 10625
rect 35348 10616 35400 10668
rect 29828 10591 29880 10600
rect 29828 10557 29837 10591
rect 29837 10557 29871 10591
rect 29871 10557 29880 10591
rect 29828 10548 29880 10557
rect 30380 10591 30432 10600
rect 30380 10557 30389 10591
rect 30389 10557 30423 10591
rect 30423 10557 30432 10591
rect 30380 10548 30432 10557
rect 25872 10455 25924 10464
rect 25872 10421 25881 10455
rect 25881 10421 25915 10455
rect 25915 10421 25924 10455
rect 25872 10412 25924 10421
rect 27344 10455 27396 10464
rect 27344 10421 27353 10455
rect 27353 10421 27387 10455
rect 27387 10421 27396 10455
rect 27344 10412 27396 10421
rect 27896 10455 27948 10464
rect 27896 10421 27905 10455
rect 27905 10421 27939 10455
rect 27939 10421 27948 10455
rect 27896 10412 27948 10421
rect 28080 10455 28132 10464
rect 28080 10421 28089 10455
rect 28089 10421 28123 10455
rect 28123 10421 28132 10455
rect 28080 10412 28132 10421
rect 29092 10455 29144 10464
rect 29092 10421 29101 10455
rect 29101 10421 29135 10455
rect 29135 10421 29144 10455
rect 29092 10412 29144 10421
rect 29184 10412 29236 10464
rect 29644 10412 29696 10464
rect 30840 10412 30892 10464
rect 34152 10548 34204 10600
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10508 10208 10560 10260
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 10600 10004 10652 10056
rect 12440 10208 12492 10260
rect 12532 10251 12584 10260
rect 12532 10217 12541 10251
rect 12541 10217 12575 10251
rect 12575 10217 12584 10251
rect 12532 10208 12584 10217
rect 12624 10208 12676 10260
rect 13912 10208 13964 10260
rect 14648 10208 14700 10260
rect 16396 10208 16448 10260
rect 17868 10208 17920 10260
rect 21272 10208 21324 10260
rect 21640 10208 21692 10260
rect 22744 10208 22796 10260
rect 11520 10072 11572 10124
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 13176 10004 13228 10056
rect 9220 9979 9272 9988
rect 9220 9945 9229 9979
rect 9229 9945 9263 9979
rect 9263 9945 9272 9979
rect 9220 9936 9272 9945
rect 14280 9979 14332 9988
rect 14280 9945 14289 9979
rect 14289 9945 14323 9979
rect 14323 9945 14332 9979
rect 14280 9936 14332 9945
rect 16856 10072 16908 10124
rect 17224 10115 17276 10124
rect 17224 10081 17233 10115
rect 17233 10081 17267 10115
rect 17267 10081 17276 10115
rect 17224 10072 17276 10081
rect 16304 10004 16356 10056
rect 16948 10004 17000 10056
rect 17500 10004 17552 10056
rect 17776 10140 17828 10192
rect 17960 10072 18012 10124
rect 18512 10072 18564 10124
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 19984 9936 20036 9988
rect 21824 10072 21876 10124
rect 20996 10047 21048 10056
rect 20996 10013 21004 10047
rect 21004 10013 21038 10047
rect 21038 10013 21048 10047
rect 20996 10004 21048 10013
rect 21088 10047 21140 10056
rect 21088 10013 21097 10047
rect 21097 10013 21131 10047
rect 21131 10013 21140 10047
rect 21088 10004 21140 10013
rect 28080 10208 28132 10260
rect 28908 10251 28960 10260
rect 28908 10217 28917 10251
rect 28917 10217 28951 10251
rect 28951 10217 28960 10251
rect 28908 10208 28960 10217
rect 30380 10208 30432 10260
rect 30932 10208 30984 10260
rect 32864 10208 32916 10260
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25872 10072 25924 10124
rect 29736 10140 29788 10192
rect 25780 10047 25832 10056
rect 25780 10013 25789 10047
rect 25789 10013 25823 10047
rect 25823 10013 25832 10047
rect 25780 10004 25832 10013
rect 26608 10004 26660 10056
rect 22192 9936 22244 9988
rect 23940 9936 23992 9988
rect 28448 10072 28500 10124
rect 28816 10072 28868 10124
rect 27160 10047 27212 10056
rect 27160 10013 27169 10047
rect 27169 10013 27203 10047
rect 27203 10013 27212 10047
rect 27160 10004 27212 10013
rect 27344 10047 27396 10056
rect 27344 10013 27353 10047
rect 27353 10013 27387 10047
rect 27387 10013 27396 10047
rect 27344 10004 27396 10013
rect 16764 9911 16816 9920
rect 16764 9877 16773 9911
rect 16773 9877 16807 9911
rect 16807 9877 16816 9911
rect 16764 9868 16816 9877
rect 23296 9868 23348 9920
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 25320 9868 25372 9920
rect 27896 9936 27948 9988
rect 25964 9868 26016 9920
rect 27528 9911 27580 9920
rect 27528 9877 27537 9911
rect 27537 9877 27571 9911
rect 27571 9877 27580 9911
rect 27528 9868 27580 9877
rect 28264 9868 28316 9920
rect 29184 10004 29236 10056
rect 29644 10072 29696 10124
rect 30840 10115 30892 10124
rect 30840 10081 30849 10115
rect 30849 10081 30883 10115
rect 30883 10081 30892 10115
rect 30840 10072 30892 10081
rect 30380 10049 30432 10056
rect 30380 10015 30389 10049
rect 30389 10015 30423 10049
rect 30423 10015 30432 10049
rect 30380 10004 30432 10015
rect 31300 9936 31352 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 9220 9664 9272 9716
rect 9772 9664 9824 9716
rect 10508 9664 10560 9716
rect 10784 9664 10836 9716
rect 12440 9664 12492 9716
rect 12716 9664 12768 9716
rect 22192 9707 22244 9716
rect 22192 9673 22201 9707
rect 22201 9673 22235 9707
rect 22235 9673 22244 9707
rect 22192 9664 22244 9673
rect 24032 9707 24084 9716
rect 24032 9673 24041 9707
rect 24041 9673 24075 9707
rect 24075 9673 24084 9707
rect 24032 9664 24084 9673
rect 25780 9707 25832 9716
rect 25780 9673 25789 9707
rect 25789 9673 25823 9707
rect 25823 9673 25832 9707
rect 25780 9664 25832 9673
rect 25964 9664 26016 9716
rect 11520 9528 11572 9580
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 14004 9528 14056 9580
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 15936 9460 15988 9512
rect 25412 9639 25464 9648
rect 25412 9605 25421 9639
rect 25421 9605 25455 9639
rect 25455 9605 25464 9639
rect 25412 9596 25464 9605
rect 26056 9596 26108 9648
rect 27988 9707 28040 9716
rect 27988 9673 27997 9707
rect 27997 9673 28031 9707
rect 28031 9673 28040 9707
rect 27988 9664 28040 9673
rect 29000 9664 29052 9716
rect 29092 9664 29144 9716
rect 30380 9664 30432 9716
rect 31300 9664 31352 9716
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 22008 9528 22060 9580
rect 23020 9571 23072 9580
rect 23020 9537 23029 9571
rect 23029 9537 23063 9571
rect 23063 9537 23072 9571
rect 23020 9528 23072 9537
rect 23296 9571 23348 9580
rect 23296 9537 23305 9571
rect 23305 9537 23339 9571
rect 23339 9537 23348 9571
rect 23296 9528 23348 9537
rect 23940 9528 23992 9580
rect 28172 9571 28224 9580
rect 28172 9537 28181 9571
rect 28181 9537 28215 9571
rect 28215 9537 28224 9571
rect 28172 9528 28224 9537
rect 14556 9392 14608 9444
rect 10324 9324 10376 9376
rect 10692 9324 10744 9376
rect 10968 9324 11020 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 15476 9324 15528 9376
rect 18052 9324 18104 9376
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 28264 9460 28316 9512
rect 27344 9392 27396 9444
rect 25320 9324 25372 9376
rect 29644 9324 29696 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 11520 9163 11572 9172
rect 11520 9129 11529 9163
rect 11529 9129 11563 9163
rect 11563 9129 11572 9163
rect 11520 9120 11572 9129
rect 14556 9120 14608 9172
rect 15476 9120 15528 9172
rect 15936 9163 15988 9172
rect 15936 9129 15945 9163
rect 15945 9129 15979 9163
rect 15979 9129 15988 9163
rect 15936 9120 15988 9129
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 17224 9120 17276 9172
rect 10692 8916 10744 8968
rect 12256 8916 12308 8968
rect 10968 8780 11020 8832
rect 14740 8891 14792 8900
rect 14740 8857 14749 8891
rect 14749 8857 14783 8891
rect 14783 8857 14792 8891
rect 14740 8848 14792 8857
rect 18972 9120 19024 9172
rect 19708 9120 19760 9172
rect 20076 9120 20128 9172
rect 17684 8916 17736 8968
rect 17776 8959 17828 8968
rect 17776 8925 17785 8959
rect 17785 8925 17819 8959
rect 17819 8925 17828 8959
rect 17776 8916 17828 8925
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 20260 9095 20312 9104
rect 20260 9061 20269 9095
rect 20269 9061 20303 9095
rect 20303 9061 20312 9095
rect 20260 9052 20312 9061
rect 21088 8984 21140 9036
rect 22100 9027 22152 9036
rect 22100 8993 22109 9027
rect 22109 8993 22143 9027
rect 22143 8993 22152 9027
rect 22100 8984 22152 8993
rect 23020 8984 23072 9036
rect 18144 8891 18196 8900
rect 18144 8857 18153 8891
rect 18153 8857 18187 8891
rect 18187 8857 18196 8891
rect 18144 8848 18196 8857
rect 17500 8780 17552 8832
rect 25228 9095 25280 9104
rect 25228 9061 25237 9095
rect 25237 9061 25271 9095
rect 25271 9061 25280 9095
rect 25228 9052 25280 9061
rect 24492 8984 24544 9036
rect 26056 9052 26108 9104
rect 28172 9120 28224 9172
rect 29644 9120 29696 9172
rect 31300 9163 31352 9172
rect 31300 9129 31309 9163
rect 31309 9129 31343 9163
rect 31343 9129 31352 9163
rect 31300 9120 31352 9129
rect 26608 9052 26660 9104
rect 27436 9052 27488 9104
rect 28632 9052 28684 9104
rect 27344 9027 27396 9036
rect 27344 8993 27353 9027
rect 27353 8993 27387 9027
rect 27387 8993 27396 9027
rect 27344 8984 27396 8993
rect 25136 8916 25188 8968
rect 27528 8916 27580 8968
rect 28264 8959 28316 8968
rect 28264 8925 28273 8959
rect 28273 8925 28307 8959
rect 28307 8925 28316 8959
rect 28264 8916 28316 8925
rect 20996 8780 21048 8832
rect 21272 8780 21324 8832
rect 23204 8823 23256 8832
rect 23204 8789 23213 8823
rect 23213 8789 23247 8823
rect 23247 8789 23256 8823
rect 23204 8780 23256 8789
rect 24676 8780 24728 8832
rect 29000 8916 29052 8968
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 26700 8823 26752 8832
rect 26700 8789 26709 8823
rect 26709 8789 26743 8823
rect 26743 8789 26752 8823
rect 26700 8780 26752 8789
rect 27620 8780 27672 8832
rect 27988 8780 28040 8832
rect 28908 8891 28960 8900
rect 28908 8857 28917 8891
rect 28917 8857 28951 8891
rect 28951 8857 28960 8891
rect 28908 8848 28960 8857
rect 30104 8848 30156 8900
rect 29828 8780 29880 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 15016 8576 15068 8628
rect 15568 8576 15620 8628
rect 16764 8576 16816 8628
rect 17776 8576 17828 8628
rect 12624 8508 12676 8560
rect 14372 8508 14424 8560
rect 18144 8508 18196 8560
rect 23204 8576 23256 8628
rect 26056 8576 26108 8628
rect 26700 8576 26752 8628
rect 27988 8576 28040 8628
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 30104 8619 30156 8628
rect 30104 8585 30113 8619
rect 30113 8585 30147 8619
rect 30147 8585 30156 8619
rect 30104 8576 30156 8585
rect 23572 8508 23624 8560
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 13176 8236 13228 8288
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 16856 8372 16908 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 17684 8372 17736 8424
rect 17960 8372 18012 8424
rect 15476 8304 15528 8356
rect 18144 8304 18196 8356
rect 21088 8440 21140 8492
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 21824 8440 21876 8492
rect 19708 8415 19760 8424
rect 19708 8381 19717 8415
rect 19717 8381 19751 8415
rect 19751 8381 19760 8415
rect 19708 8372 19760 8381
rect 22008 8372 22060 8424
rect 23480 8372 23532 8424
rect 25596 8508 25648 8560
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 25136 8304 25188 8356
rect 25504 8415 25556 8424
rect 25504 8381 25513 8415
rect 25513 8381 25547 8415
rect 25547 8381 25556 8415
rect 25504 8372 25556 8381
rect 27620 8440 27672 8492
rect 28908 8440 28960 8492
rect 27436 8415 27488 8424
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 29184 8440 29236 8492
rect 30472 8508 30524 8560
rect 29736 8440 29788 8492
rect 38200 8483 38252 8492
rect 38200 8449 38209 8483
rect 38209 8449 38243 8483
rect 38243 8449 38252 8483
rect 38200 8440 38252 8449
rect 27988 8304 28040 8356
rect 38384 8347 38436 8356
rect 38384 8313 38393 8347
rect 38393 8313 38427 8347
rect 38427 8313 38436 8347
rect 38384 8304 38436 8313
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 26608 8279 26660 8288
rect 26608 8245 26617 8279
rect 26617 8245 26651 8279
rect 26651 8245 26660 8279
rect 26608 8236 26660 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11888 8032 11940 8084
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 15476 8032 15528 8084
rect 17132 8032 17184 8084
rect 18144 8032 18196 8084
rect 10692 7964 10744 8016
rect 12716 7828 12768 7880
rect 19708 8032 19760 8084
rect 21456 8032 21508 8084
rect 23572 8075 23624 8084
rect 23572 8041 23581 8075
rect 23581 8041 23615 8075
rect 23615 8041 23624 8075
rect 23572 8032 23624 8041
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13452 7760 13504 7812
rect 15844 7803 15896 7812
rect 15844 7769 15853 7803
rect 15853 7769 15887 7803
rect 15887 7769 15896 7803
rect 15844 7760 15896 7769
rect 18328 7760 18380 7812
rect 20260 7828 20312 7880
rect 14188 7692 14240 7744
rect 18052 7692 18104 7744
rect 21088 7760 21140 7812
rect 22100 7896 22152 7948
rect 29000 8032 29052 8084
rect 26608 7896 26660 7948
rect 27988 7896 28040 7948
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 27252 7760 27304 7812
rect 21272 7692 21324 7744
rect 28908 7828 28960 7880
rect 29000 7692 29052 7744
rect 29184 7692 29236 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 15844 7488 15896 7540
rect 16672 7488 16724 7540
rect 17132 7488 17184 7540
rect 23480 7488 23532 7540
rect 27252 7488 27304 7540
rect 18328 7352 18380 7404
rect 29736 7352 29788 7404
rect 18052 7148 18104 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 15474 39200 15530 40000
rect 17406 39200 17462 40000
rect 19338 39200 19394 40000
rect 21914 39200 21970 40000
rect 23202 39200 23258 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 15488 37466 15516 39200
rect 17420 37466 17448 39200
rect 19352 37466 19380 39200
rect 21928 37466 21956 39200
rect 15476 37460 15528 37466
rect 15476 37402 15528 37408
rect 17408 37460 17460 37466
rect 17408 37402 17460 37408
rect 19340 37460 19392 37466
rect 19340 37402 19392 37408
rect 21916 37460 21968 37466
rect 21916 37402 21968 37408
rect 15660 37188 15712 37194
rect 15660 37130 15712 37136
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 19524 37188 19576 37194
rect 19524 37130 19576 37136
rect 22376 37188 22428 37194
rect 22376 37130 22428 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 15672 35894 15700 37130
rect 17328 35894 17356 37130
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 15580 35866 15700 35894
rect 17236 35866 17356 35894
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 15580 31754 15608 35866
rect 15488 31726 15608 31754
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 7564 31272 7616 31278
rect 7564 31214 7616 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 7576 30938 7604 31214
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 8220 30938 8248 31078
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 6380 30258 6408 30534
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 3422 30016 3478 30025
rect 3422 29951 3478 29960
rect 3332 26920 3384 26926
rect 3332 26862 3384 26868
rect 3344 26586 3372 26862
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 1676 25696 1728 25702
rect 1676 25638 1728 25644
rect 938 25256 994 25265
rect 938 25191 994 25200
rect 952 25158 980 25191
rect 940 25152 992 25158
rect 940 25094 992 25100
rect 1688 24818 1716 25638
rect 2792 25498 2820 25842
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 2780 25492 2832 25498
rect 2780 25434 2832 25440
rect 3160 25430 3188 25638
rect 3344 25498 3372 26522
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3148 25424 3200 25430
rect 3148 25366 3200 25372
rect 3240 25356 3292 25362
rect 3240 25298 3292 25304
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 1964 24954 1992 25230
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 2136 24880 2188 24886
rect 2136 24822 2188 24828
rect 1676 24812 1728 24818
rect 1676 24754 1728 24760
rect 1124 24608 1176 24614
rect 1122 24576 1124 24585
rect 1176 24576 1178 24585
rect 1122 24511 1178 24520
rect 2044 24132 2096 24138
rect 2044 24074 2096 24080
rect 2056 23866 2084 24074
rect 2148 23866 2176 24822
rect 2884 24818 2912 25162
rect 3252 24886 3280 25298
rect 3240 24880 3292 24886
rect 3240 24822 3292 24828
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 3252 24410 3280 24822
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3252 24206 3280 24346
rect 3344 24206 3372 24754
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3252 23866 3280 24006
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 2136 23860 2188 23866
rect 2136 23802 2188 23808
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 2884 22778 2912 23054
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21554 3280 21830
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3436 19446 3464 29951
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 6276 29640 6328 29646
rect 6276 29582 6328 29588
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5368 28558 5396 29446
rect 5828 29306 5856 29582
rect 6092 29572 6144 29578
rect 6092 29514 6144 29520
rect 6000 29504 6052 29510
rect 6000 29446 6052 29452
rect 6012 29306 6040 29446
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 6000 29300 6052 29306
rect 6000 29242 6052 29248
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 5552 28626 5580 28902
rect 6104 28626 6132 29514
rect 6288 29170 6316 29582
rect 7116 29510 7144 30534
rect 7208 29578 7236 30670
rect 7484 30394 7512 30670
rect 7472 30388 7524 30394
rect 7472 30330 7524 30336
rect 7380 30048 7432 30054
rect 7380 29990 7432 29996
rect 7392 29646 7420 29990
rect 7852 29782 7880 30738
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 12256 30728 12308 30734
rect 12256 30670 12308 30676
rect 8392 30592 8444 30598
rect 8392 30534 8444 30540
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8404 30326 8432 30534
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 7840 29776 7892 29782
rect 7840 29718 7892 29724
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 7196 29572 7248 29578
rect 7196 29514 7248 29520
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 6368 29232 6420 29238
rect 6368 29174 6420 29180
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 6380 28626 6408 29174
rect 8312 29170 8340 29582
rect 8496 29578 8524 30534
rect 10612 30394 10640 30670
rect 10784 30592 10836 30598
rect 10784 30534 10836 30540
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 10600 30388 10652 30394
rect 10600 30330 10652 30336
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 8484 29572 8536 29578
rect 8484 29514 8536 29520
rect 9588 29572 9640 29578
rect 9588 29514 9640 29520
rect 8668 29504 8720 29510
rect 8668 29446 8720 29452
rect 6644 29164 6696 29170
rect 6644 29106 6696 29112
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 6460 29028 6512 29034
rect 6460 28970 6512 28976
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 6092 28620 6144 28626
rect 6092 28562 6144 28568
rect 6368 28620 6420 28626
rect 6368 28562 6420 28568
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5552 27878 5580 28562
rect 5816 28484 5868 28490
rect 5816 28426 5868 28432
rect 5828 28218 5856 28426
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5552 27674 5580 27814
rect 4068 27668 4120 27674
rect 4068 27610 4120 27616
rect 5540 27668 5592 27674
rect 5540 27610 5592 27616
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3804 26450 3832 27406
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3608 26308 3660 26314
rect 3608 26250 3660 26256
rect 3516 25900 3568 25906
rect 3516 25842 3568 25848
rect 3528 25498 3556 25842
rect 3620 25498 3648 26250
rect 3804 25906 3832 26386
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3792 25900 3844 25906
rect 3792 25842 3844 25848
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3516 25492 3568 25498
rect 3516 25434 3568 25440
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3712 24954 3740 25638
rect 3700 24948 3752 24954
rect 3700 24890 3752 24896
rect 3804 24818 3832 25842
rect 3896 25294 3924 26182
rect 4080 25838 4108 27610
rect 4160 27396 4212 27402
rect 4160 27338 4212 27344
rect 4172 27130 4200 27338
rect 5264 27328 5316 27334
rect 5264 27270 5316 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5276 27130 5304 27270
rect 5552 27130 5580 27610
rect 6092 27328 6144 27334
rect 6092 27270 6144 27276
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 6104 26994 6132 27270
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5632 26852 5684 26858
rect 5632 26794 5684 26800
rect 4620 26784 4672 26790
rect 4620 26726 4672 26732
rect 5540 26784 5592 26790
rect 5540 26726 5592 26732
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 4448 26042 4476 26318
rect 4632 26042 4660 26726
rect 4804 26240 4856 26246
rect 4804 26182 4856 26188
rect 4816 26042 4844 26182
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5552 26042 5580 26726
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4620 26036 4672 26042
rect 4620 25978 4672 25984
rect 4804 26036 4856 26042
rect 4804 25978 4856 25984
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5644 25906 5672 26794
rect 6104 26586 6132 26930
rect 6092 26580 6144 26586
rect 6092 26522 6144 26528
rect 6380 26450 6408 28562
rect 6472 28218 6500 28970
rect 6564 28762 6592 29038
rect 6656 28966 6684 29106
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 7288 28960 7340 28966
rect 7288 28902 7340 28908
rect 7472 28960 7524 28966
rect 7472 28902 7524 28908
rect 6552 28756 6604 28762
rect 6552 28698 6604 28704
rect 6644 28484 6696 28490
rect 6644 28426 6696 28432
rect 6656 28218 6684 28426
rect 7300 28218 7328 28902
rect 6460 28212 6512 28218
rect 6460 28154 6512 28160
rect 6644 28212 6696 28218
rect 6644 28154 6696 28160
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 6472 27674 6500 28154
rect 6920 28144 6972 28150
rect 6920 28086 6972 28092
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 6368 26444 6420 26450
rect 6368 26386 6420 26392
rect 5632 25900 5684 25906
rect 5632 25842 5684 25848
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 4080 25362 4108 25774
rect 6932 25770 6960 28086
rect 7484 27878 7512 28902
rect 8036 28762 8064 29038
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7380 27328 7432 27334
rect 7380 27270 7432 27276
rect 7392 27130 7420 27270
rect 7380 27124 7432 27130
rect 7380 27066 7432 27072
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7208 26382 7236 26726
rect 7196 26376 7248 26382
rect 7196 26318 7248 26324
rect 7852 25906 7880 26862
rect 8220 26586 8248 26930
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 5276 25294 5304 25638
rect 3884 25288 3936 25294
rect 3884 25230 3936 25236
rect 5264 25288 5316 25294
rect 5264 25230 5316 25236
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4816 24886 4844 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3712 24206 3740 24550
rect 3804 24274 3832 24754
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3792 24268 3844 24274
rect 3792 24210 3844 24216
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 3620 22642 3648 22918
rect 3804 22778 3832 24210
rect 3896 23866 3924 24686
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 5460 24410 5488 25230
rect 5552 24954 5580 25230
rect 7852 25226 7880 25842
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 7840 25220 7892 25226
rect 7840 25162 7892 25168
rect 5540 24948 5592 24954
rect 5540 24890 5592 24896
rect 6184 24812 6236 24818
rect 6184 24754 6236 24760
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5552 24614 5580 24686
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4160 24064 4212 24070
rect 4080 24012 4160 24018
rect 4080 24006 4212 24012
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 4080 23990 4200 24006
rect 4080 23866 4108 23990
rect 3884 23860 3936 23866
rect 3884 23802 3936 23808
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4724 23662 4752 24006
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4816 23594 4844 24278
rect 5552 24206 5580 24550
rect 6196 24410 6224 24754
rect 6828 24676 6880 24682
rect 6828 24618 6880 24624
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 5356 24200 5408 24206
rect 5356 24142 5408 24148
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5368 23866 5396 24142
rect 6840 24070 6868 24618
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7392 24410 7420 24550
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 5460 23866 5488 24006
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 6840 23798 6868 24006
rect 7668 23866 7696 24074
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 6828 23792 6880 23798
rect 6828 23734 6880 23740
rect 7852 23730 7880 25162
rect 8036 23730 8064 25298
rect 8220 24818 8248 25706
rect 8312 24818 8340 29106
rect 8680 28558 8708 29446
rect 8944 29164 8996 29170
rect 8944 29106 8996 29112
rect 8956 28762 8984 29106
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 9600 28626 9628 29514
rect 9692 29306 9720 29582
rect 10796 29578 10824 30534
rect 11256 30326 11284 30534
rect 11808 30326 11836 30670
rect 12268 30394 12296 30670
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12256 30388 12308 30394
rect 12256 30330 12308 30336
rect 11244 30320 11296 30326
rect 11244 30262 11296 30268
rect 11796 30320 11848 30326
rect 11796 30262 11848 30268
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 12716 30252 12768 30258
rect 12716 30194 12768 30200
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 10784 29572 10836 29578
rect 10784 29514 10836 29520
rect 11072 29510 11100 30126
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9692 28558 9720 29242
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9588 28416 9640 28422
rect 9588 28358 9640 28364
rect 9600 28150 9628 28358
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 9220 28076 9272 28082
rect 9220 28018 9272 28024
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8496 27538 8524 27814
rect 8484 27532 8536 27538
rect 8484 27474 8536 27480
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8404 26314 8432 27406
rect 8496 26382 8524 27474
rect 9232 26586 9260 28018
rect 9416 27674 9444 28018
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9404 27668 9456 27674
rect 9404 27610 9456 27616
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9508 26586 9536 26726
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 9496 26580 9548 26586
rect 9496 26522 9548 26528
rect 9692 26450 9720 27950
rect 9784 27470 9812 27950
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9772 26852 9824 26858
rect 9772 26794 9824 26800
rect 9784 26586 9812 26794
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9680 26444 9732 26450
rect 9680 26386 9732 26392
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 9692 26042 9720 26386
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9876 26042 9904 26318
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8680 25498 8708 25774
rect 10060 25702 10088 29106
rect 11072 29102 11100 29446
rect 11164 29306 11192 30194
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 11152 29300 11204 29306
rect 11152 29242 11204 29248
rect 12360 29102 12388 29990
rect 12452 29850 12480 30126
rect 12728 29850 12756 30194
rect 12440 29844 12492 29850
rect 12440 29786 12492 29792
rect 12716 29844 12768 29850
rect 12716 29786 12768 29792
rect 12912 29714 12940 30534
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13740 29714 13768 30194
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 14108 29714 14136 29990
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 11060 29096 11112 29102
rect 11060 29038 11112 29044
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 10692 28484 10744 28490
rect 10692 28426 10744 28432
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10152 26994 10180 27814
rect 10244 27130 10272 28018
rect 10416 27872 10468 27878
rect 10416 27814 10468 27820
rect 10428 27470 10456 27814
rect 10416 27464 10468 27470
rect 10416 27406 10468 27412
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10140 26988 10192 26994
rect 10140 26930 10192 26936
rect 10336 26926 10364 27270
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10508 26852 10560 26858
rect 10428 26812 10508 26840
rect 10428 26450 10456 26812
rect 10508 26794 10560 26800
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10704 26042 10732 28426
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10796 26994 10824 28154
rect 11072 27470 11100 29038
rect 12360 28626 12388 29038
rect 12636 28762 12664 29038
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 13280 28694 13308 29582
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 13360 29504 13412 29510
rect 13360 29446 13412 29452
rect 13372 29238 13400 29446
rect 14752 29306 14780 29514
rect 14740 29300 14792 29306
rect 14740 29242 14792 29248
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 15108 29232 15160 29238
rect 15108 29174 15160 29180
rect 14556 29096 14608 29102
rect 14556 29038 14608 29044
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 13268 28688 13320 28694
rect 13268 28630 13320 28636
rect 12348 28620 12400 28626
rect 12348 28562 12400 28568
rect 14200 28558 14228 28970
rect 14280 28960 14332 28966
rect 14280 28902 14332 28908
rect 14292 28558 14320 28902
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14280 28552 14332 28558
rect 14280 28494 14332 28500
rect 12072 28484 12124 28490
rect 12072 28426 12124 28432
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 12084 28218 12112 28426
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 11072 27062 11100 27406
rect 11060 27056 11112 27062
rect 11060 26998 11112 27004
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10980 26382 11008 26862
rect 11072 26586 11100 26998
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 9416 25226 9444 25638
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 9404 25220 9456 25226
rect 9404 25162 9456 25168
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 8312 24274 8340 24754
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 8036 23322 8064 23666
rect 8588 23662 8616 24006
rect 9692 23730 9720 24006
rect 9220 23724 9272 23730
rect 9496 23724 9548 23730
rect 9272 23684 9496 23712
rect 9220 23666 9272 23672
rect 9496 23666 9548 23672
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 9048 23474 9076 23598
rect 9496 23588 9548 23594
rect 9496 23530 9548 23536
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9508 23474 9536 23530
rect 9048 23446 9536 23474
rect 9600 23322 9628 23530
rect 9692 23322 9720 23666
rect 9876 23594 9904 25434
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 9968 24274 9996 25230
rect 10796 24954 10824 25230
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 24410 10088 24686
rect 10704 24614 10732 24754
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 10704 23798 10732 24550
rect 10692 23792 10744 23798
rect 10692 23734 10744 23740
rect 10888 23730 10916 24754
rect 10980 24698 11008 25434
rect 11164 24886 11192 26250
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11256 25294 11284 25978
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11336 25152 11388 25158
rect 11336 25094 11388 25100
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11348 24954 11376 25094
rect 11440 24954 11468 25094
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11152 24880 11204 24886
rect 11152 24822 11204 24828
rect 10980 24670 11100 24698
rect 11072 24614 11100 24670
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 10980 24070 11008 24550
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 4528 23112 4580 23118
rect 4528 23054 4580 23060
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 4540 22778 4568 23054
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 6380 22778 6408 23054
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 3804 22234 3832 22714
rect 3974 22536 4030 22545
rect 3974 22471 4030 22480
rect 4540 22522 4568 22714
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 4540 22494 4752 22522
rect 3988 22234 4016 22471
rect 4540 22438 4568 22494
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 4528 22432 4580 22438
rect 4528 22374 4580 22380
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21350 4016 21830
rect 4080 21554 4108 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4724 21486 4752 22494
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4816 21690 4844 21898
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21690 5304 22578
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5460 22386 5488 22510
rect 5540 22500 5592 22506
rect 5540 22442 5592 22448
rect 5368 22358 5488 22386
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 5264 21684 5316 21690
rect 5264 21626 5316 21632
rect 4712 21480 4764 21486
rect 4712 21422 4764 21428
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4724 21146 4752 21422
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 5092 20942 5120 21286
rect 5276 21010 5304 21626
rect 5368 21146 5396 22358
rect 5552 22250 5580 22442
rect 5460 22222 5580 22250
rect 5828 22234 5856 22578
rect 6092 22432 6144 22438
rect 6092 22374 6144 22380
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 5816 22228 5868 22234
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5460 20942 5488 22222
rect 5816 22170 5868 22176
rect 5724 21888 5776 21894
rect 5724 21830 5776 21836
rect 5736 21690 5764 21830
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5828 21622 5856 22170
rect 5816 21616 5868 21622
rect 5816 21558 5868 21564
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5552 21146 5580 21422
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6104 20942 6132 22374
rect 6932 22030 6960 22374
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 7208 21554 7236 22918
rect 9048 22658 9076 23054
rect 9692 22778 9720 23258
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9876 22778 9904 22918
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8864 22630 9076 22658
rect 11072 22642 11100 24142
rect 11060 22636 11112 22642
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 7300 21690 7328 22510
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7576 21962 7604 22374
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7288 21684 7340 21690
rect 7288 21626 7340 21632
rect 8128 21554 8156 22510
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8128 21350 8156 21490
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 21010 8156 21286
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 5448 20936 5500 20942
rect 5448 20878 5500 20884
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4080 20505 4108 20538
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 8312 19854 8340 21966
rect 8404 21690 8432 22510
rect 8496 22386 8524 22578
rect 8760 22568 8812 22574
rect 8760 22510 8812 22516
rect 8668 22432 8720 22438
rect 8496 22358 8616 22386
rect 8668 22374 8720 22380
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8496 21962 8524 22102
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8496 21570 8524 21898
rect 8404 21554 8524 21570
rect 8392 21548 8524 21554
rect 8444 21542 8524 21548
rect 8392 21490 8444 21496
rect 8588 21418 8616 22358
rect 8680 21486 8708 22374
rect 8772 22166 8800 22510
rect 8760 22160 8812 22166
rect 8760 22102 8812 22108
rect 8864 21690 8892 22630
rect 11060 22578 11112 22584
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9048 21894 9076 22374
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 8956 21690 8984 21830
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 9048 21622 9076 21830
rect 10060 21622 10088 22374
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 9048 21146 9076 21558
rect 10152 21146 10180 22510
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10796 22030 10824 22374
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19922 9352 20198
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8300 19848 8352 19854
rect 4066 19816 4122 19825
rect 8300 19790 8352 19796
rect 4066 19751 4122 19760
rect 4080 19514 4108 19751
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4066 18456 4122 18465
rect 4874 18459 5182 18468
rect 4066 18391 4122 18400
rect 4080 18222 4108 18391
rect 8312 18222 8340 19790
rect 9784 18442 9812 20402
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9876 19786 9904 20198
rect 10980 19854 11008 21966
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20466 11100 20742
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 9968 19514 9996 19654
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10704 19378 10732 19654
rect 10980 19378 11008 19790
rect 11164 19378 11192 24822
rect 11532 24818 11560 25638
rect 11624 25430 11652 25842
rect 11900 25702 11928 26930
rect 11992 26382 12020 27406
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12452 26858 12480 27270
rect 12636 27130 12664 27406
rect 13096 27130 13124 28018
rect 13188 27674 13216 28426
rect 13728 28212 13780 28218
rect 13832 28200 13860 28494
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14016 28218 14044 28358
rect 13780 28172 13860 28200
rect 14004 28212 14056 28218
rect 13728 28154 13780 28160
rect 14004 28154 14056 28160
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13280 27538 13308 27950
rect 13268 27532 13320 27538
rect 13268 27474 13320 27480
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 13280 26994 13308 27474
rect 13372 27334 13400 28018
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13544 27396 13596 27402
rect 13544 27338 13596 27344
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12544 26790 12572 26930
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 12544 25906 12572 26726
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11612 25424 11664 25430
rect 11612 25366 11664 25372
rect 12268 25294 12296 25774
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12452 25226 12480 25842
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12636 25498 12664 25638
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11256 24138 11284 24550
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11624 23866 11652 24074
rect 11716 23866 11744 24754
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12360 23866 12388 24074
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12544 23186 12572 23666
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11808 22574 11836 22918
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 12440 22704 12492 22710
rect 12440 22646 12492 22652
rect 11900 22574 11928 22646
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11888 22568 11940 22574
rect 11888 22510 11940 22516
rect 12452 22234 12480 22646
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12544 22030 12572 23122
rect 12636 22982 12664 25434
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12728 25158 12756 25298
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 13188 24070 13216 26862
rect 13372 25838 13400 27270
rect 13556 27130 13584 27338
rect 13544 27124 13596 27130
rect 13544 27066 13596 27072
rect 13648 26042 13676 27474
rect 14384 27470 14412 27814
rect 14568 27470 14596 29038
rect 14740 27940 14792 27946
rect 14740 27882 14792 27888
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14660 27538 14688 27814
rect 14752 27674 14780 27882
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13726 27160 13782 27169
rect 13832 27130 13860 27270
rect 14292 27130 14320 27406
rect 14384 27282 14412 27406
rect 14384 27254 14504 27282
rect 13726 27095 13728 27104
rect 13780 27095 13782 27104
rect 13820 27124 13872 27130
rect 13728 27066 13780 27072
rect 13820 27066 13872 27072
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14476 26994 14504 27254
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14752 26926 14780 27610
rect 15120 27606 15148 29174
rect 15212 29170 15240 29242
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15212 28218 15240 29106
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 15396 27470 15424 27814
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 13912 26920 13964 26926
rect 13912 26862 13964 26868
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 13728 26376 13780 26382
rect 13728 26318 13780 26324
rect 13740 26042 13768 26318
rect 13924 26042 13952 26862
rect 15028 26382 15056 27406
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15212 26586 15240 26930
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15016 26376 15068 26382
rect 15016 26318 15068 26324
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13372 24818 13400 25774
rect 13464 25498 13492 25842
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13648 24886 13676 25978
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15028 25498 15056 25638
rect 15016 25492 15068 25498
rect 15016 25434 15068 25440
rect 15304 25294 15332 27406
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15396 25498 15424 26930
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 14476 24954 14504 25230
rect 14832 25220 14884 25226
rect 14832 25162 14884 25168
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 13820 24948 13872 24954
rect 13820 24890 13872 24896
rect 14464 24948 14516 24954
rect 14464 24890 14516 24896
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13832 24818 13860 24890
rect 14844 24834 14872 25162
rect 15396 24954 15424 25162
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15396 24834 15424 24890
rect 14752 24818 14872 24834
rect 15304 24818 15424 24834
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14740 24812 14872 24818
rect 14792 24806 14872 24812
rect 15108 24812 15160 24818
rect 14740 24754 14792 24760
rect 15108 24754 15160 24760
rect 15292 24812 15424 24818
rect 15344 24806 15424 24812
rect 15292 24754 15344 24760
rect 13556 24614 13584 24754
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13924 24342 13952 24754
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 12912 23866 12940 24006
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 11532 21690 11560 21966
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 12072 21616 12124 21622
rect 12072 21558 12124 21564
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11808 21146 11836 21422
rect 12084 21146 12112 21558
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20330 11652 20878
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20324 11664 20330
rect 11612 20266 11664 20272
rect 11716 19718 11744 20402
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 12530 20360 12586 20369
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11900 19854 11928 20198
rect 11992 19990 12020 20334
rect 12530 20295 12532 20304
rect 12584 20295 12586 20304
rect 12532 20266 12584 20272
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 12544 19922 12572 20266
rect 12636 19990 12664 22918
rect 12808 21344 12860 21350
rect 12728 21304 12808 21332
rect 12728 20398 12756 21304
rect 12808 21286 12860 21292
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 20262 12756 20334
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12728 19854 12756 20198
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11152 19372 11204 19378
rect 11204 19320 11376 19334
rect 11152 19314 11376 19320
rect 10980 18986 11008 19314
rect 11164 19306 11376 19314
rect 10888 18970 11008 18986
rect 10876 18964 11008 18970
rect 10928 18958 11008 18964
rect 10876 18906 10928 18912
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9692 18414 9812 18442
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 8312 16998 8340 18158
rect 8772 17882 8800 18158
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 9692 17678 9720 18414
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9784 17882 9812 18294
rect 9876 18086 9904 18566
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 9876 17882 9904 18022
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 10244 17678 10272 18022
rect 10888 17746 10916 18906
rect 10876 17740 10928 17746
rect 10876 17682 10928 17688
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 8312 16182 8340 16934
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 2778 15736 2834 15745
rect 4214 15739 4522 15748
rect 2778 15671 2834 15680
rect 2792 15434 2820 15671
rect 2780 15428 2832 15434
rect 2780 15370 2832 15376
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 7760 14074 7788 15982
rect 8036 15706 8064 15982
rect 9140 15978 9168 17478
rect 9232 16794 9260 17614
rect 10244 16794 10272 17614
rect 11348 17270 11376 19306
rect 12728 18834 12756 19790
rect 12992 19440 13044 19446
rect 12990 19408 12992 19417
rect 13044 19408 13046 19417
rect 12990 19343 13046 19352
rect 13096 18834 13124 20470
rect 13188 18970 13216 24006
rect 13280 23866 13308 24006
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13556 23186 13584 24210
rect 13924 23866 13952 24278
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13636 22772 13688 22778
rect 13832 22760 13860 23122
rect 13924 22778 13952 23462
rect 14568 23186 14596 24754
rect 14752 23594 14780 24754
rect 15120 24426 15148 24754
rect 15488 24614 15516 31726
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15580 30190 15608 30670
rect 15568 30184 15620 30190
rect 15568 30126 15620 30132
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15764 29646 15792 29990
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 16488 29572 16540 29578
rect 16488 29514 16540 29520
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16500 29238 16528 29514
rect 16868 29306 16896 29514
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 15752 28076 15804 28082
rect 15752 28018 15804 28024
rect 15660 27464 15712 27470
rect 15660 27406 15712 27412
rect 15672 27130 15700 27406
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15764 26994 15792 28018
rect 16316 27878 16344 28494
rect 16408 28150 16436 28562
rect 16500 28150 16528 29174
rect 17052 29170 17080 29446
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 16764 28620 16816 28626
rect 16764 28562 16816 28568
rect 16396 28144 16448 28150
rect 16396 28086 16448 28092
rect 16488 28144 16540 28150
rect 16488 28086 16540 28092
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16316 27062 16344 27814
rect 16776 27470 16804 28562
rect 17052 28558 17080 29106
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 17144 27606 17172 29106
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 16948 27532 17000 27538
rect 16948 27474 17000 27480
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16304 27056 16356 27062
rect 16304 26998 16356 27004
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15580 26246 15608 26930
rect 15672 26382 15700 26930
rect 15764 26382 15792 26930
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15764 25294 15792 26318
rect 16316 25294 16344 26998
rect 16592 26586 16620 27406
rect 16960 27169 16988 27474
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 17038 27296 17094 27305
rect 17038 27231 17094 27240
rect 16946 27160 17002 27169
rect 17052 27130 17080 27231
rect 16946 27095 17002 27104
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 17038 27024 17094 27033
rect 16960 26994 17038 27010
rect 16948 26988 17038 26994
rect 17000 26982 17038 26988
rect 17038 26959 17094 26968
rect 16948 26930 17000 26936
rect 16946 26888 17002 26897
rect 16946 26823 16948 26832
rect 17000 26823 17002 26832
rect 16948 26794 17000 26800
rect 16580 26580 16632 26586
rect 16580 26522 16632 26528
rect 16856 26444 16908 26450
rect 16856 26386 16908 26392
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16592 25702 16620 26250
rect 16868 26042 16896 26386
rect 16960 26382 16988 26794
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16776 25498 16804 25842
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 15764 24954 15792 25230
rect 15752 24948 15804 24954
rect 15752 24890 15804 24896
rect 17052 24886 17080 25298
rect 17144 25158 17172 27338
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 15120 24398 15240 24426
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14844 23662 14872 24006
rect 15212 23730 15240 24398
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 15016 23588 15068 23594
rect 15016 23530 15068 23536
rect 14556 23180 14608 23186
rect 14556 23122 14608 23128
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 13688 22732 13860 22760
rect 13912 22772 13964 22778
rect 13636 22714 13688 22720
rect 13912 22714 13964 22720
rect 14476 22710 14504 22918
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13556 22094 13584 22374
rect 13556 22066 13676 22094
rect 13268 21956 13320 21962
rect 13268 21898 13320 21904
rect 13280 21350 13308 21898
rect 13648 21690 13676 22066
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14016 21894 14044 22034
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13280 18970 13308 20334
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13372 18834 13400 19858
rect 13556 19378 13584 20402
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10980 16658 11008 17070
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 9956 16584 10008 16590
rect 9402 16552 9458 16561
rect 9956 16526 10008 16532
rect 9402 16487 9404 16496
rect 9456 16487 9458 16496
rect 9404 16458 9456 16464
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 8312 14006 8340 14214
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 4066 13696 4122 13705
rect 4066 13631 4122 13640
rect 4080 13530 4108 13631
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8680 13530 8708 13942
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 8864 12238 8892 12582
rect 8956 12238 8984 14010
rect 9140 13258 9168 15914
rect 9968 15910 9996 16526
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9876 15502 9904 15846
rect 9968 15502 9996 15846
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 15314 9996 15438
rect 10060 15366 10088 16050
rect 9876 15286 9996 15314
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 14074 9720 14214
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9692 13326 9720 14010
rect 9876 13938 9904 15286
rect 10336 14482 10364 16594
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 15706 10456 16390
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10704 15570 10732 16526
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16250 10824 16390
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 11164 16182 11192 16594
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11164 15638 11192 16118
rect 11532 16114 11560 18362
rect 11624 17746 11652 18702
rect 12176 18426 12204 18770
rect 13556 18766 13584 19314
rect 13648 19174 13676 21626
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13740 19854 13768 20198
rect 14016 20058 14044 20334
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 13912 19984 13964 19990
rect 14108 19938 14136 20878
rect 13964 19932 14136 19938
rect 13912 19926 14136 19932
rect 13924 19910 14136 19926
rect 14200 19922 14228 21490
rect 14464 21344 14516 21350
rect 14384 21304 14464 21332
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13740 19378 13768 19654
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 14108 19310 14136 19910
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19514 14320 19790
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 13004 18290 13032 18634
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11624 17338 11652 17682
rect 12544 17678 12572 18158
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17338 12756 17478
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 11624 16114 11652 17274
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11992 16590 12020 16934
rect 12728 16794 12756 17274
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12072 16176 12124 16182
rect 12072 16118 12124 16124
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 11532 15502 11560 16050
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15570 12020 15846
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11164 15094 11192 15302
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9876 13326 9904 13874
rect 9968 13530 9996 13874
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4066 11656 4122 11665
rect 4066 11591 4068 11600
rect 4120 11591 4122 11600
rect 4068 11562 4120 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 8956 10130 8984 12174
rect 9140 11694 9168 13194
rect 10060 12782 10088 14418
rect 11164 14414 11192 15030
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11532 14482 11560 14962
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11532 14074 11560 14418
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11900 13462 11928 13874
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11898 9720 12106
rect 9876 12102 9904 12718
rect 10060 12434 10088 12718
rect 10060 12406 10272 12434
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9876 11762 9904 12038
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11082 9168 11630
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 10244 10606 10272 12406
rect 10336 11694 10364 13262
rect 11900 12782 11928 13398
rect 11992 12986 12020 15370
rect 12084 15366 12112 16118
rect 12176 15910 12204 16458
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 13870 12112 15302
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11992 12782 12020 12922
rect 12176 12782 12204 15438
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14074 12664 14350
rect 12912 14346 12940 17818
rect 13004 17678 13032 18226
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13372 16114 13400 16458
rect 13556 16114 13584 16526
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 12900 14340 12952 14346
rect 12820 14300 12900 14328
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11808 12306 11836 12718
rect 12268 12442 12296 13194
rect 12348 12980 12400 12986
rect 12532 12980 12584 12986
rect 12348 12922 12400 12928
rect 12452 12940 12532 12968
rect 12360 12832 12388 12922
rect 12452 12832 12480 12940
rect 12532 12922 12584 12928
rect 12820 12850 12848 14300
rect 12900 14282 12952 14288
rect 13004 14278 13032 14758
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13462 13032 14214
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 13004 13326 13032 13398
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 12986 12940 13194
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12360 12804 12480 12832
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12256 12436 12308 12442
rect 12452 12434 12480 12582
rect 12452 12406 12572 12434
rect 12256 12378 12308 12384
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 9232 9722 9260 9930
rect 9784 9722 9812 10406
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 10336 9382 10364 11630
rect 10704 11150 10732 12038
rect 11808 11898 11836 12242
rect 12268 12102 12296 12378
rect 12544 12238 12572 12406
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12256 12096 12308 12102
rect 12256 12038 12308 12044
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11808 11234 11836 11834
rect 11808 11206 12020 11234
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10266 10548 10610
rect 10796 10606 10824 11018
rect 11716 10810 11744 11086
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11808 10674 11836 11206
rect 11992 11150 12020 11206
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10520 9722 10548 10202
rect 10612 10062 10640 10406
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10796 9722 10824 10542
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 11532 9586 11560 10066
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 10704 8974 10732 9318
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 10704 8022 10732 8910
rect 10980 8838 11008 9318
rect 11532 9178 11560 9522
rect 12268 9518 12296 12038
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12360 10606 12388 11222
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12452 10742 12480 11086
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12452 10266 12480 10678
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12544 10266 12572 10474
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10266 12664 10406
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12820 10062 12848 12786
rect 13188 10062 13216 14350
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13326 13308 13670
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 12986 13400 13398
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13464 12374 13492 13194
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13648 12238 13676 19110
rect 14384 18426 14412 21304
rect 14464 21286 14516 21292
rect 14660 20942 14688 21898
rect 15028 21622 15056 23530
rect 15212 22778 15240 23666
rect 16776 23594 16804 24754
rect 17144 23866 17172 25094
rect 17236 24614 17264 35866
rect 19536 31754 19564 37130
rect 19536 31726 19656 31754
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17604 30258 17632 30534
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17604 29850 17632 30194
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17592 29572 17644 29578
rect 17592 29514 17644 29520
rect 17604 29306 17632 29514
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17512 29102 17540 29242
rect 18052 29232 18104 29238
rect 18052 29174 18104 29180
rect 17500 29096 17552 29102
rect 17500 29038 17552 29044
rect 17960 28960 18012 28966
rect 17960 28902 18012 28908
rect 17972 28558 18000 28902
rect 18064 28626 18092 29174
rect 18156 29102 18184 29990
rect 19524 29232 19576 29238
rect 19524 29174 19576 29180
rect 18144 29096 18196 29102
rect 18512 29096 18564 29102
rect 18196 29044 18368 29050
rect 18144 29038 18368 29044
rect 18512 29038 18564 29044
rect 18156 29022 18368 29038
rect 18236 28960 18288 28966
rect 18236 28902 18288 28908
rect 18248 28762 18276 28902
rect 18340 28762 18368 29022
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18524 28694 18552 29038
rect 19536 28762 19564 29174
rect 19524 28756 19576 28762
rect 19524 28698 19576 28704
rect 18512 28688 18564 28694
rect 18512 28630 18564 28636
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17316 27056 17368 27062
rect 17316 26998 17368 27004
rect 17328 26790 17356 26998
rect 17420 26994 17448 28494
rect 18524 28490 18552 28630
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18604 28484 18656 28490
rect 18604 28426 18656 28432
rect 18524 28150 18552 28426
rect 18616 28218 18644 28426
rect 19156 28416 19208 28422
rect 19156 28358 19208 28364
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19168 28218 19196 28358
rect 19260 28218 19288 28358
rect 18604 28212 18656 28218
rect 18604 28154 18656 28160
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 18512 28144 18564 28150
rect 18512 28086 18564 28092
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18696 28076 18748 28082
rect 18696 28018 18748 28024
rect 19156 28076 19208 28082
rect 19156 28018 19208 28024
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18052 27396 18104 27402
rect 18052 27338 18104 27344
rect 17682 27296 17738 27305
rect 17682 27231 17738 27240
rect 17696 26994 17724 27231
rect 18064 26994 18092 27338
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17512 26382 17540 26794
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17788 26246 17816 26930
rect 18064 26586 18092 26930
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 17776 26240 17828 26246
rect 17776 26182 17828 26188
rect 18248 25906 18276 27406
rect 18328 27396 18380 27402
rect 18328 27338 18380 27344
rect 18340 27130 18368 27338
rect 18432 27130 18460 28018
rect 18708 27674 18736 28018
rect 18696 27668 18748 27674
rect 18696 27610 18748 27616
rect 19064 27396 19116 27402
rect 19064 27338 19116 27344
rect 18328 27124 18380 27130
rect 18328 27066 18380 27072
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18788 27056 18840 27062
rect 19076 27033 19104 27338
rect 19168 27334 19196 28018
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19156 27328 19208 27334
rect 19156 27270 19208 27276
rect 18788 26998 18840 27004
rect 19062 27024 19118 27033
rect 18420 26920 18472 26926
rect 18420 26862 18472 26868
rect 18432 26042 18460 26862
rect 18708 26518 18736 26998
rect 18800 26897 18828 26998
rect 19062 26959 19118 26968
rect 18786 26888 18842 26897
rect 18786 26823 18842 26832
rect 19168 26790 19196 27270
rect 19156 26784 19208 26790
rect 19156 26726 19208 26732
rect 18696 26512 18748 26518
rect 18696 26454 18748 26460
rect 18420 26036 18472 26042
rect 18420 25978 18472 25984
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 17316 25764 17368 25770
rect 17316 25706 17368 25712
rect 17328 25498 17356 25706
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17592 25696 17644 25702
rect 17592 25638 17644 25644
rect 17512 25498 17540 25638
rect 17604 25498 17632 25638
rect 17316 25492 17368 25498
rect 17316 25434 17368 25440
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17960 24268 18012 24274
rect 17960 24210 18012 24216
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17132 23860 17184 23866
rect 17132 23802 17184 23808
rect 16764 23588 16816 23594
rect 16764 23530 16816 23536
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15764 23050 15792 23462
rect 16776 23322 16804 23530
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15580 21894 15608 22374
rect 16580 22024 16632 22030
rect 16578 21992 16580 22001
rect 16632 21992 16634 22001
rect 16578 21927 16634 21936
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15568 21888 15620 21894
rect 15568 21830 15620 21836
rect 15752 21888 15804 21894
rect 15752 21830 15804 21836
rect 15016 21616 15068 21622
rect 15016 21558 15068 21564
rect 15120 21554 15148 21830
rect 15580 21690 15608 21830
rect 15764 21690 15792 21830
rect 16592 21690 16620 21927
rect 15292 21684 15344 21690
rect 15568 21684 15620 21690
rect 15344 21644 15516 21672
rect 15292 21626 15344 21632
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15200 21412 15252 21418
rect 15200 21354 15252 21360
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14936 20942 14964 21286
rect 15108 21072 15160 21078
rect 15108 21014 15160 21020
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14660 20058 14688 20198
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14752 19854 14780 20266
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14476 18766 14504 19314
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14464 18760 14516 18766
rect 14464 18702 14516 18708
rect 14476 18426 14504 18702
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 17814 14320 18158
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13740 15706 13768 16662
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13740 15570 13768 15642
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13832 15502 13860 16730
rect 14108 15910 14136 17478
rect 14292 17202 14320 17750
rect 14568 17678 14596 18838
rect 14752 18834 14780 19790
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14936 18630 14964 19790
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14660 17202 14688 18566
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17678 14872 17818
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14292 16794 14320 17138
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 16794 14504 16934
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14660 16708 14688 17138
rect 14568 16680 14688 16708
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 16250 14320 16526
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14568 15570 14596 16680
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14660 16250 14688 16390
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14752 16130 14780 17546
rect 14936 17202 14964 18566
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 14660 16114 14780 16130
rect 14648 16108 14780 16114
rect 14700 16102 14780 16108
rect 14648 16050 14700 16056
rect 14936 15706 14964 17138
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14550 13768 14826
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13832 14074 13860 15438
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13924 14958 13952 15302
rect 14752 15162 14780 15438
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14414 13952 14894
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14618 14136 14758
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 14108 14074 14136 14554
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14476 14006 14504 14962
rect 14936 14550 14964 15302
rect 15028 14958 15056 20402
rect 15120 20398 15148 21014
rect 15212 20754 15240 21354
rect 15304 20942 15332 21354
rect 15488 21350 15516 21644
rect 15568 21626 15620 21632
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 15580 21554 15608 21626
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15396 20754 15424 20810
rect 15672 20806 15700 21422
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 15212 20726 15424 20754
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 15212 20058 15240 20538
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15856 19854 15884 20742
rect 16592 20602 16620 20878
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15120 18766 15148 19450
rect 15396 18766 15424 19722
rect 15580 19514 15608 19790
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15488 18834 15516 19246
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 16132 18766 16160 19790
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16316 19514 16344 19654
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16224 19394 16252 19450
rect 16672 19440 16724 19446
rect 16670 19408 16672 19417
rect 16724 19408 16726 19417
rect 16224 19378 16436 19394
rect 16224 19372 16448 19378
rect 16224 19366 16396 19372
rect 16670 19343 16726 19352
rect 16396 19314 16448 19320
rect 16776 18766 16804 21286
rect 16868 20874 16896 22510
rect 17144 22166 17172 23802
rect 17328 23186 17356 24142
rect 17972 23322 18000 24210
rect 18432 23662 18460 25842
rect 19168 25838 19196 26726
rect 19352 26042 19380 27950
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19536 27130 19564 27406
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19340 26036 19392 26042
rect 19340 25978 19392 25984
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19156 25832 19208 25838
rect 19156 25774 19208 25780
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 19076 24954 19104 25094
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 19076 24818 19104 24890
rect 19168 24818 19196 25774
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 18892 24410 18920 24754
rect 19260 24682 19288 25842
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18892 23798 18920 24074
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19168 23866 19196 24006
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 18880 23792 18932 23798
rect 18880 23734 18932 23740
rect 18972 23792 19024 23798
rect 18972 23734 19024 23740
rect 18420 23656 18472 23662
rect 18420 23598 18472 23604
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17328 22574 17356 23122
rect 18248 23118 18276 23462
rect 18984 23118 19012 23734
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18236 23112 18288 23118
rect 18236 23054 18288 23060
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17972 22778 18000 22918
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 18156 22234 18184 23054
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 22710 18644 22918
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 19076 22438 19104 23462
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 17132 22160 17184 22166
rect 17132 22102 17184 22108
rect 17040 21344 17092 21350
rect 17144 21332 17172 22102
rect 17512 21554 17540 22170
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17092 21304 17172 21332
rect 17040 21286 17092 21292
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16868 20398 16896 20810
rect 17316 20800 17368 20806
rect 17420 20754 17448 21490
rect 17684 21140 17736 21146
rect 17788 21128 17816 21490
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17736 21100 17816 21128
rect 17684 21082 17736 21088
rect 17368 20748 17448 20754
rect 17316 20742 17448 20748
rect 17328 20726 17448 20742
rect 17420 20398 17448 20726
rect 17788 20398 17816 21100
rect 17972 20942 18000 21286
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18708 20874 18736 21898
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18708 20777 18736 20810
rect 18694 20768 18750 20777
rect 18694 20703 18750 20712
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 17408 20392 17460 20398
rect 17500 20392 17552 20398
rect 17408 20334 17460 20340
rect 17498 20360 17500 20369
rect 17776 20392 17828 20398
rect 17552 20360 17554 20369
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 15396 18290 15424 18702
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 16132 18086 16160 18702
rect 16316 18426 16344 18702
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16776 18358 16804 18702
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16776 18154 16804 18294
rect 17420 18154 17448 20334
rect 17554 20318 17724 20346
rect 17776 20334 17828 20340
rect 17498 20295 17554 20304
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17604 18766 17632 19926
rect 17696 19446 17724 20318
rect 17788 19854 17816 20334
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 20058 17908 20198
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17684 19440 17736 19446
rect 17684 19382 17736 19388
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17338 15148 17614
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16040 16250 16068 16458
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16132 16114 16160 18022
rect 17696 17678 17724 19382
rect 17972 18970 18000 20402
rect 18064 20262 18092 20402
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18156 18766 18184 19110
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17788 18426 17816 18702
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 18156 18222 18184 18566
rect 18340 18358 18368 18566
rect 18328 18352 18380 18358
rect 18328 18294 18380 18300
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 17066 17080 17478
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 14832 14340 14884 14346
rect 14832 14282 14884 14288
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13832 13530 13860 13874
rect 14016 13530 14044 13874
rect 14476 13530 14504 13942
rect 14568 13870 14596 14214
rect 14844 13870 14872 14282
rect 14936 14074 14964 14486
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15028 13938 15056 14894
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 13740 13326 13768 13466
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 14476 13190 14504 13466
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14568 12986 14596 13670
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12442 13768 12718
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 14844 11218 14872 13670
rect 15120 12434 15148 16050
rect 16960 15502 16988 17002
rect 17052 16046 17080 17002
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16960 15026 16988 15438
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16684 14618 16712 14894
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15212 14414 15240 14486
rect 16960 14482 16988 14962
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15752 14408 15804 14414
rect 16120 14408 16172 14414
rect 15804 14368 16120 14396
rect 15752 14350 15804 14356
rect 16120 14350 16172 14356
rect 15212 13938 15240 14350
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 14074 15700 14214
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 14936 12406 15148 12434
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 10606 13584 11086
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13924 10266 13952 10474
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12728 9722 12756 9998
rect 12440 9716 12492 9722
rect 12716 9716 12768 9722
rect 12492 9676 12572 9704
rect 12440 9658 12492 9664
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 12268 8974 12296 9454
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 10980 800 11008 8774
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 8090 11928 8366
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 12544 7868 12572 9676
rect 12716 9658 12768 9664
rect 14016 9586 14044 10950
rect 14292 10674 14320 10950
rect 14384 10674 14412 11154
rect 14844 11014 14872 11154
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14660 10266 14688 10610
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12636 8090 12664 8502
rect 14292 8362 14320 9930
rect 14936 9586 14964 12406
rect 15488 12322 15516 12582
rect 15304 12306 15516 12322
rect 15292 12300 15516 12306
rect 15344 12294 15516 12300
rect 15292 12242 15344 12248
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8566 14412 9318
rect 14568 9178 14596 9386
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 14752 8430 14780 8842
rect 15028 8634 15056 12174
rect 16132 11354 16160 14350
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16316 11898 16344 12106
rect 16684 11898 16712 12786
rect 16868 12442 16896 12786
rect 16856 12436 16908 12442
rect 17052 12434 17080 15982
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17144 14958 17172 15506
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17144 14414 17172 14894
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 12986 17172 14350
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 14006 17356 14282
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17236 12714 17264 13262
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17052 12406 17356 12434
rect 16856 12378 16908 12384
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 17144 11830 17172 12106
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17328 11694 17356 12406
rect 17420 11762 17448 17206
rect 18432 17202 18460 19790
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18524 18970 18552 19314
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18616 18630 18644 19654
rect 18800 18766 18828 21490
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18604 18624 18656 18630
rect 18604 18566 18656 18572
rect 18616 18086 18644 18566
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18800 17678 18828 18702
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18892 17354 18920 21830
rect 19076 20262 19104 22374
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18984 19514 19012 19858
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18800 17338 18920 17354
rect 18800 17332 18932 17338
rect 18800 17326 18880 17332
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17696 16590 17724 16934
rect 17788 16658 17816 16934
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17880 16454 17908 17070
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17880 16182 17908 16390
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 14958 17816 15302
rect 18432 15162 18460 16050
rect 18800 15978 18828 17326
rect 18880 17274 18932 17280
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 16726 18920 17138
rect 18984 16998 19012 19450
rect 19076 19334 19104 20198
rect 19076 19306 19196 19334
rect 19168 18902 19196 19306
rect 19260 19242 19288 24618
rect 19444 23186 19472 25638
rect 19628 24614 19656 31726
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 21548 30048 21600 30054
rect 21548 29990 21600 29996
rect 19996 29646 20024 29990
rect 21560 29646 21588 29990
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 21548 29640 21600 29646
rect 21548 29582 21600 29588
rect 19996 29306 20024 29582
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 19984 29300 20036 29306
rect 19984 29242 20036 29248
rect 19996 28558 20024 29242
rect 20456 28558 20484 29446
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19720 26790 19748 27814
rect 19996 27470 20024 28494
rect 21088 28484 21140 28490
rect 21088 28426 21140 28432
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 21008 28150 21036 28358
rect 20996 28144 21048 28150
rect 20996 28086 21048 28092
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 20916 27674 20944 28018
rect 20904 27668 20956 27674
rect 20904 27610 20956 27616
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19800 27328 19852 27334
rect 19800 27270 19852 27276
rect 19812 26858 19840 27270
rect 19800 26852 19852 26858
rect 19800 26794 19852 26800
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19720 26586 19748 26726
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19996 25702 20024 27406
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20548 27130 20576 27338
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20720 27056 20772 27062
rect 20720 26998 20772 27004
rect 20352 26852 20404 26858
rect 20352 26794 20404 26800
rect 20364 26314 20392 26794
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 20088 25294 20116 25978
rect 20180 25906 20208 26250
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 20180 25158 20208 25842
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 20180 24954 20208 25094
rect 20168 24948 20220 24954
rect 20168 24890 20220 24896
rect 20272 24818 20300 25230
rect 20364 25158 20392 26250
rect 20732 25906 20760 26998
rect 21008 26926 21036 28086
rect 21100 27062 21128 28426
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 22020 28014 22048 28086
rect 22008 28008 22060 28014
rect 22008 27950 22060 27956
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21284 27130 21312 27338
rect 22020 27334 22048 27950
rect 22204 27946 22232 29446
rect 22388 28150 22416 37130
rect 23216 35894 23244 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 23216 35866 23796 35894
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 22376 28144 22428 28150
rect 22376 28086 22428 28092
rect 22652 28144 22704 28150
rect 22652 28086 22704 28092
rect 22192 27940 22244 27946
rect 22192 27882 22244 27888
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21088 27056 21140 27062
rect 21088 26998 21140 27004
rect 22020 26994 22048 27270
rect 22480 27130 22508 27814
rect 22560 27532 22612 27538
rect 22560 27474 22612 27480
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21732 26920 21784 26926
rect 21732 26862 21784 26868
rect 21008 26246 21036 26862
rect 20996 26240 21048 26246
rect 20996 26182 21048 26188
rect 21192 25974 21220 26862
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 21180 25968 21232 25974
rect 21180 25910 21232 25916
rect 20720 25900 20772 25906
rect 20720 25842 20772 25848
rect 20732 25498 20760 25842
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20628 25424 20680 25430
rect 20824 25378 20852 25910
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 20916 25498 20944 25842
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20680 25372 20852 25378
rect 20628 25366 20852 25372
rect 20640 25350 20852 25366
rect 20352 25152 20404 25158
rect 20352 25094 20404 25100
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19628 22778 19656 23666
rect 20088 23662 20116 24006
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19812 23186 19840 23462
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 20088 22574 20116 23598
rect 20364 22642 20392 25094
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20628 23520 20680 23526
rect 20628 23462 20680 23468
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20352 22636 20404 22642
rect 20352 22578 20404 22584
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 22030 19380 22374
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 21146 19748 21286
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19536 20534 19564 20742
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19628 19378 19656 19654
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19248 19236 19300 19242
rect 19248 19178 19300 19184
rect 19156 18896 19208 18902
rect 19156 18838 19208 18844
rect 19168 18290 19196 18838
rect 19720 18834 19748 19314
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19432 18624 19484 18630
rect 19484 18572 19564 18578
rect 19432 18566 19564 18572
rect 19444 18550 19564 18566
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19536 18222 19564 18550
rect 19720 18426 19748 18770
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19536 17678 19564 18158
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16250 19012 16390
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18788 15972 18840 15978
rect 18788 15914 18840 15920
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17604 14618 17632 14894
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17788 14498 17816 14894
rect 17604 14470 17816 14498
rect 17604 14346 17632 14470
rect 17776 14408 17828 14414
rect 17880 14396 17908 14894
rect 17972 14618 18000 14894
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17972 14482 18000 14554
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18616 14414 18644 15030
rect 19156 14884 19208 14890
rect 19156 14826 19208 14832
rect 19168 14414 19196 14826
rect 17828 14368 17908 14396
rect 18236 14408 18288 14414
rect 17776 14350 17828 14356
rect 18236 14350 18288 14356
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19156 14408 19208 14414
rect 19156 14350 19208 14356
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17696 13920 17724 14282
rect 17788 14074 17816 14350
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17776 13932 17828 13938
rect 17696 13892 17776 13920
rect 17776 13874 17828 13880
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17788 13326 17816 13874
rect 18064 13394 18092 13874
rect 18248 13530 18276 14350
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18432 14074 18460 14214
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18800 13938 18828 14214
rect 19076 14074 19104 14350
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 18248 12850 18276 13466
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18432 12442 18460 12650
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11830 17908 12038
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17408 11756 17460 11762
rect 17408 11698 17460 11704
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15396 10810 15424 10950
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15580 10470 15608 11086
rect 16132 10674 16160 11154
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17236 10674 17264 11086
rect 16120 10668 16172 10674
rect 17224 10668 17276 10674
rect 16172 10628 16436 10656
rect 16120 10610 16172 10616
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10062 16344 10406
rect 16408 10266 16436 10628
rect 17224 10610 17276 10616
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 17236 10130 17264 10610
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 9178 15516 9318
rect 15948 9178 15976 9454
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 15488 8362 15516 9114
rect 16776 8634 16804 9862
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 13188 7886 13216 8230
rect 12716 7880 12768 7886
rect 12544 7840 12716 7868
rect 12716 7822 12768 7828
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13464 7818 13492 8298
rect 15488 8090 15516 8298
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15580 7954 15608 8570
rect 16868 8430 16896 10066
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16960 9178 16988 9998
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17224 9172 17276 9178
rect 17328 9160 17356 11630
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17420 10674 17448 11154
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10674 17908 11018
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10742 18092 10950
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 17408 10668 17460 10674
rect 17868 10668 17920 10674
rect 17408 10610 17460 10616
rect 17788 10628 17868 10656
rect 17420 10180 17448 10610
rect 17788 10198 17816 10628
rect 17868 10610 17920 10616
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17880 10266 17908 10474
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 10192 17828 10198
rect 17420 10152 17540 10180
rect 17512 10062 17540 10152
rect 17776 10134 17828 10140
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17276 9132 17356 9160
rect 17224 9114 17276 9120
rect 17236 8430 17264 9114
rect 17512 8838 17540 9998
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17696 8430 17724 8910
rect 17788 8634 17816 8910
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17972 8430 18000 10066
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 8974 18092 9318
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18156 8566 18184 8842
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 800 14228 7686
rect 15856 7546 15884 7754
rect 16684 7546 16712 8230
rect 17144 8090 17172 8366
rect 18156 8362 18184 8502
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 8090 18184 8298
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17144 7546 17172 8026
rect 18340 7818 18368 12378
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18432 10674 18460 11086
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18524 10674 18552 10950
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18432 10062 18460 10610
rect 18524 10130 18552 10610
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 18064 7206 18092 7686
rect 18340 7410 18368 7754
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 800 18092 7142
rect 18708 800 18736 12038
rect 18800 10538 18828 13874
rect 19076 12782 19104 14010
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18984 9178 19012 11494
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19260 2774 19288 16594
rect 19904 16590 19932 22510
rect 20088 22098 20116 22510
rect 20548 22166 20576 22714
rect 20640 22166 20668 23462
rect 20732 22574 20760 24754
rect 20824 22710 20852 25350
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21192 24818 21220 25230
rect 21284 24818 21312 25842
rect 21468 24886 21496 25842
rect 21456 24880 21508 24886
rect 21456 24822 21508 24828
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21192 23322 21220 24754
rect 21468 24614 21496 24822
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 23866 21588 24550
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21180 23316 21232 23322
rect 21180 23258 21232 23264
rect 21192 22778 21220 23258
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21468 22778 21496 22918
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 20628 22160 20680 22166
rect 20628 22102 20680 22108
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 20088 21418 20116 22034
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 20180 20806 20208 21422
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 19996 20534 20024 20742
rect 20640 20602 20668 22102
rect 20732 21894 20760 22510
rect 20824 22234 20852 22646
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20732 21554 20760 21830
rect 20916 21554 20944 22510
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20732 20602 20760 21490
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20628 20596 20680 20602
rect 20628 20538 20680 20544
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 20824 20466 20852 20810
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19996 17746 20024 18158
rect 20272 17814 20300 18226
rect 20456 18086 20484 18634
rect 20548 18426 20576 19110
rect 20640 18970 20668 19314
rect 20824 19174 20852 20402
rect 20916 19446 20944 21490
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21008 20058 21036 21422
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 21100 20602 21128 20810
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20260 17808 20312 17814
rect 20260 17750 20312 17756
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 20640 17610 20668 18906
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20732 17134 20760 18770
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16794 20760 17070
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16250 19656 16390
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19904 15978 19932 16526
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 16182 20760 16390
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 19352 13870 19380 14486
rect 19628 14074 19656 14758
rect 19720 14074 19748 14894
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19628 11762 19656 12038
rect 19720 11830 19748 13194
rect 19812 12850 19840 15914
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 20088 15570 20116 15846
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20088 15026 20116 15506
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 15026 20576 15302
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 19996 14618 20024 14962
rect 20088 14618 20116 14962
rect 20640 14770 20668 15506
rect 20732 15502 20760 16118
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20720 14816 20772 14822
rect 20640 14764 20720 14770
rect 20640 14758 20772 14764
rect 20640 14742 20760 14758
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20640 14278 20668 14742
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20824 13870 20852 19110
rect 20916 18630 20944 19382
rect 21192 19310 21220 21354
rect 21560 21010 21588 23054
rect 21744 22642 21772 26862
rect 22284 26512 22336 26518
rect 22284 26454 22336 26460
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 24410 21864 24550
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21928 24206 21956 25638
rect 22020 24614 22048 26182
rect 22112 25702 22140 26250
rect 22296 25906 22324 26454
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22388 26042 22416 26182
rect 22572 26058 22600 27474
rect 22664 27130 22692 28086
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22848 27674 22876 28018
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 23492 27470 23520 27882
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22836 27328 22888 27334
rect 22836 27270 22888 27276
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 22756 26790 22784 27270
rect 22848 26994 22876 27270
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 23388 26784 23440 26790
rect 23388 26726 23440 26732
rect 22756 26450 22784 26726
rect 22744 26444 22796 26450
rect 22744 26386 22796 26392
rect 22376 26036 22428 26042
rect 22572 26030 22692 26058
rect 22376 25978 22428 25984
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22112 25498 22140 25638
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 24750 22140 25230
rect 22296 24886 22324 25842
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22388 25498 22416 25638
rect 22572 25498 22600 25842
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22572 24954 22600 25434
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22284 24880 22336 24886
rect 22284 24822 22336 24828
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21744 21434 21772 22578
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 21928 21622 21956 21830
rect 22020 21690 22048 24550
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22388 23662 22416 24006
rect 22664 23730 22692 26030
rect 22756 25294 22784 26386
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 22928 26240 22980 26246
rect 22928 26182 22980 26188
rect 22940 25294 22968 26182
rect 23308 26042 23336 26318
rect 23400 26246 23428 26726
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23572 26240 23624 26246
rect 23572 26182 23624 26188
rect 23296 26036 23348 26042
rect 23296 25978 23348 25984
rect 23308 25294 23336 25978
rect 23400 25974 23428 26182
rect 23584 25974 23612 26182
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 23400 25498 23428 25910
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23400 24410 23428 24754
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22100 23044 22152 23050
rect 22100 22986 22152 22992
rect 22284 23044 22336 23050
rect 22284 22986 22336 22992
rect 22112 22234 22140 22986
rect 22296 22778 22324 22986
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21916 21616 21968 21622
rect 21916 21558 21968 21564
rect 21744 21406 21956 21434
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21192 18698 21220 19246
rect 21836 18834 21864 19314
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20916 18358 20944 18566
rect 20904 18352 20956 18358
rect 20904 18294 20956 18300
rect 20916 17610 20944 18294
rect 21100 18154 21128 18566
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14618 21128 14758
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 12986 21036 13670
rect 21100 13394 21128 13874
rect 21284 13870 21312 15370
rect 21376 14822 21404 17818
rect 21560 17610 21588 18634
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21744 18222 21772 18566
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21468 16794 21496 17138
rect 21652 16810 21680 17750
rect 21744 17678 21772 18158
rect 21836 17814 21864 18770
rect 21928 17898 21956 21406
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 19990 22140 20334
rect 22204 20330 22232 22442
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 19378 22140 19926
rect 22388 19514 22416 23598
rect 22664 22778 22692 23666
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 22030 22508 22374
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22664 20942 22692 22510
rect 22848 21690 22876 22578
rect 23032 22098 23060 24074
rect 23768 23866 23796 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23952 27130 23980 27406
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 23952 25906 23980 27066
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 28908 26308 28960 26314
rect 28908 26250 28960 26256
rect 26976 26240 27028 26246
rect 26976 26182 27028 26188
rect 28264 26240 28316 26246
rect 28264 26182 28316 26188
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25294 25176 25774
rect 26988 25294 27016 26182
rect 28276 25702 28304 26182
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28264 25696 28316 25702
rect 28264 25638 28316 25644
rect 28080 25424 28132 25430
rect 28080 25366 28132 25372
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 25148 24614 25176 25230
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 25700 24954 25728 25162
rect 26436 24954 26464 25162
rect 25688 24948 25740 24954
rect 25688 24890 25740 24896
rect 26424 24948 26476 24954
rect 26424 24890 26476 24896
rect 26148 24812 26200 24818
rect 26148 24754 26200 24760
rect 24308 24608 24360 24614
rect 24308 24550 24360 24556
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 24320 24206 24348 24550
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 24320 23186 24348 24142
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24688 23866 24716 24074
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 25148 23730 25176 24210
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 24308 23180 24360 23186
rect 24308 23122 24360 23128
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23400 22642 23428 22986
rect 24596 22778 24624 23462
rect 25148 23066 25176 23666
rect 25240 23322 25268 24550
rect 25424 24138 25452 24550
rect 26160 24410 26188 24754
rect 26148 24404 26200 24410
rect 26148 24346 26200 24352
rect 26988 24274 27016 25230
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27172 24682 27200 25094
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27172 24410 27200 24618
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 26976 24268 27028 24274
rect 26976 24210 27028 24216
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 25412 24132 25464 24138
rect 25412 24074 25464 24080
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 26068 23662 26096 24006
rect 26424 23724 26476 23730
rect 26424 23666 26476 23672
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 25872 23588 25924 23594
rect 25872 23530 25924 23536
rect 25884 23322 25912 23530
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 25872 23316 25924 23322
rect 25872 23258 25924 23264
rect 25240 23225 25268 23258
rect 25226 23216 25282 23225
rect 25226 23151 25282 23160
rect 25148 23038 25268 23066
rect 25240 22982 25268 23038
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 23388 22636 23440 22642
rect 23388 22578 23440 22584
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 24032 22432 24084 22438
rect 24032 22374 24084 22380
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22572 20466 22600 20878
rect 23308 20534 23336 22374
rect 23768 22098 23796 22374
rect 23756 22092 23808 22098
rect 23756 22034 23808 22040
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23400 20874 23428 21286
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23584 20466 23612 21966
rect 23940 21888 23992 21894
rect 23940 21830 23992 21836
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22480 19281 22508 20334
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 22848 19922 22876 20266
rect 23400 19990 23428 20266
rect 23492 20058 23520 20402
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23388 19984 23440 19990
rect 23388 19926 23440 19932
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22848 19378 22876 19858
rect 23584 19417 23612 20198
rect 23570 19408 23626 19417
rect 22836 19372 22888 19378
rect 23570 19343 23626 19352
rect 22836 19314 22888 19320
rect 22466 19272 22522 19281
rect 22466 19207 22522 19216
rect 22480 18970 22508 19207
rect 22848 18970 22876 19314
rect 23584 19258 23612 19343
rect 23492 19230 23612 19258
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 23216 18766 23244 19110
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23216 18630 23244 18702
rect 23204 18624 23256 18630
rect 23204 18566 23256 18572
rect 23308 18426 23336 19110
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23492 18154 23520 19230
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 21928 17882 22324 17898
rect 21928 17876 22336 17882
rect 21928 17870 22284 17876
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21732 17672 21784 17678
rect 21732 17614 21784 17620
rect 21732 17536 21784 17542
rect 21928 17524 21956 17870
rect 22284 17818 22336 17824
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 21784 17496 21956 17524
rect 21732 17478 21784 17484
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21652 16794 21772 16810
rect 21456 16788 21508 16794
rect 21652 16788 21784 16794
rect 21652 16782 21732 16788
rect 21456 16730 21508 16736
rect 21732 16730 21784 16736
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21560 15366 21588 15846
rect 21548 15360 21600 15366
rect 21548 15302 21600 15308
rect 21560 15026 21588 15302
rect 21836 15162 21864 17070
rect 22020 16658 22048 17546
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23296 17536 23348 17542
rect 23296 17478 23348 17484
rect 22204 16658 22232 17478
rect 22756 17338 22784 17478
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 22020 16182 22048 16594
rect 23032 16590 23060 17478
rect 23216 17202 23244 17478
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23308 17134 23336 17478
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21560 14482 21588 14962
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 19800 12708 19852 12714
rect 19800 12650 19852 12656
rect 19812 11830 19840 12650
rect 20548 12238 20576 12786
rect 20824 12714 20852 12786
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20732 12238 20760 12378
rect 20824 12238 20852 12650
rect 21100 12646 21128 13330
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 21008 12306 21036 12582
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20536 12232 20588 12238
rect 19982 12200 20038 12209
rect 20536 12174 20588 12180
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 19982 12135 20038 12144
rect 19708 11824 19760 11830
rect 19708 11766 19760 11772
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19996 11762 20024 12135
rect 20732 11898 20760 12174
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20824 11830 20852 12038
rect 20916 11898 20944 12174
rect 21008 11898 21036 12242
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20996 11892 21048 11898
rect 21100 11880 21128 12582
rect 21180 11892 21232 11898
rect 21100 11852 21180 11880
rect 20996 11834 21048 11840
rect 21180 11834 21232 11840
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 9586 19932 10406
rect 19996 9994 20024 11698
rect 21284 10266 21312 13262
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21376 12442 21404 12786
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11558 21496 12038
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21652 10266 21680 10406
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21836 10130 21864 15098
rect 22112 15094 22140 15506
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22112 14346 22140 15030
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14414 22324 14758
rect 22480 14618 22508 16390
rect 22572 15978 22600 16526
rect 22560 15972 22612 15978
rect 22560 15914 22612 15920
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22100 14340 22152 14346
rect 22100 14282 22152 14288
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22204 13938 22232 14214
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22388 13530 22416 14350
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22572 13326 22600 15914
rect 23216 14890 23244 16934
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 23308 14929 23336 16458
rect 23584 15502 23612 19110
rect 23676 18426 23704 21558
rect 23952 21554 23980 21830
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23768 17898 23796 20742
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23860 18970 23888 20402
rect 24044 19514 24072 22374
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 24412 21486 24440 22102
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21554 24532 21830
rect 24492 21548 24544 21554
rect 24492 21490 24544 21496
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 20534 24164 21286
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 19786 24164 20470
rect 24780 20262 24808 21490
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24780 19922 24808 20198
rect 24872 19990 24900 20402
rect 25044 20256 25096 20262
rect 25044 20198 25096 20204
rect 25056 20058 25084 20198
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24032 19508 24084 19514
rect 23952 19468 24032 19496
rect 23952 19378 23980 19468
rect 24032 19450 24084 19456
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 23940 19168 23992 19174
rect 23940 19110 23992 19116
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23952 18426 23980 19110
rect 24044 18970 24072 19246
rect 24032 18964 24084 18970
rect 24032 18906 24084 18912
rect 24136 18834 24164 19314
rect 24860 18896 24912 18902
rect 24860 18838 24912 18844
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 24872 18358 24900 18838
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 23768 17870 23888 17898
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23768 17338 23796 17682
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23662 16552 23718 16561
rect 23662 16487 23718 16496
rect 23676 16182 23704 16487
rect 23664 16176 23716 16182
rect 23664 16118 23716 16124
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 23768 15570 23796 16050
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23584 15094 23612 15438
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23572 14952 23624 14958
rect 23294 14920 23350 14929
rect 23204 14884 23256 14890
rect 23572 14894 23624 14900
rect 23294 14855 23350 14864
rect 23204 14826 23256 14832
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22756 13326 22784 14282
rect 23032 13938 23060 14350
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 22112 12458 22140 13262
rect 22572 12986 22600 13262
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 22020 12430 22140 12458
rect 22756 12442 22784 12786
rect 22744 12436 22796 12442
rect 22020 12374 22048 12430
rect 22848 12434 22876 13262
rect 22940 12986 22968 13262
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 22928 12436 22980 12442
rect 22848 12406 22928 12434
rect 22744 12378 22796 12384
rect 22928 12378 22980 12384
rect 22008 12368 22060 12374
rect 23032 12322 23060 13874
rect 23124 13530 23152 13874
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 22008 12310 22060 12316
rect 22940 12294 23060 12322
rect 22836 12232 22888 12238
rect 22940 12209 22968 12294
rect 23124 12238 23152 13262
rect 23112 12232 23164 12238
rect 22836 12174 22888 12180
rect 22926 12200 22982 12209
rect 22848 11082 22876 12174
rect 23112 12174 23164 12180
rect 22926 12135 22982 12144
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22296 10674 22324 10950
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22756 10606 22784 10950
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22756 10266 22784 10542
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19720 9178 19748 9522
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 9178 20116 9318
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19720 8090 19748 8366
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 20272 7886 20300 9046
rect 21008 8838 21036 9998
rect 21100 9042 21128 9998
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21100 8498 21128 8978
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 21100 7818 21128 8434
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21284 7750 21312 8774
rect 21836 8498 21864 10066
rect 23216 10010 23244 14826
rect 23308 14482 23336 14855
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 14074 23336 14214
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23296 12096 23348 12102
rect 23492 12050 23520 14418
rect 23584 14074 23612 14894
rect 23768 14822 23796 15506
rect 23860 15502 23888 17870
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24044 17338 24072 17614
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24872 17066 24900 18294
rect 25240 17882 25268 22918
rect 25320 22636 25372 22642
rect 25320 22578 25372 22584
rect 25332 21146 25360 22578
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25332 20466 25360 20878
rect 25412 20800 25464 20806
rect 25412 20742 25464 20748
rect 25424 20602 25452 20742
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 20466 25544 21082
rect 25792 21026 25820 22510
rect 25976 22234 26004 22510
rect 25964 22228 26016 22234
rect 25964 22170 26016 22176
rect 26068 21554 26096 23598
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 23254 26188 23462
rect 26148 23248 26200 23254
rect 26148 23190 26200 23196
rect 26436 22778 26464 23666
rect 27264 23662 27292 24210
rect 27540 24206 27568 24890
rect 28092 24818 28120 25366
rect 28276 24818 28304 25638
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 27252 23656 27304 23662
rect 27252 23598 27304 23604
rect 26516 22976 26568 22982
rect 26516 22918 26568 22924
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26528 22642 26556 22918
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 26528 22030 26556 22578
rect 27080 22098 27108 22578
rect 27068 22092 27120 22098
rect 27264 22094 27292 23598
rect 27540 23322 27568 24142
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 28000 23594 28028 24006
rect 28092 23730 28120 24142
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 27988 23588 28040 23594
rect 27988 23530 28040 23536
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27540 23118 27568 23258
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27436 22976 27488 22982
rect 27620 22976 27672 22982
rect 27436 22918 27488 22924
rect 27540 22924 27620 22930
rect 27540 22918 27672 22924
rect 27448 22778 27476 22918
rect 27540 22902 27660 22918
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27540 22642 27568 22902
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27264 22066 27568 22094
rect 27068 22034 27120 22040
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25884 21146 25912 21286
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 25792 20998 25912 21026
rect 26068 21010 26096 21490
rect 26528 21486 26556 21966
rect 26516 21480 26568 21486
rect 26516 21422 26568 21428
rect 25688 20936 25740 20942
rect 25688 20878 25740 20884
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25412 20324 25464 20330
rect 25412 20266 25464 20272
rect 25424 19378 25452 20266
rect 25608 19854 25636 20810
rect 25700 20466 25728 20878
rect 25780 20868 25832 20874
rect 25780 20810 25832 20816
rect 25792 20602 25820 20810
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25700 19514 25728 20402
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25332 18426 25360 19314
rect 25424 18970 25452 19314
rect 25884 19310 25912 20998
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25412 18692 25464 18698
rect 25412 18634 25464 18640
rect 25320 18420 25372 18426
rect 25320 18362 25372 18368
rect 25424 18170 25452 18634
rect 25884 18222 25912 19246
rect 26068 18902 26096 20742
rect 26344 20466 26372 20742
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26148 20324 26200 20330
rect 26148 20266 26200 20272
rect 26160 19854 26188 20266
rect 26344 19854 26372 20402
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 26976 20256 27028 20262
rect 26976 20198 27028 20204
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 26804 19854 26832 20198
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26988 19378 27016 20198
rect 27448 19854 27476 20198
rect 27540 19990 27568 22066
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 27632 21078 27660 21286
rect 27620 21072 27672 21078
rect 27620 21014 27672 21020
rect 27632 20466 27660 21014
rect 28000 20942 28028 23530
rect 28184 23322 28212 24074
rect 28368 24070 28396 25842
rect 28448 24948 28500 24954
rect 28448 24890 28500 24896
rect 28460 24614 28488 24890
rect 28920 24818 28948 26250
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 30564 26240 30616 26246
rect 30564 26182 30616 26188
rect 29196 25906 29224 26182
rect 30576 26042 30604 26182
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30564 26036 30616 26042
rect 30564 25978 30616 25984
rect 35440 26036 35492 26042
rect 35440 25978 35492 25984
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 29736 25832 29788 25838
rect 29736 25774 29788 25780
rect 29748 25498 29776 25774
rect 29736 25492 29788 25498
rect 29736 25434 29788 25440
rect 29552 25288 29604 25294
rect 29552 25230 29604 25236
rect 29564 24954 29592 25230
rect 29552 24948 29604 24954
rect 29552 24890 29604 24896
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28448 24608 28500 24614
rect 28448 24550 28500 24556
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28828 24274 28856 24550
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28356 24064 28408 24070
rect 28356 24006 28408 24012
rect 28632 24064 28684 24070
rect 28632 24006 28684 24012
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 28368 23202 28396 24006
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 28276 23174 28396 23202
rect 28184 22778 28212 23122
rect 28276 23050 28304 23174
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 28368 22778 28396 23054
rect 28460 22778 28488 23054
rect 28644 23050 28672 24006
rect 28828 23866 28856 24210
rect 28920 24206 28948 24754
rect 29000 24676 29052 24682
rect 29000 24618 29052 24624
rect 29012 24410 29040 24618
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 30392 24274 30420 25978
rect 30472 25968 30524 25974
rect 35452 25945 35480 25978
rect 30472 25910 30524 25916
rect 35438 25936 35494 25945
rect 30484 25498 30512 25910
rect 35438 25871 35494 25880
rect 33324 25832 33376 25838
rect 33324 25774 33376 25780
rect 31208 25696 31260 25702
rect 31208 25638 31260 25644
rect 30472 25492 30524 25498
rect 30472 25434 30524 25440
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30564 24880 30616 24886
rect 30564 24822 30616 24828
rect 30472 24812 30524 24818
rect 30472 24754 30524 24760
rect 29460 24268 29512 24274
rect 29460 24210 29512 24216
rect 30380 24268 30432 24274
rect 30380 24210 30432 24216
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28920 23866 28948 24006
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28828 23118 28856 23462
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28632 23044 28684 23050
rect 28632 22986 28684 22992
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 28356 22772 28408 22778
rect 28356 22714 28408 22720
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 28644 22012 28672 22986
rect 28920 22642 28948 23122
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 29368 22976 29420 22982
rect 29368 22918 29420 22924
rect 28908 22636 28960 22642
rect 28908 22578 28960 22584
rect 28724 22568 28776 22574
rect 28776 22528 28856 22556
rect 28724 22510 28776 22516
rect 28724 22024 28776 22030
rect 28644 21984 28724 22012
rect 28724 21966 28776 21972
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28460 20942 28488 21082
rect 28552 21078 28580 21830
rect 28632 21616 28684 21622
rect 28828 21604 28856 22528
rect 28908 22500 28960 22506
rect 28908 22442 28960 22448
rect 28920 22098 28948 22442
rect 28908 22092 28960 22098
rect 29104 22094 29132 22918
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 29196 22234 29224 22578
rect 29380 22574 29408 22918
rect 29472 22642 29500 24210
rect 30484 24206 30512 24754
rect 30472 24200 30524 24206
rect 30472 24142 30524 24148
rect 30288 24064 30340 24070
rect 30288 24006 30340 24012
rect 30472 24064 30524 24070
rect 30472 24006 30524 24012
rect 30300 23866 30328 24006
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 29736 23180 29788 23186
rect 29736 23122 29788 23128
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29564 22778 29592 22918
rect 29552 22772 29604 22778
rect 29552 22714 29604 22720
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29368 22568 29420 22574
rect 29368 22510 29420 22516
rect 29184 22228 29236 22234
rect 29184 22170 29236 22176
rect 29104 22066 29316 22094
rect 28908 22034 28960 22040
rect 29288 22030 29316 22066
rect 29748 22030 29776 23122
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 29920 22568 29972 22574
rect 29920 22510 29972 22516
rect 29932 22438 29960 22510
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29932 22166 29960 22374
rect 29920 22160 29972 22166
rect 29920 22102 29972 22108
rect 30208 22094 30236 22578
rect 30300 22234 30328 22578
rect 30392 22234 30420 22578
rect 30288 22228 30340 22234
rect 30288 22170 30340 22176
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30024 22066 30236 22094
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29736 22024 29788 22030
rect 29736 21966 29788 21972
rect 29276 21888 29328 21894
rect 29276 21830 29328 21836
rect 28684 21576 28856 21604
rect 28632 21558 28684 21564
rect 28540 21072 28592 21078
rect 28540 21014 28592 21020
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28540 20936 28592 20942
rect 28644 20924 28672 21558
rect 28828 21078 28856 21576
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28592 20896 28672 20924
rect 28724 20936 28776 20942
rect 28540 20878 28592 20884
rect 28724 20878 28776 20884
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 27724 20602 27752 20742
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27528 19984 27580 19990
rect 27528 19926 27580 19932
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27068 19712 27120 19718
rect 27068 19654 27120 19660
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26056 18896 26108 18902
rect 26056 18838 26108 18844
rect 25332 18154 25452 18170
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25320 18148 25452 18154
rect 25372 18142 25452 18148
rect 25320 18090 25372 18096
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25332 17678 25360 18090
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25700 17202 25728 17682
rect 25792 17202 25820 17818
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 24860 17060 24912 17066
rect 24860 17002 24912 17008
rect 24676 16584 24728 16590
rect 24674 16552 24676 16561
rect 24728 16552 24730 16561
rect 26068 16522 26096 18838
rect 27080 18766 27108 19654
rect 27540 19292 27568 19926
rect 27724 19922 27752 20538
rect 28000 20398 28028 20878
rect 28356 20868 28408 20874
rect 28356 20810 28408 20816
rect 28368 20602 28396 20810
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 27988 20392 28040 20398
rect 27988 20334 28040 20340
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 28460 19854 28488 20878
rect 28632 20800 28684 20806
rect 28736 20754 28764 20878
rect 28684 20748 28764 20754
rect 28632 20742 28764 20748
rect 28644 20726 28764 20742
rect 28736 20602 28764 20726
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 29288 20466 29316 21830
rect 30024 20466 30052 22066
rect 30380 21888 30432 21894
rect 30380 21830 30432 21836
rect 30392 21690 30420 21830
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 30392 21146 30420 21626
rect 30380 21140 30432 21146
rect 30380 21082 30432 21088
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30116 20466 30144 20878
rect 30288 20868 30340 20874
rect 30288 20810 30340 20816
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29276 20460 29328 20466
rect 29276 20402 29328 20408
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 29012 19786 29040 20402
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 29104 19718 29132 20402
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29736 20256 29788 20262
rect 29736 20198 29788 20204
rect 29656 20058 29684 20198
rect 29644 20052 29696 20058
rect 29644 19994 29696 20000
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 29092 19712 29144 19718
rect 29092 19654 29144 19660
rect 27724 19310 27752 19654
rect 28722 19408 28778 19417
rect 28722 19343 28778 19352
rect 27712 19304 27764 19310
rect 27540 19281 27660 19292
rect 27540 19272 27674 19281
rect 27540 19264 27618 19272
rect 27712 19246 27764 19252
rect 27618 19207 27674 19216
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27540 18834 27568 19110
rect 27528 18828 27580 18834
rect 27528 18770 27580 18776
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26160 18426 26188 18634
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 26608 18080 26660 18086
rect 26608 18022 26660 18028
rect 26620 17610 26648 18022
rect 26608 17604 26660 17610
rect 26608 17546 26660 17552
rect 24674 16487 24730 16496
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25424 16182 25452 16390
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 24860 15904 24912 15910
rect 24860 15846 24912 15852
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23756 14816 23808 14822
rect 23756 14758 23808 14764
rect 23768 14278 23796 14758
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23676 14074 23704 14214
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23768 13938 23796 14214
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 23756 12232 23808 12238
rect 23754 12200 23756 12209
rect 23808 12200 23810 12209
rect 23754 12135 23810 12144
rect 23296 12038 23348 12044
rect 23308 11354 23336 12038
rect 23400 12022 23520 12050
rect 23400 11354 23428 12022
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23400 11218 23428 11290
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23400 10538 23428 11018
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 22192 9988 22244 9994
rect 23216 9982 23428 10010
rect 23952 9994 23980 15846
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24412 14414 24440 15438
rect 24872 14414 24900 15846
rect 24400 14408 24452 14414
rect 24320 14368 24400 14396
rect 24320 13462 24348 14368
rect 24400 14350 24452 14356
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 25424 14362 25452 16118
rect 25872 16040 25924 16046
rect 25872 15982 25924 15988
rect 25504 15904 25556 15910
rect 25556 15852 25636 15858
rect 25504 15846 25636 15852
rect 25516 15830 25636 15846
rect 25608 15366 25636 15830
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25608 15026 25636 15302
rect 25884 15162 25912 15982
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25504 14408 25556 14414
rect 25424 14356 25504 14362
rect 25424 14350 25556 14356
rect 25424 14334 25544 14350
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24308 13456 24360 13462
rect 24308 13398 24360 13404
rect 24320 12918 24348 13398
rect 24964 13394 24992 13670
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24952 13388 25004 13394
rect 24952 13330 25004 13336
rect 24308 12912 24360 12918
rect 24308 12854 24360 12860
rect 24412 11354 24440 13330
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12986 24808 13262
rect 24964 12986 24992 13330
rect 25136 13184 25188 13190
rect 25136 13126 25188 13132
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25148 12850 25176 13126
rect 25228 12912 25280 12918
rect 25228 12854 25280 12860
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 25136 12844 25188 12850
rect 25136 12786 25188 12792
rect 24780 12434 24808 12786
rect 25044 12640 25096 12646
rect 25044 12582 25096 12588
rect 24780 12406 24900 12434
rect 24872 11762 24900 12406
rect 25056 12306 25084 12582
rect 25044 12300 25096 12306
rect 25044 12242 25096 12248
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 22192 9930 22244 9936
rect 22204 9722 22232 9930
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 23308 9586 23336 9862
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21468 8090 21496 8434
rect 22020 8430 22048 9522
rect 23032 9042 23060 9522
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 22112 7954 22140 8978
rect 23204 8832 23256 8838
rect 23204 8774 23256 8780
rect 23216 8634 23244 8774
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 19260 2746 19380 2774
rect 19352 800 19380 2746
rect 21284 800 21312 7686
rect 23308 2774 23336 9522
rect 23400 8922 23428 9982
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23952 9586 23980 9930
rect 24044 9722 24072 10474
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24320 9674 24348 11290
rect 25240 11218 25268 12854
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24688 10810 24716 11086
rect 24780 10810 24808 11154
rect 25228 11076 25280 11082
rect 25228 11018 25280 11024
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 25240 10674 25268 11018
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 24320 9646 24532 9674
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24504 9042 24532 9646
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 25148 8974 25176 9862
rect 25240 9110 25268 10610
rect 25332 10062 25360 12242
rect 25424 12102 25452 14334
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25608 13802 25636 13874
rect 25596 13796 25648 13802
rect 25596 13738 25648 13744
rect 25504 13728 25556 13734
rect 25504 13670 25556 13676
rect 25516 12850 25544 13670
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25504 12844 25556 12850
rect 25504 12786 25556 12792
rect 25504 12436 25556 12442
rect 25608 12434 25636 12922
rect 25700 12918 25728 13126
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 25872 12708 25924 12714
rect 25872 12650 25924 12656
rect 25556 12406 25636 12434
rect 25504 12378 25556 12384
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25412 11620 25464 11626
rect 25412 11562 25464 11568
rect 25424 10674 25452 11562
rect 25516 10674 25544 12378
rect 25884 12170 25912 12650
rect 25976 12238 26004 12718
rect 26068 12442 26096 16458
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 14618 26188 16390
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26436 15162 26464 16050
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 26896 14414 26924 14554
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 26988 13802 27016 18702
rect 27080 16454 27108 18702
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 18426 27568 18566
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27632 18222 27660 19207
rect 28736 18970 28764 19343
rect 28724 18964 28776 18970
rect 28724 18906 28776 18912
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27344 18080 27396 18086
rect 27344 18022 27396 18028
rect 27356 17882 27384 18022
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 27540 17134 27568 17478
rect 27528 17128 27580 17134
rect 27528 17070 27580 17076
rect 27896 17128 27948 17134
rect 27896 17070 27948 17076
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27252 16108 27304 16114
rect 27252 16050 27304 16056
rect 27264 15434 27292 16050
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 15162 27292 15370
rect 27540 15366 27568 17070
rect 27908 16794 27936 17070
rect 28368 16998 28396 17478
rect 28644 17270 28672 17478
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28356 16992 28408 16998
rect 28356 16934 28408 16940
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 27988 15972 28040 15978
rect 27988 15914 28040 15920
rect 28000 15502 28028 15914
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15638 28212 15846
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27712 15088 27764 15094
rect 27712 15030 27764 15036
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14618 27384 14962
rect 27528 14952 27580 14958
rect 27526 14920 27528 14929
rect 27580 14920 27582 14929
rect 27526 14855 27582 14864
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 27080 14074 27108 14350
rect 27252 14272 27304 14278
rect 27252 14214 27304 14220
rect 27528 14272 27580 14278
rect 27528 14214 27580 14220
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27264 14074 27292 14214
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27540 14006 27568 14214
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27632 13938 27660 14214
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 26976 13796 27028 13802
rect 26976 13738 27028 13744
rect 27264 13530 27292 13874
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27448 12918 27476 13806
rect 27620 13728 27672 13734
rect 27620 13670 27672 13676
rect 27632 13530 27660 13670
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 27724 13326 27752 15030
rect 28276 14890 28304 15370
rect 28368 14890 28396 16934
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28552 15094 28580 15574
rect 29000 15360 29052 15366
rect 29000 15302 29052 15308
rect 28540 15088 28592 15094
rect 28540 15030 28592 15036
rect 29012 15026 29040 15302
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28264 14884 28316 14890
rect 28264 14826 28316 14832
rect 28356 14884 28408 14890
rect 28356 14826 28408 14832
rect 28736 14550 28764 14894
rect 28908 14884 28960 14890
rect 28908 14826 28960 14832
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28828 14618 28856 14758
rect 28816 14612 28868 14618
rect 28816 14554 28868 14560
rect 28724 14544 28776 14550
rect 28724 14486 28776 14492
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27908 13326 27936 13670
rect 28000 13530 28028 14350
rect 28448 13932 28500 13938
rect 28448 13874 28500 13880
rect 27988 13524 28040 13530
rect 27988 13466 28040 13472
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27436 12912 27488 12918
rect 27436 12854 27488 12860
rect 27528 12844 27580 12850
rect 27528 12786 27580 12792
rect 26056 12436 26108 12442
rect 26056 12378 26108 12384
rect 27160 12436 27212 12442
rect 27160 12378 27212 12384
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25320 9920 25372 9926
rect 25320 9862 25372 9868
rect 25332 9382 25360 9862
rect 25424 9654 25452 10406
rect 25412 9648 25464 9654
rect 25412 9590 25464 9596
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25228 9104 25280 9110
rect 25228 9046 25280 9052
rect 25136 8968 25188 8974
rect 23400 8894 23520 8922
rect 25136 8910 25188 8916
rect 23492 8430 23520 8894
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 23572 8560 23624 8566
rect 23572 8502 23624 8508
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23492 7886 23520 8366
rect 23584 8090 23612 8502
rect 24688 8498 24716 8774
rect 25608 8566 25636 12038
rect 26160 11898 26188 12174
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26068 11778 26096 11834
rect 26068 11762 26188 11778
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 26068 11756 26200 11762
rect 26068 11750 26148 11756
rect 25700 11354 25728 11698
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 25884 11354 25912 11630
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 26068 10742 26096 11750
rect 26148 11698 26200 11704
rect 26056 10736 26108 10742
rect 26056 10678 26108 10684
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25884 10130 25912 10406
rect 25872 10124 25924 10130
rect 25872 10066 25924 10072
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25792 9722 25820 9998
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25976 9722 26004 9862
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 26068 9654 26096 10678
rect 26620 10062 26648 11834
rect 26976 11212 27028 11218
rect 26976 11154 27028 11160
rect 26988 10742 27016 11154
rect 26976 10736 27028 10742
rect 26976 10678 27028 10684
rect 27172 10062 27200 12378
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27448 10810 27476 12038
rect 27540 11626 27568 12786
rect 27632 12782 27660 13126
rect 27724 12986 27752 13262
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27816 12782 27844 13262
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27908 12714 27936 13126
rect 28000 12986 28028 13466
rect 28080 13252 28132 13258
rect 28080 13194 28132 13200
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27896 12708 27948 12714
rect 27896 12650 27948 12656
rect 28000 12434 28028 12786
rect 27816 12406 28028 12434
rect 27816 12170 27844 12406
rect 28092 12238 28120 13194
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 27804 12164 27856 12170
rect 27804 12106 27856 12112
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 28184 11150 28212 12786
rect 28264 12776 28316 12782
rect 28264 12718 28316 12724
rect 28276 11558 28304 12718
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 27540 10538 27568 10610
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27896 10464 27948 10470
rect 27896 10406 27948 10412
rect 27356 10062 27384 10406
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 27160 10056 27212 10062
rect 27160 9998 27212 10004
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 26068 9110 26096 9590
rect 26620 9110 26648 9998
rect 27908 9994 27936 10406
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27528 9920 27580 9926
rect 27528 9862 27580 9868
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 26056 9104 26108 9110
rect 26056 9046 26108 9052
rect 26608 9104 26660 9110
rect 26608 9046 26660 9052
rect 26068 8634 26096 9046
rect 27356 9042 27384 9386
rect 27436 9104 27488 9110
rect 27436 9046 27488 9052
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 26700 8832 26752 8838
rect 26700 8774 26752 8780
rect 26712 8634 26740 8774
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 25596 8560 25648 8566
rect 25596 8502 25648 8508
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 25504 8424 25556 8430
rect 25608 8412 25636 8502
rect 27448 8430 27476 9046
rect 27540 8974 27568 9862
rect 28000 9722 28028 10610
rect 28092 10470 28120 11018
rect 28184 10810 28212 11086
rect 28264 11008 28316 11014
rect 28264 10950 28316 10956
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 28092 10266 28120 10406
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 28276 9926 28304 10950
rect 28368 10674 28396 10950
rect 28460 10674 28488 13874
rect 28644 13870 28672 14418
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28736 13326 28764 14282
rect 28920 14278 28948 14826
rect 29104 14618 29132 19654
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 17746 29224 18702
rect 29472 18222 29500 19382
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29460 18216 29512 18222
rect 29460 18158 29512 18164
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29368 17672 29420 17678
rect 29368 17614 29420 17620
rect 29276 17060 29328 17066
rect 29276 17002 29328 17008
rect 29288 16658 29316 17002
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29288 16425 29316 16458
rect 29274 16416 29330 16425
rect 29274 16351 29330 16360
rect 29380 16046 29408 17614
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 29196 15706 29224 15846
rect 29288 15706 29316 15846
rect 29184 15700 29236 15706
rect 29184 15642 29236 15648
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29472 15434 29500 18158
rect 29564 17882 29592 18226
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29552 17740 29604 17746
rect 29552 17682 29604 17688
rect 29564 17202 29592 17682
rect 29552 17196 29604 17202
rect 29552 17138 29604 17144
rect 29460 15428 29512 15434
rect 29460 15370 29512 15376
rect 29092 14612 29144 14618
rect 29092 14554 29144 14560
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 29196 14498 29224 14554
rect 29012 14470 29224 14498
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28724 13320 28776 13326
rect 28724 13262 28776 13268
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 28644 11150 28672 11494
rect 28736 11354 28764 13262
rect 28816 12436 28868 12442
rect 28816 12378 28868 12384
rect 28724 11348 28776 11354
rect 28724 11290 28776 11296
rect 28828 11234 28856 12378
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28920 11354 28948 11494
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 28736 11206 28856 11234
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28736 10674 28764 11206
rect 28816 11008 28868 11014
rect 28816 10950 28868 10956
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28724 10668 28776 10674
rect 28724 10610 28776 10616
rect 28460 10130 28488 10610
rect 28828 10130 28856 10950
rect 28920 10810 28948 10950
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 28920 10266 28948 10610
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28816 10124 28868 10130
rect 28816 10066 28868 10072
rect 28264 9920 28316 9926
rect 28264 9862 28316 9868
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28184 9178 28212 9522
rect 28276 9518 28304 9862
rect 29012 9722 29040 14470
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29288 12986 29316 13874
rect 29472 13308 29500 15370
rect 29564 14006 29592 17138
rect 29656 14958 29684 19722
rect 29748 19514 29776 20198
rect 29932 20058 29960 20402
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 30024 18970 30052 20402
rect 30300 20330 30328 20810
rect 30484 20346 30512 24006
rect 30576 22778 30604 24822
rect 30668 24750 30696 25094
rect 31220 24954 31248 25638
rect 31208 24948 31260 24954
rect 31208 24890 31260 24896
rect 32220 24880 32272 24886
rect 32220 24822 32272 24828
rect 30656 24744 30708 24750
rect 30656 24686 30708 24692
rect 30668 24614 30696 24686
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 31116 24608 31168 24614
rect 31116 24550 31168 24556
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 30668 24070 30696 24550
rect 31128 24274 31156 24550
rect 31116 24268 31168 24274
rect 31116 24210 31168 24216
rect 31680 24138 31708 24550
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30656 23520 30708 23526
rect 30656 23462 30708 23468
rect 30840 23520 30892 23526
rect 30840 23462 30892 23468
rect 30668 23118 30696 23462
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30748 22976 30800 22982
rect 30748 22918 30800 22924
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30760 22710 30788 22918
rect 30852 22778 30880 23462
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30748 22704 30800 22710
rect 30748 22646 30800 22652
rect 31300 22568 31352 22574
rect 31300 22510 31352 22516
rect 30748 22432 30800 22438
rect 30748 22374 30800 22380
rect 30760 22098 30788 22374
rect 31312 22166 31340 22510
rect 31300 22160 31352 22166
rect 31300 22102 31352 22108
rect 30748 22092 30800 22098
rect 30748 22034 30800 22040
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30668 21690 30696 21898
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 31312 20466 31340 22102
rect 31760 22024 31812 22030
rect 31760 21966 31812 21972
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 31772 21690 31800 21966
rect 32140 21690 32168 21966
rect 32232 21894 32260 24822
rect 33140 24744 33192 24750
rect 33140 24686 33192 24692
rect 32588 24200 32640 24206
rect 32588 24142 32640 24148
rect 32600 23866 32628 24142
rect 33152 24070 33180 24686
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 32600 23594 32628 23802
rect 33152 23798 33180 24006
rect 33140 23792 33192 23798
rect 33140 23734 33192 23740
rect 32588 23588 32640 23594
rect 32588 23530 32640 23536
rect 32600 23474 32628 23530
rect 32864 23520 32916 23526
rect 32600 23446 32720 23474
rect 32864 23462 32916 23468
rect 32588 22432 32640 22438
rect 32588 22374 32640 22380
rect 32600 22234 32628 22374
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32692 22094 32720 23446
rect 32876 23186 32904 23462
rect 33152 23254 33180 23734
rect 33140 23248 33192 23254
rect 33140 23190 33192 23196
rect 32864 23180 32916 23186
rect 32864 23122 32916 23128
rect 32876 22760 32904 23122
rect 32956 22772 33008 22778
rect 32876 22732 32956 22760
rect 32876 22438 32904 22732
rect 32956 22714 33008 22720
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32692 22066 32812 22094
rect 32588 22024 32640 22030
rect 32416 21972 32588 21978
rect 32416 21966 32640 21972
rect 32416 21950 32628 21966
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 31484 21344 31536 21350
rect 31484 21286 31536 21292
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31496 20942 31524 21286
rect 31588 21078 31616 21286
rect 31576 21072 31628 21078
rect 31576 21014 31628 21020
rect 31484 20936 31536 20942
rect 31484 20878 31536 20884
rect 31392 20868 31444 20874
rect 31392 20810 31444 20816
rect 31404 20466 31432 20810
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 31300 20460 31352 20466
rect 31300 20402 31352 20408
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 30288 20324 30340 20330
rect 30288 20266 30340 20272
rect 30392 20318 30512 20346
rect 30300 19786 30328 20266
rect 30288 19780 30340 19786
rect 30288 19722 30340 19728
rect 30012 18964 30064 18970
rect 30012 18906 30064 18912
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29840 16794 29868 17138
rect 29920 17128 29972 17134
rect 29920 17070 29972 17076
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29932 16561 29960 17070
rect 29918 16552 29974 16561
rect 30024 16522 30052 18906
rect 30392 18834 30420 20318
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30484 19854 30512 20198
rect 30852 20058 30880 20402
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30840 20052 30892 20058
rect 30840 19994 30892 20000
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30564 19440 30616 19446
rect 30564 19382 30616 19388
rect 30576 18970 30604 19382
rect 30564 18964 30616 18970
rect 30564 18906 30616 18912
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30760 18170 30788 19994
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 31036 19514 31064 19654
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 30840 18624 30892 18630
rect 30840 18566 30892 18572
rect 30852 18358 30880 18566
rect 30840 18352 30892 18358
rect 30840 18294 30892 18300
rect 30760 18142 30880 18170
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30196 17740 30248 17746
rect 30196 17682 30248 17688
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30116 16590 30144 17478
rect 30208 17134 30236 17682
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30196 17128 30248 17134
rect 30196 17070 30248 17076
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 29918 16487 29974 16496
rect 30012 16516 30064 16522
rect 29932 16250 29960 16487
rect 30012 16458 30064 16464
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 30024 16130 30052 16458
rect 29748 16102 30052 16130
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29748 14618 29776 16102
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29932 15366 29960 15982
rect 29920 15360 29972 15366
rect 29920 15302 29972 15308
rect 30104 15360 30156 15366
rect 30104 15302 30156 15308
rect 29932 15026 29960 15302
rect 30116 15162 30144 15302
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30012 15088 30064 15094
rect 30208 15042 30236 17070
rect 30576 16590 30604 17614
rect 30760 17542 30788 18022
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30668 17338 30696 17478
rect 30656 17332 30708 17338
rect 30656 17274 30708 17280
rect 30564 16584 30616 16590
rect 30564 16526 30616 16532
rect 30472 16516 30524 16522
rect 30472 16458 30524 16464
rect 30484 15638 30512 16458
rect 30852 16182 30880 18142
rect 31312 17678 31340 20402
rect 31404 19854 31432 20402
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31312 16998 31340 17614
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 31036 16794 31064 16934
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31588 16658 31616 21014
rect 31956 20602 31984 21490
rect 32416 21486 32444 21950
rect 32404 21480 32456 21486
rect 32404 21422 32456 21428
rect 31944 20596 31996 20602
rect 31944 20538 31996 20544
rect 32036 19848 32088 19854
rect 32036 19790 32088 19796
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32048 19514 32076 19790
rect 32036 19508 32088 19514
rect 32036 19450 32088 19456
rect 32232 19446 32260 19790
rect 32416 19786 32444 21422
rect 32784 19922 32812 22066
rect 32864 22024 32916 22030
rect 32864 21966 32916 21972
rect 32876 21690 32904 21966
rect 32864 21684 32916 21690
rect 32864 21626 32916 21632
rect 32968 20330 32996 22510
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 33060 21554 33088 21830
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 33152 21146 33180 21830
rect 33140 21140 33192 21146
rect 33140 21082 33192 21088
rect 33048 20800 33100 20806
rect 33048 20742 33100 20748
rect 32956 20324 33008 20330
rect 32956 20266 33008 20272
rect 32772 19916 32824 19922
rect 32772 19858 32824 19864
rect 32404 19780 32456 19786
rect 32404 19722 32456 19728
rect 32588 19780 32640 19786
rect 32588 19722 32640 19728
rect 32600 19514 32628 19722
rect 32588 19508 32640 19514
rect 32588 19450 32640 19456
rect 32220 19440 32272 19446
rect 32220 19382 32272 19388
rect 32784 19334 32812 19858
rect 32968 19700 32996 20266
rect 33060 19854 33088 20742
rect 33140 20460 33192 20466
rect 33140 20402 33192 20408
rect 33152 20058 33180 20402
rect 33140 20052 33192 20058
rect 33140 19994 33192 20000
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 32968 19672 33088 19700
rect 32692 19306 32812 19334
rect 32956 19372 33008 19378
rect 32956 19314 33008 19320
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32312 18080 32364 18086
rect 32312 18022 32364 18028
rect 32220 17536 32272 17542
rect 32220 17478 32272 17484
rect 32232 17338 32260 17478
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31680 16794 31708 17070
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 31024 16652 31076 16658
rect 31024 16594 31076 16600
rect 31576 16652 31628 16658
rect 31576 16594 31628 16600
rect 31036 16538 31064 16594
rect 31036 16510 31156 16538
rect 31128 16454 31156 16510
rect 32128 16516 32180 16522
rect 32128 16458 32180 16464
rect 31024 16448 31076 16454
rect 31024 16390 31076 16396
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31392 16448 31444 16454
rect 31392 16390 31444 16396
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30656 16108 30708 16114
rect 30656 16050 30708 16056
rect 30472 15632 30524 15638
rect 30472 15574 30524 15580
rect 30668 15502 30696 16050
rect 31036 15638 31064 16390
rect 31116 16108 31168 16114
rect 31116 16050 31168 16056
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31024 15632 31076 15638
rect 31024 15574 31076 15580
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30064 15036 30236 15042
rect 30012 15030 30236 15036
rect 29920 15020 29972 15026
rect 30024 15014 30236 15030
rect 29920 14962 29972 14968
rect 29736 14612 29788 14618
rect 29736 14554 29788 14560
rect 29748 14006 29776 14554
rect 29552 14000 29604 14006
rect 29552 13942 29604 13948
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 29552 13320 29604 13326
rect 29472 13280 29552 13308
rect 29552 13262 29604 13268
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29460 12776 29512 12782
rect 29460 12718 29512 12724
rect 29472 12306 29500 12718
rect 29460 12300 29512 12306
rect 29460 12242 29512 12248
rect 29092 10464 29144 10470
rect 29092 10406 29144 10412
rect 29184 10464 29236 10470
rect 29184 10406 29236 10412
rect 29104 9722 29132 10406
rect 29196 10062 29224 10406
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 28172 9172 28224 9178
rect 28172 9114 28224 9120
rect 28276 8974 28304 9454
rect 28632 9104 28684 9110
rect 28632 9046 28684 9052
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 28264 8968 28316 8974
rect 28264 8910 28316 8916
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27632 8498 27660 8774
rect 28000 8634 28028 8774
rect 28644 8634 28672 9046
rect 29564 8974 29592 13262
rect 29828 13252 29880 13258
rect 29828 13194 29880 13200
rect 29840 12986 29868 13194
rect 30104 13184 30156 13190
rect 30104 13126 30156 13132
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 30116 12918 30144 13126
rect 30104 12912 30156 12918
rect 30104 12854 30156 12860
rect 30208 12782 30236 15014
rect 30668 14958 30696 15438
rect 30656 14952 30708 14958
rect 30656 14894 30708 14900
rect 31128 14618 31156 16050
rect 31312 15910 31340 16050
rect 31404 16046 31432 16390
rect 32140 16250 32168 16458
rect 32128 16244 32180 16250
rect 32128 16186 32180 16192
rect 32324 16046 32352 18022
rect 32508 17882 32536 18226
rect 32692 18086 32720 19306
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32968 17882 32996 19314
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 32508 17746 32536 17818
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32404 17604 32456 17610
rect 32404 17546 32456 17552
rect 32864 17604 32916 17610
rect 32864 17546 32916 17552
rect 32416 17270 32444 17546
rect 32876 17354 32904 17546
rect 32600 17326 32904 17354
rect 32600 17270 32628 17326
rect 32404 17264 32456 17270
rect 32404 17206 32456 17212
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32772 17264 32824 17270
rect 32772 17206 32824 17212
rect 32404 17060 32456 17066
rect 32784 17048 32812 17206
rect 32456 17020 32812 17048
rect 32404 17002 32456 17008
rect 32876 16998 32904 17326
rect 32864 16992 32916 16998
rect 32864 16934 32916 16940
rect 32968 16794 32996 17818
rect 33060 17626 33088 19672
rect 33336 19310 33364 25774
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35440 25424 35492 25430
rect 35440 25366 35492 25372
rect 35452 25265 35480 25366
rect 35438 25256 35494 25265
rect 35438 25191 35494 25200
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35346 24576 35402 24585
rect 34934 24508 35242 24517
rect 35346 24511 35402 24520
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35360 24410 35388 24511
rect 33600 24404 33652 24410
rect 33600 24346 33652 24352
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 33612 23730 33640 24346
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33704 23254 33732 23666
rect 33876 23520 33928 23526
rect 33796 23480 33876 23508
rect 33692 23248 33744 23254
rect 33692 23190 33744 23196
rect 33796 22760 33824 23480
rect 33876 23462 33928 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 35452 23225 35480 23258
rect 35438 23216 35494 23225
rect 35438 23151 35494 23160
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 33612 22732 33824 22760
rect 33612 22234 33640 22732
rect 33692 22636 33744 22642
rect 33692 22578 33744 22584
rect 33600 22228 33652 22234
rect 33600 22170 33652 22176
rect 33704 22030 33732 22578
rect 33692 22024 33744 22030
rect 33692 21966 33744 21972
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 33520 21690 33548 21830
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 33704 20466 33732 21966
rect 33796 21894 33824 22732
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 33784 21888 33836 21894
rect 33784 21830 33836 21836
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 34336 20460 34388 20466
rect 34336 20402 34388 20408
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 33428 19514 33456 19858
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33796 19514 33824 19654
rect 34348 19514 34376 20402
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35530 19816 35586 19825
rect 35530 19751 35532 19760
rect 35584 19751 35586 19760
rect 35532 19722 35584 19728
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33784 19508 33836 19514
rect 33784 19450 33836 19456
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 33324 19304 33376 19310
rect 33324 19246 33376 19252
rect 33336 18222 33364 19246
rect 35438 19136 35494 19145
rect 34934 19068 35242 19077
rect 35438 19071 35494 19080
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35452 18902 35480 19071
rect 35440 18896 35492 18902
rect 35440 18838 35492 18844
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35346 18320 35402 18329
rect 35346 18255 35348 18264
rect 35400 18255 35402 18264
rect 35348 18226 35400 18232
rect 33324 18216 33376 18222
rect 33324 18158 33376 18164
rect 34336 18080 34388 18086
rect 34336 18022 34388 18028
rect 34348 17882 34376 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 34336 17876 34388 17882
rect 34336 17818 34388 17824
rect 33520 17678 33548 17818
rect 34060 17808 34112 17814
rect 34058 17776 34060 17785
rect 34112 17776 34114 17785
rect 34058 17711 34114 17720
rect 33508 17672 33560 17678
rect 33060 17598 33180 17626
rect 33508 17614 33560 17620
rect 33048 17536 33100 17542
rect 33048 17478 33100 17484
rect 33060 17338 33088 17478
rect 33048 17332 33100 17338
rect 33048 17274 33100 17280
rect 33152 17218 33180 17598
rect 33692 17536 33744 17542
rect 33692 17478 33744 17484
rect 33060 17190 33180 17218
rect 33232 17196 33284 17202
rect 33060 16998 33088 17190
rect 33232 17138 33284 17144
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 32956 16788 33008 16794
rect 32956 16730 33008 16736
rect 33244 16726 33272 17138
rect 33232 16720 33284 16726
rect 33232 16662 33284 16668
rect 32954 16552 33010 16561
rect 32954 16487 32956 16496
rect 33008 16487 33010 16496
rect 32956 16458 33008 16464
rect 32404 16448 32456 16454
rect 32404 16390 32456 16396
rect 32416 16114 32444 16390
rect 32968 16250 32996 16458
rect 33244 16250 33272 16662
rect 33704 16590 33732 17478
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 38844 17128 38896 17134
rect 38842 17096 38844 17105
rect 38896 17096 38898 17105
rect 38842 17031 38898 17040
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 33704 16454 33732 16526
rect 33508 16448 33560 16454
rect 33508 16390 33560 16396
rect 33692 16448 33744 16454
rect 33692 16390 33744 16396
rect 32956 16244 33008 16250
rect 32956 16186 33008 16192
rect 33232 16244 33284 16250
rect 33232 16186 33284 16192
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 32312 16040 32364 16046
rect 32312 15982 32364 15988
rect 31300 15904 31352 15910
rect 31300 15846 31352 15852
rect 31496 15366 31524 15982
rect 32324 15638 32352 15982
rect 33520 15910 33548 16390
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 33508 15904 33560 15910
rect 33508 15846 33560 15852
rect 33784 15904 33836 15910
rect 33784 15846 33836 15852
rect 33796 15638 33824 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 37292 15745 37320 16050
rect 37278 15736 37334 15745
rect 35440 15700 35492 15706
rect 37278 15671 37334 15680
rect 35440 15642 35492 15648
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 33784 15632 33836 15638
rect 33784 15574 33836 15580
rect 31576 15428 31628 15434
rect 31576 15370 31628 15376
rect 31484 15360 31536 15366
rect 31484 15302 31536 15308
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30392 13258 30420 14214
rect 30564 13932 30616 13938
rect 30564 13874 30616 13880
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30380 13252 30432 13258
rect 30380 13194 30432 13200
rect 30484 12986 30512 13670
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 30576 12782 30604 13874
rect 30852 13530 30880 14350
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 31404 13938 31432 14214
rect 31496 14074 31524 15302
rect 31588 14618 31616 15370
rect 31576 14612 31628 14618
rect 31576 14554 31628 14560
rect 32128 14544 32180 14550
rect 32128 14486 32180 14492
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 31576 14340 31628 14346
rect 31576 14282 31628 14288
rect 31588 14074 31616 14282
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 31392 13932 31444 13938
rect 31392 13874 31444 13880
rect 31220 13530 31248 13874
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 31208 13524 31260 13530
rect 31208 13466 31260 13472
rect 30852 12850 30880 13466
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 31404 12442 31432 13874
rect 31864 13530 31892 14350
rect 32048 14074 32076 14350
rect 32036 14068 32088 14074
rect 32036 14010 32088 14016
rect 32036 13932 32088 13938
rect 32140 13920 32168 14486
rect 32088 13892 32168 13920
rect 32220 13932 32272 13938
rect 32036 13874 32088 13880
rect 32220 13874 32272 13880
rect 31852 13524 31904 13530
rect 31852 13466 31904 13472
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 31392 12436 31444 12442
rect 31392 12378 31444 12384
rect 31772 12374 31800 13126
rect 31956 12918 31984 13262
rect 32048 12918 32076 13874
rect 32232 13394 32260 13874
rect 32220 13388 32272 13394
rect 32220 13330 32272 13336
rect 31944 12912 31996 12918
rect 31944 12854 31996 12860
rect 32036 12912 32088 12918
rect 32036 12854 32088 12860
rect 31852 12640 31904 12646
rect 31852 12582 31904 12588
rect 31760 12368 31812 12374
rect 31760 12310 31812 12316
rect 31864 12306 31892 12582
rect 31852 12300 31904 12306
rect 31852 12242 31904 12248
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31220 11676 31248 12038
rect 31680 11898 31708 12038
rect 31668 11892 31720 11898
rect 31668 11834 31720 11840
rect 31864 11762 31892 12242
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 31392 11688 31444 11694
rect 31220 11648 31392 11676
rect 31392 11630 31444 11636
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30484 11150 30512 11494
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30932 11008 30984 11014
rect 30932 10950 30984 10956
rect 30944 10742 30972 10950
rect 31404 10810 31432 11630
rect 31956 11626 31984 12854
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32140 12442 32168 12786
rect 32128 12436 32180 12442
rect 32128 12378 32180 12384
rect 32220 12232 32272 12238
rect 32324 12220 32352 15574
rect 35452 15065 35480 15642
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35438 15056 35494 15065
rect 35438 14991 35494 15000
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 32496 14476 32548 14482
rect 32496 14418 32548 14424
rect 32508 13938 32536 14418
rect 35624 14408 35676 14414
rect 35622 14376 35624 14385
rect 35676 14376 35678 14385
rect 35622 14311 35678 14320
rect 33048 14272 33100 14278
rect 33048 14214 33100 14220
rect 33060 14074 33088 14214
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 33048 14068 33100 14074
rect 33048 14010 33100 14016
rect 32496 13932 32548 13938
rect 32496 13874 32548 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32272 12192 32352 12220
rect 32220 12174 32272 12180
rect 32128 12164 32180 12170
rect 32128 12106 32180 12112
rect 32140 11830 32168 12106
rect 32128 11824 32180 11830
rect 32128 11766 32180 11772
rect 31944 11620 31996 11626
rect 31944 11562 31996 11568
rect 32232 11354 32260 12174
rect 32600 11898 32628 12786
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34518 12336 34574 12345
rect 34518 12271 34574 12280
rect 34532 12238 34560 12271
rect 34152 12232 34204 12238
rect 34152 12174 34204 12180
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 32588 11892 32640 11898
rect 32588 11834 32640 11840
rect 32220 11348 32272 11354
rect 32220 11290 32272 11296
rect 32128 11076 32180 11082
rect 32128 11018 32180 11024
rect 32140 10810 32168 11018
rect 31392 10804 31444 10810
rect 31392 10746 31444 10752
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 30932 10736 30984 10742
rect 30932 10678 30984 10684
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29656 10130 29684 10406
rect 29748 10198 29776 10610
rect 29828 10600 29880 10606
rect 29828 10542 29880 10548
rect 30380 10600 30432 10606
rect 30380 10542 30432 10548
rect 29736 10192 29788 10198
rect 29736 10134 29788 10140
rect 29644 10124 29696 10130
rect 29644 10066 29696 10072
rect 29644 9376 29696 9382
rect 29644 9318 29696 9324
rect 29656 9178 29684 9318
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28920 8498 28948 8842
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 25556 8384 25636 8412
rect 27436 8424 27488 8430
rect 25504 8366 25556 8372
rect 27436 8366 27488 8372
rect 25136 8356 25188 8362
rect 25136 8298 25188 8304
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23492 7546 23520 7822
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23216 2746 23336 2774
rect 23216 800 23244 2746
rect 25148 800 25176 8298
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26620 7954 26648 8230
rect 28000 7954 28028 8298
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 28920 7886 28948 8434
rect 29012 8090 29040 8910
rect 29840 8838 29868 10542
rect 30392 10266 30420 10542
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30380 10260 30432 10266
rect 30380 10202 30432 10208
rect 30852 10130 30880 10406
rect 30944 10266 30972 10678
rect 31300 10668 31352 10674
rect 31300 10610 31352 10616
rect 32864 10668 32916 10674
rect 32864 10610 32916 10616
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30392 9722 30420 9998
rect 30380 9716 30432 9722
rect 30852 9674 30880 10066
rect 31312 9994 31340 10610
rect 32876 10266 32904 10610
rect 34164 10606 34192 12174
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 38200 11348 38252 11354
rect 38200 11290 38252 11296
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 34152 10600 34204 10606
rect 34152 10542 34204 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10305 35388 10610
rect 35346 10296 35402 10305
rect 32864 10260 32916 10266
rect 35346 10231 35402 10240
rect 32864 10202 32916 10208
rect 31300 9988 31352 9994
rect 31300 9930 31352 9936
rect 31312 9722 31340 9930
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 30380 9658 30432 9664
rect 30484 9646 30880 9674
rect 31300 9716 31352 9722
rect 31300 9658 31352 9664
rect 30104 8900 30156 8906
rect 30104 8842 30156 8848
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 30116 8634 30144 8842
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30484 8566 30512 9646
rect 31312 9178 31340 9658
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 31300 9172 31352 9178
rect 31300 9114 31352 9120
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 30472 8560 30524 8566
rect 30472 8502 30524 8508
rect 38212 8498 38240 11290
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 27252 7812 27304 7818
rect 27252 7754 27304 7760
rect 27264 7546 27292 7754
rect 29196 7750 29224 8434
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 29012 800 29040 7686
rect 29748 7410 29776 8434
rect 38384 8356 38436 8362
rect 38384 8298 38436 8304
rect 38396 8265 38424 8298
rect 38382 8256 38438 8265
rect 34934 8188 35242 8197
rect 38382 8191 38438 8200
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 10966 0 11022 800
rect 14186 0 14242 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 23202 0 23258 800
rect 25134 0 25190 800
rect 28998 0 29054 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 3422 29960 3478 30016
rect 938 25200 994 25256
rect 1122 24556 1124 24576
rect 1124 24556 1176 24576
rect 1176 24556 1178 24576
rect 1122 24520 1178 24556
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 3974 22480 4030 22536
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4066 20440 4122 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19760 4122 19816
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4066 18400 4122 18456
rect 13726 27124 13782 27160
rect 13726 27104 13728 27124
rect 13728 27104 13780 27124
rect 13780 27104 13782 27124
rect 12530 20324 12586 20360
rect 12530 20304 12532 20324
rect 12532 20304 12584 20324
rect 12584 20304 12586 20324
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 2778 15680 2834 15736
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 12990 19388 12992 19408
rect 12992 19388 13044 19408
rect 13044 19388 13046 19408
rect 12990 19352 13046 19388
rect 17038 27240 17094 27296
rect 16946 27104 17002 27160
rect 17038 26968 17094 27024
rect 16946 26852 17002 26888
rect 16946 26832 16948 26852
rect 16948 26832 17000 26852
rect 17000 26832 17002 26852
rect 9402 16516 9458 16552
rect 9402 16496 9404 16516
rect 9404 16496 9456 16516
rect 9456 16496 9458 16516
rect 4066 13640 4122 13696
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4066 11620 4122 11656
rect 4066 11600 4068 11620
rect 4068 11600 4120 11620
rect 4120 11600 4122 11620
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 17682 27240 17738 27296
rect 19062 26968 19118 27024
rect 18786 26832 18842 26888
rect 16578 21972 16580 21992
rect 16580 21972 16632 21992
rect 16632 21972 16634 21992
rect 16578 21936 16634 21972
rect 16670 19388 16672 19408
rect 16672 19388 16724 19408
rect 16724 19388 16726 19408
rect 16670 19352 16726 19388
rect 18694 20712 18750 20768
rect 17498 20340 17500 20360
rect 17500 20340 17552 20360
rect 17552 20340 17554 20360
rect 17498 20304 17554 20340
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 25226 23160 25282 23216
rect 23570 19352 23626 19408
rect 22466 19216 22522 19272
rect 19982 12144 20038 12200
rect 23662 16496 23718 16552
rect 23294 14864 23350 14920
rect 22926 12144 22982 12200
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35438 25880 35494 25936
rect 24674 16532 24676 16552
rect 24676 16532 24728 16552
rect 24728 16532 24730 16552
rect 24674 16496 24730 16532
rect 28722 19352 28778 19408
rect 27618 19216 27674 19272
rect 23754 12180 23756 12200
rect 23756 12180 23808 12200
rect 23808 12180 23810 12200
rect 23754 12144 23810 12180
rect 27526 14900 27528 14920
rect 27528 14900 27580 14920
rect 27580 14900 27582 14920
rect 27526 14864 27582 14900
rect 29274 16360 29330 16416
rect 29918 16496 29974 16552
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35438 25200 35494 25256
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35346 24520 35402 24576
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35438 23160 35494 23216
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35530 19780 35586 19816
rect 35530 19760 35532 19780
rect 35532 19760 35584 19780
rect 35584 19760 35586 19780
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35438 19080 35494 19136
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 35346 18284 35402 18320
rect 35346 18264 35348 18284
rect 35348 18264 35400 18284
rect 35400 18264 35402 18284
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34058 17756 34060 17776
rect 34060 17756 34112 17776
rect 34112 17756 34114 17776
rect 34058 17720 34114 17756
rect 32954 16516 33010 16552
rect 32954 16496 32956 16516
rect 32956 16496 33008 16516
rect 33008 16496 33010 16516
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 38842 17076 38844 17096
rect 38844 17076 38896 17096
rect 38896 17076 38898 17096
rect 38842 17040 38898 17076
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 37278 15680 37334 15736
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35438 15000 35494 15056
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 35622 14356 35624 14376
rect 35624 14356 35676 14376
rect 35676 14356 35678 14376
rect 35622 14320 35678 14356
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34518 12280 34574 12336
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35346 10240 35402 10296
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 38382 8200 38438 8256
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 0 30018 800 30048
rect 3417 30018 3483 30021
rect 0 30016 3483 30018
rect 0 29960 3422 30016
rect 3478 29960 3483 30016
rect 0 29958 3483 29960
rect 0 29928 800 29958
rect 3417 29955 3483 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 17033 27298 17099 27301
rect 17677 27298 17743 27301
rect 17033 27296 17743 27298
rect 17033 27240 17038 27296
rect 17094 27240 17682 27296
rect 17738 27240 17743 27296
rect 17033 27238 17743 27240
rect 17033 27235 17099 27238
rect 17677 27235 17743 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 13721 27162 13787 27165
rect 16941 27162 17007 27165
rect 13721 27160 17007 27162
rect 13721 27104 13726 27160
rect 13782 27104 16946 27160
rect 17002 27104 17007 27160
rect 13721 27102 17007 27104
rect 13721 27099 13787 27102
rect 16941 27099 17007 27102
rect 17033 27026 17099 27029
rect 19057 27026 19123 27029
rect 17033 27024 19123 27026
rect 17033 26968 17038 27024
rect 17094 26968 19062 27024
rect 19118 26968 19123 27024
rect 17033 26966 19123 26968
rect 17033 26963 17099 26966
rect 19057 26963 19123 26966
rect 16941 26890 17007 26893
rect 18781 26890 18847 26893
rect 16941 26888 18847 26890
rect 16941 26832 16946 26888
rect 17002 26832 18786 26888
rect 18842 26832 18847 26888
rect 16941 26830 18847 26832
rect 16941 26827 17007 26830
rect 18781 26827 18847 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 35433 25938 35499 25941
rect 39200 25938 40000 25968
rect 35433 25936 40000 25938
rect 35433 25880 35438 25936
rect 35494 25880 40000 25936
rect 35433 25878 40000 25880
rect 35433 25875 35499 25878
rect 39200 25848 40000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 35433 25258 35499 25261
rect 39200 25258 40000 25288
rect 35433 25256 40000 25258
rect 35433 25200 35438 25256
rect 35494 25200 40000 25256
rect 35433 25198 40000 25200
rect 35433 25195 35499 25198
rect 39200 25168 40000 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 0 24578 800 24608
rect 1117 24578 1183 24581
rect 0 24576 1183 24578
rect 0 24520 1122 24576
rect 1178 24520 1183 24576
rect 0 24518 1183 24520
rect 0 24488 800 24518
rect 1117 24515 1183 24518
rect 35341 24578 35407 24581
rect 39200 24578 40000 24608
rect 35341 24576 40000 24578
rect 35341 24520 35346 24576
rect 35402 24520 40000 24576
rect 35341 24518 40000 24520
rect 35341 24515 35407 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 40000 24518
rect 34930 24447 35246 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 25078 23156 25084 23220
rect 25148 23218 25154 23220
rect 25221 23218 25287 23221
rect 25148 23216 25287 23218
rect 25148 23160 25226 23216
rect 25282 23160 25287 23216
rect 25148 23158 25287 23160
rect 25148 23156 25154 23158
rect 25221 23155 25287 23158
rect 35433 23218 35499 23221
rect 39200 23218 40000 23248
rect 35433 23216 40000 23218
rect 35433 23160 35438 23216
rect 35494 23160 40000 23216
rect 35433 23158 40000 23160
rect 35433 23155 35499 23158
rect 39200 23128 40000 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 0 22538 800 22568
rect 3969 22538 4035 22541
rect 0 22536 4035 22538
rect 0 22480 3974 22536
rect 4030 22480 4035 22536
rect 0 22478 4035 22480
rect 0 22448 800 22478
rect 3969 22475 4035 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 16573 21994 16639 21997
rect 2730 21992 16639 21994
rect 2730 21936 16578 21992
rect 16634 21936 16639 21992
rect 2730 21934 16639 21936
rect 0 21858 800 21888
rect 2730 21858 2790 21934
rect 16573 21931 16639 21934
rect 0 21798 2790 21858
rect 0 21768 800 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 18689 20772 18755 20773
rect 18638 20708 18644 20772
rect 18708 20770 18755 20772
rect 18708 20768 18800 20770
rect 18750 20712 18800 20768
rect 18708 20710 18800 20712
rect 18708 20708 18755 20710
rect 18689 20707 18755 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 0 20498 800 20528
rect 4061 20498 4127 20501
rect 0 20496 4127 20498
rect 0 20440 4066 20496
rect 4122 20440 4127 20496
rect 0 20438 4127 20440
rect 0 20408 800 20438
rect 4061 20435 4127 20438
rect 12525 20362 12591 20365
rect 17493 20362 17559 20365
rect 12525 20360 17559 20362
rect 12525 20304 12530 20360
rect 12586 20304 17498 20360
rect 17554 20304 17559 20360
rect 12525 20302 17559 20304
rect 12525 20299 12591 20302
rect 17493 20299 17559 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 4061 19818 4127 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 800 19758
rect 4061 19755 4127 19758
rect 35525 19818 35591 19821
rect 39200 19818 40000 19848
rect 35525 19816 40000 19818
rect 35525 19760 35530 19816
rect 35586 19760 40000 19816
rect 35525 19758 40000 19760
rect 35525 19755 35591 19758
rect 39200 19728 40000 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 12985 19410 13051 19413
rect 16665 19410 16731 19413
rect 12985 19408 16731 19410
rect 12985 19352 12990 19408
rect 13046 19352 16670 19408
rect 16726 19352 16731 19408
rect 12985 19350 16731 19352
rect 12985 19347 13051 19350
rect 16665 19347 16731 19350
rect 23565 19410 23631 19413
rect 28717 19410 28783 19413
rect 23565 19408 28783 19410
rect 23565 19352 23570 19408
rect 23626 19352 28722 19408
rect 28778 19352 28783 19408
rect 23565 19350 28783 19352
rect 23565 19347 23631 19350
rect 28717 19347 28783 19350
rect 22461 19274 22527 19277
rect 27613 19274 27679 19277
rect 22461 19272 27679 19274
rect 22461 19216 22466 19272
rect 22522 19216 27618 19272
rect 27674 19216 27679 19272
rect 22461 19214 27679 19216
rect 22461 19211 22527 19214
rect 27613 19211 27679 19214
rect 35433 19138 35499 19141
rect 39200 19138 40000 19168
rect 35433 19136 40000 19138
rect 35433 19080 35438 19136
rect 35494 19080 40000 19136
rect 35433 19078 40000 19080
rect 35433 19075 35499 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 40000 19078
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4061 18458 4127 18461
rect 39200 18458 40000 18488
rect 0 18456 4127 18458
rect 0 18400 4066 18456
rect 4122 18400 4127 18456
rect 0 18398 4127 18400
rect 0 18368 800 18398
rect 4061 18395 4127 18398
rect 36126 18398 40000 18458
rect 35341 18322 35407 18325
rect 36126 18322 36186 18398
rect 39200 18368 40000 18398
rect 35341 18320 36186 18322
rect 35341 18264 35346 18320
rect 35402 18264 36186 18320
rect 35341 18262 36186 18264
rect 35341 18259 35407 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 34053 17778 34119 17781
rect 39200 17778 40000 17808
rect 34053 17776 40000 17778
rect 34053 17720 34058 17776
rect 34114 17720 40000 17776
rect 34053 17718 40000 17720
rect 34053 17715 34119 17718
rect 39200 17688 40000 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 38837 17098 38903 17101
rect 39200 17098 40000 17128
rect 38837 17096 40000 17098
rect 38837 17040 38842 17096
rect 38898 17040 40000 17096
rect 38837 17038 40000 17040
rect 38837 17035 38903 17038
rect 39200 17008 40000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 9397 16554 9463 16557
rect 18638 16554 18644 16556
rect 9397 16552 18644 16554
rect 9397 16496 9402 16552
rect 9458 16496 18644 16552
rect 9397 16494 18644 16496
rect 9397 16491 9463 16494
rect 18638 16492 18644 16494
rect 18708 16554 18714 16556
rect 23657 16554 23723 16557
rect 18708 16552 23723 16554
rect 18708 16496 23662 16552
rect 23718 16496 23723 16552
rect 18708 16494 23723 16496
rect 18708 16492 18714 16494
rect 23657 16491 23723 16494
rect 24669 16554 24735 16557
rect 25078 16554 25084 16556
rect 24669 16552 25084 16554
rect 24669 16496 24674 16552
rect 24730 16496 25084 16552
rect 24669 16494 25084 16496
rect 24669 16491 24735 16494
rect 25078 16492 25084 16494
rect 25148 16492 25154 16556
rect 29913 16554 29979 16557
rect 32949 16554 33015 16557
rect 29913 16552 33015 16554
rect 29913 16496 29918 16552
rect 29974 16496 32954 16552
rect 33010 16496 33015 16552
rect 29913 16494 33015 16496
rect 29913 16491 29979 16494
rect 32949 16491 33015 16494
rect 33182 16494 36186 16554
rect 29269 16418 29335 16421
rect 33182 16418 33242 16494
rect 29269 16416 33242 16418
rect 29269 16360 29274 16416
rect 29330 16360 33242 16416
rect 29269 16358 33242 16360
rect 36126 16418 36186 16494
rect 39200 16418 40000 16448
rect 36126 16358 40000 16418
rect 29269 16355 29335 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 39200 16328 40000 16358
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 2773 15738 2839 15741
rect 0 15736 2839 15738
rect 0 15680 2778 15736
rect 2834 15680 2839 15736
rect 0 15678 2839 15680
rect 0 15648 800 15678
rect 2773 15675 2839 15678
rect 37273 15738 37339 15741
rect 39200 15738 40000 15768
rect 37273 15736 40000 15738
rect 37273 15680 37278 15736
rect 37334 15680 40000 15736
rect 37273 15678 40000 15680
rect 37273 15675 37339 15678
rect 39200 15648 40000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 35433 15058 35499 15061
rect 39200 15058 40000 15088
rect 35433 15056 40000 15058
rect 35433 15000 35438 15056
rect 35494 15000 40000 15056
rect 35433 14998 40000 15000
rect 35433 14995 35499 14998
rect 39200 14968 40000 14998
rect 23289 14922 23355 14925
rect 27521 14922 27587 14925
rect 23289 14920 27587 14922
rect 23289 14864 23294 14920
rect 23350 14864 27526 14920
rect 27582 14864 27587 14920
rect 23289 14862 27587 14864
rect 23289 14859 23355 14862
rect 27521 14859 27587 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 35617 14378 35683 14381
rect 39200 14378 40000 14408
rect 35617 14376 40000 14378
rect 35617 14320 35622 14376
rect 35678 14320 40000 14376
rect 35617 14318 40000 14320
rect 35617 14315 35683 14318
rect 39200 14288 40000 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 0 13698 800 13728
rect 4061 13698 4127 13701
rect 0 13696 4127 13698
rect 0 13640 4066 13696
rect 4122 13640 4127 13696
rect 0 13638 4127 13640
rect 0 13608 800 13638
rect 4061 13635 4127 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 34513 12338 34579 12341
rect 39200 12338 40000 12368
rect 34513 12336 40000 12338
rect 34513 12280 34518 12336
rect 34574 12280 40000 12336
rect 34513 12278 40000 12280
rect 34513 12275 34579 12278
rect 39200 12248 40000 12278
rect 19977 12202 20043 12205
rect 22921 12202 22987 12205
rect 23749 12202 23815 12205
rect 19977 12200 23815 12202
rect 19977 12144 19982 12200
rect 20038 12144 22926 12200
rect 22982 12144 23754 12200
rect 23810 12144 23815 12200
rect 19977 12142 23815 12144
rect 19977 12139 20043 12142
rect 22921 12139 22987 12142
rect 23749 12139 23815 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 0 11658 800 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 800 11598
rect 4061 11595 4127 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 35341 10298 35407 10301
rect 39200 10298 40000 10328
rect 35341 10296 40000 10298
rect 35341 10240 35346 10296
rect 35402 10240 40000 10296
rect 35341 10238 40000 10240
rect 35341 10235 35407 10238
rect 39200 10208 40000 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 38377 8258 38443 8261
rect 39200 8258 40000 8288
rect 38377 8256 40000 8258
rect 38377 8200 38382 8256
rect 38438 8200 40000 8256
rect 38377 8198 40000 8200
rect 38377 8195 38443 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 40000 8198
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 25084 23156 25148 23220
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 18644 20768 18708 20772
rect 18644 20712 18694 20768
rect 18694 20712 18708 20768
rect 18644 20708 18708 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 18644 16492 18708 16556
rect 25084 16492 25148 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 25083 23220 25149 23221
rect 25083 23156 25084 23220
rect 25148 23156 25149 23220
rect 25083 23155 25149 23156
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 18643 20772 18709 20773
rect 18643 20708 18644 20772
rect 18708 20708 18709 20772
rect 18643 20707 18709 20708
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 18646 16557 18706 20707
rect 25086 16557 25146 23155
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 18643 16556 18709 16557
rect 18643 16492 18644 16556
rect 18708 16492 18709 16556
rect 18643 16491 18709 16492
rect 25083 16556 25149 16557
rect 25083 16492 25084 16556
rect 25148 16492 25149 16556
rect 25083 16491 25149 16492
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 38872 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 38872 36920
rect 1056 36642 38872 36684
rect 1056 36260 38872 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 38872 36260
rect 1056 35982 38872 36024
rect 1056 6284 38872 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 38872 6284
rect 1056 6006 38872 6048
rect 1056 5624 38872 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 38872 5624
rect 1056 5346 38872 5388
use sky130_fd_sc_hd__and3b_1  _0676_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 22264 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0677_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20056 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0678_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 21436 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0679_
timestamp 1694700623
transform -1 0 20792 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 23000 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0681_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 22540 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0682_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20516 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0683_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19872 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0684_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15272 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0685_
timestamp 1694700623
transform 1 0 14720 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0686_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 17480 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0687_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0688_
timestamp 1694700623
transform 1 0 18308 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0689_
timestamp 1694700623
transform 1 0 16928 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0690_
timestamp 1694700623
transform -1 0 18216 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0691_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 17664 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0692_
timestamp 1694700623
transform -1 0 16560 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1694700623
transform 1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0694_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0695_
timestamp 1694700623
transform 1 0 12144 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0696_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0697_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1694700623
transform -1 0 13064 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0699_
timestamp 1694700623
transform -1 0 12052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0700_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 20424 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0701_
timestamp 1694700623
transform -1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0702_
timestamp 1694700623
transform -1 0 20056 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0703_
timestamp 1694700623
transform -1 0 13984 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0704_
timestamp 1694700623
transform 1 0 14076 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0705_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16652 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 16192 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0707_
timestamp 1694700623
transform -1 0 16560 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15088 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0710_
timestamp 1694700623
transform -1 0 19872 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0711_
timestamp 1694700623
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13708 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12328 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0715_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13432 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0716_
timestamp 1694700623
transform 1 0 11592 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0717_
timestamp 1694700623
transform 1 0 12328 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0718_
timestamp 1694700623
transform 1 0 13248 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0719_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13432 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14260 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0721_
timestamp 1694700623
transform -1 0 13524 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0722_
timestamp 1694700623
transform 1 0 15548 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1694700623
transform 1 0 15180 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1694700623
transform -1 0 16192 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0725_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14536 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 1694700623
transform -1 0 15640 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0727_
timestamp 1694700623
transform 1 0 14996 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0728_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 15732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0729_
timestamp 1694700623
transform -1 0 15640 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0730_
timestamp 1694700623
transform 1 0 16100 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0731_
timestamp 1694700623
transform -1 0 17572 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0732_
timestamp 1694700623
transform -1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0733_
timestamp 1694700623
transform 1 0 17480 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0735_
timestamp 1694700623
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0736_
timestamp 1694700623
transform -1 0 17388 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1694700623
transform -1 0 19320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0738_
timestamp 1694700623
transform -1 0 19044 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1694700623
transform -1 0 19044 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0740_
timestamp 1694700623
transform -1 0 18400 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0741_
timestamp 1694700623
transform 1 0 18124 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0742_
timestamp 1694700623
transform -1 0 18952 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0743_
timestamp 1694700623
transform -1 0 18860 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1694700623
transform -1 0 22540 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1694700623
transform 1 0 21252 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0746_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20424 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1694700623
transform 1 0 22448 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0748_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 22448 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0749_
timestamp 1694700623
transform -1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0750_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19688 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0751_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1694700623
transform 1 0 19412 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 1694700623
transform -1 0 19872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1694700623
transform 1 0 18032 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 1694700623
transform 1 0 17940 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1694700623
transform 1 0 12880 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 1694700623
transform 1 0 11592 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1694700623
transform 1 0 12144 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0759_
timestamp 1694700623
transform 1 0 11684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1694700623
transform 1 0 14168 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 1694700623
transform 1 0 13892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1694700623
transform 1 0 16652 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0763_
timestamp 1694700623
transform 1 0 15824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1694700623
transform 1 0 18216 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0765_
timestamp 1694700623
transform 1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0766_
timestamp 1694700623
transform -1 0 25484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0767_
timestamp 1694700623
transform 1 0 22816 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0768_
timestamp 1694700623
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0769_
timestamp 1694700623
transform 1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1694700623
transform -1 0 24932 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1694700623
transform -1 0 26036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0772_
timestamp 1694700623
transform 1 0 24932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0773_
timestamp 1694700623
transform 1 0 25300 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0774_
timestamp 1694700623
transform -1 0 25852 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 1694700623
transform 1 0 26036 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _0776_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 27508 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1694700623
transform 1 0 27416 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0778_
timestamp 1694700623
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0779_
timestamp 1694700623
transform 1 0 11776 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0780_
timestamp 1694700623
transform -1 0 14720 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0781_
timestamp 1694700623
transform 1 0 10672 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0782_
timestamp 1694700623
transform 1 0 10764 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0783_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11132 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0784_
timestamp 1694700623
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0785_
timestamp 1694700623
transform 1 0 11224 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0786_
timestamp 1694700623
transform 1 0 12328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _0787_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11224 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_2  _0788_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13708 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0789_
timestamp 1694700623
transform -1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0790_
timestamp 1694700623
transform 1 0 11868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0791_
timestamp 1694700623
transform 1 0 12880 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1694700623
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1694700623
transform -1 0 13984 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0794_
timestamp 1694700623
transform 1 0 14720 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0795_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 14536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0796_
timestamp 1694700623
transform 1 0 14352 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0797_
timestamp 1694700623
transform 1 0 11592 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0798_
timestamp 1694700623
transform 1 0 12696 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1694700623
transform -1 0 19228 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0800_
timestamp 1694700623
transform -1 0 17204 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0801_
timestamp 1694700623
transform 1 0 17296 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_2  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 18032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _0803_
timestamp 1694700623
transform 1 0 12788 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0804_
timestamp 1694700623
transform -1 0 16468 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1694700623
transform -1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0806_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1694700623
transform -1 0 16008 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0808_
timestamp 1694700623
transform 1 0 15180 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _0809_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14352 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_2  _0810_
timestamp 1694700623
transform 1 0 12236 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _0811_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 13984 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0812_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14444 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0813_
timestamp 1694700623
transform -1 0 20700 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0814_
timestamp 1694700623
transform -1 0 18308 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0815_
timestamp 1694700623
transform 1 0 18216 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0816_
timestamp 1694700623
transform -1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1694700623
transform -1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0818_
timestamp 1694700623
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0819_
timestamp 1694700623
transform -1 0 17572 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0820_
timestamp 1694700623
transform -1 0 14904 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0821_
timestamp 1694700623
transform 1 0 11408 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0822_
timestamp 1694700623
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1694700623
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0824_
timestamp 1694700623
transform 1 0 14444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0825_
timestamp 1694700623
transform 1 0 10764 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1694700623
transform 1 0 11592 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1694700623
transform 1 0 11316 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0828_
timestamp 1694700623
transform -1 0 12696 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0829_
timestamp 1694700623
transform -1 0 12144 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0831_
timestamp 1694700623
transform -1 0 23920 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0832_
timestamp 1694700623
transform 1 0 20884 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0833_
timestamp 1694700623
transform -1 0 22448 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0834_
timestamp 1694700623
transform -1 0 20332 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0835_
timestamp 1694700623
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 1694700623
transform 1 0 20332 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0837_
timestamp 1694700623
transform 1 0 19412 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0838_
timestamp 1694700623
transform 1 0 19964 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1694700623
transform -1 0 17572 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0840_
timestamp 1694700623
transform -1 0 17848 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0841_
timestamp 1694700623
transform 1 0 16560 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0842_
timestamp 1694700623
transform 1 0 16652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 21160 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1694700623
transform 1 0 17756 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0845_
timestamp 1694700623
transform -1 0 19504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0846_
timestamp 1694700623
transform -1 0 20240 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 15640 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0848_
timestamp 1694700623
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0849_
timestamp 1694700623
transform -1 0 18308 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0850_
timestamp 1694700623
transform -1 0 18676 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0851_
timestamp 1694700623
transform -1 0 18216 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0853_
timestamp 1694700623
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0854_
timestamp 1694700623
transform 1 0 20516 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0855_
timestamp 1694700623
transform -1 0 21620 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0856_
timestamp 1694700623
transform 1 0 19780 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0857_
timestamp 1694700623
transform -1 0 19872 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0858_
timestamp 1694700623
transform 1 0 32936 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0859_
timestamp 1694700623
transform 1 0 32660 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0860_
timestamp 1694700623
transform 1 0 33212 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0861_
timestamp 1694700623
transform -1 0 33948 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0862_
timestamp 1694700623
transform 1 0 32384 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0863_
timestamp 1694700623
transform -1 0 32660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0864_
timestamp 1694700623
transform 1 0 28704 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0865_
timestamp 1694700623
transform 1 0 28244 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0866_
timestamp 1694700623
transform 1 0 29532 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0867_
timestamp 1694700623
transform -1 0 30268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0868_
timestamp 1694700623
transform -1 0 30176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1694700623
transform 1 0 30544 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0870_
timestamp 1694700623
transform 1 0 27968 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0871_
timestamp 1694700623
transform 1 0 28796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0872_
timestamp 1694700623
transform 1 0 32108 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0873_
timestamp 1694700623
transform 1 0 31924 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0874_
timestamp 1694700623
transform 1 0 31464 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0875_
timestamp 1694700623
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1694700623
transform -1 0 30544 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 1694700623
transform 1 0 30912 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0878_
timestamp 1694700623
transform 1 0 31280 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0879_
timestamp 1694700623
transform -1 0 32292 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0880_
timestamp 1694700623
transform -1 0 31464 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0881_
timestamp 1694700623
transform 1 0 30176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0882_
timestamp 1694700623
transform 1 0 28888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0883_
timestamp 1694700623
transform -1 0 30912 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0884_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 30452 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0885_
timestamp 1694700623
transform 1 0 27324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0886_
timestamp 1694700623
transform 1 0 25852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0887_
timestamp 1694700623
transform 1 0 27876 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1694700623
transform -1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1694700623
transform -1 0 28244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0890_
timestamp 1694700623
transform 1 0 27968 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0891_
timestamp 1694700623
transform 1 0 23552 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0892_
timestamp 1694700623
transform -1 0 25852 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0893_
timestamp 1694700623
transform 1 0 25484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1694700623
transform -1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1694700623
transform 1 0 25852 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1694700623
transform 1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1694700623
transform -1 0 25024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0898_
timestamp 1694700623
transform 1 0 23368 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1694700623
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0900_
timestamp 1694700623
transform 1 0 24564 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0901_
timestamp 1694700623
transform 1 0 25944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0902_
timestamp 1694700623
transform 1 0 27968 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0903_
timestamp 1694700623
transform 1 0 27416 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0904_
timestamp 1694700623
transform 1 0 31188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0905_
timestamp 1694700623
transform -1 0 33120 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1694700623
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 31832 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0908_
timestamp 1694700623
transform -1 0 25760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0909_
timestamp 1694700623
transform 1 0 24748 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1694700623
transform -1 0 27968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0911_
timestamp 1694700623
transform 1 0 27968 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1694700623
transform 1 0 28612 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1694700623
transform 1 0 33028 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0914_
timestamp 1694700623
transform 1 0 32292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0915_
timestamp 1694700623
transform 1 0 32844 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0916_
timestamp 1694700623
transform 1 0 33948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1694700623
transform 1 0 32936 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0918_
timestamp 1694700623
transform -1 0 33948 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1694700623
transform 1 0 32844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1694700623
transform -1 0 33396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0921_
timestamp 1694700623
transform 1 0 32108 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1694700623
transform 1 0 33856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1694700623
transform -1 0 33212 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1694700623
transform -1 0 32936 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0925_
timestamp 1694700623
transform -1 0 32108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1694700623
transform -1 0 31740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _0927_
timestamp 1694700623
transform 1 0 28336 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1694700623
transform -1 0 29072 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0929_
timestamp 1694700623
transform -1 0 28888 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0930_
timestamp 1694700623
transform 1 0 28060 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1694700623
transform 1 0 28520 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0932_
timestamp 1694700623
transform 1 0 29716 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0933_
timestamp 1694700623
transform -1 0 30728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1694700623
transform 1 0 30636 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0935_
timestamp 1694700623
transform -1 0 31004 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0936_
timestamp 1694700623
transform -1 0 30912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1694700623
transform -1 0 29992 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 28612 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0939_
timestamp 1694700623
transform 1 0 32292 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1694700623
transform 1 0 28980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0941_
timestamp 1694700623
transform -1 0 29348 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1694700623
transform -1 0 27968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1694700623
transform 1 0 27968 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0944_
timestamp 1694700623
transform -1 0 29256 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0945_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 25944 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0946_
timestamp 1694700623
transform 1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1694700623
transform 1 0 24748 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o311ai_4  _0948_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 27600 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _0949_
timestamp 1694700623
transform 1 0 23276 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0950_
timestamp 1694700623
transform 1 0 23368 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0951_
timestamp 1694700623
transform 1 0 24564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0952_
timestamp 1694700623
transform 1 0 20884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0953_
timestamp 1694700623
transform -1 0 21620 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0954_
timestamp 1694700623
transform 1 0 23920 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 21160 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp 1694700623
transform 1 0 21620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1694700623
transform -1 0 24196 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0958_
timestamp 1694700623
transform 1 0 15180 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0959_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0960_
timestamp 1694700623
transform 1 0 11592 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0961_
timestamp 1694700623
transform 1 0 12328 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0962_
timestamp 1694700623
transform -1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0963_
timestamp 1694700623
transform 1 0 17848 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1694700623
transform 1 0 20608 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1694700623
transform -1 0 22080 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0966_
timestamp 1694700623
transform 1 0 20976 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0967_
timestamp 1694700623
transform 1 0 26956 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0968_
timestamp 1694700623
transform -1 0 27968 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0969_
timestamp 1694700623
transform 1 0 32660 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0970_
timestamp 1694700623
transform -1 0 33304 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1694700623
transform -1 0 28152 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0972_
timestamp 1694700623
transform -1 0 26496 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 25944 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and4_1  _0974_
timestamp 1694700623
transform -1 0 24564 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0975_
timestamp 1694700623
transform 1 0 23276 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0976_
timestamp 1694700623
transform 1 0 23276 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0977_
timestamp 1694700623
transform -1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0978_
timestamp 1694700623
transform 1 0 20516 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0979_
timestamp 1694700623
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 21712 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _0981_
timestamp 1694700623
transform 1 0 21068 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0982_
timestamp 1694700623
transform 1 0 22448 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1694700623
transform 1 0 22080 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0984_
timestamp 1694700623
transform 1 0 28520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0985_
timestamp 1694700623
transform 1 0 25852 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0986_
timestamp 1694700623
transform -1 0 25852 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0987_
timestamp 1694700623
transform -1 0 24104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0988_
timestamp 1694700623
transform 1 0 23184 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0989_
timestamp 1694700623
transform 1 0 20700 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0990_
timestamp 1694700623
transform -1 0 24472 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 1694700623
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1694700623
transform 1 0 21344 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0993_
timestamp 1694700623
transform 1 0 25944 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0994_
timestamp 1694700623
transform -1 0 27508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 1694700623
transform 1 0 27600 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0996_
timestamp 1694700623
transform 1 0 27048 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0997_
timestamp 1694700623
transform 1 0 25576 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0998_
timestamp 1694700623
transform 1 0 20792 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 1694700623
transform 1 0 26956 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1694700623
transform 1 0 27048 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1694700623
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1694700623
transform -1 0 27232 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1003_
timestamp 1694700623
transform -1 0 25944 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1004_
timestamp 1694700623
transform 1 0 27876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1005_
timestamp 1694700623
transform 1 0 25300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1694700623
transform 1 0 26036 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1694700623
transform 1 0 24656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1008_
timestamp 1694700623
transform 1 0 29532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1009_
timestamp 1694700623
transform 1 0 30084 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1010_
timestamp 1694700623
transform 1 0 29992 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1011_
timestamp 1694700623
transform 1 0 28888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1012_
timestamp 1694700623
transform 1 0 28244 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1013_
timestamp 1694700623
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1014_
timestamp 1694700623
transform 1 0 27692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1015_
timestamp 1694700623
transform -1 0 28520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1694700623
transform 1 0 26588 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1694700623
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1018_
timestamp 1694700623
transform -1 0 30912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1019_
timestamp 1694700623
transform 1 0 29256 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1020_
timestamp 1694700623
transform -1 0 30636 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1694700623
transform 1 0 29624 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1694700623
transform -1 0 29808 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1694700623
transform 1 0 31372 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1024_
timestamp 1694700623
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1025_
timestamp 1694700623
transform 1 0 32108 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1026_
timestamp 1694700623
transform 1 0 33304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1027_
timestamp 1694700623
transform -1 0 32844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1028_
timestamp 1694700623
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1694700623
transform 1 0 32108 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1694700623
transform 1 0 31280 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1031_
timestamp 1694700623
transform -1 0 31280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1032_
timestamp 1694700623
transform -1 0 33212 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1033_
timestamp 1694700623
transform 1 0 30636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp 1694700623
transform 1 0 30084 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1694700623
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1036_
timestamp 1694700623
transform 1 0 27600 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1037_
timestamp 1694700623
transform 1 0 27968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1694700623
transform 1 0 31464 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1039_
timestamp 1694700623
transform 1 0 30452 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1040_
timestamp 1694700623
transform -1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1041_
timestamp 1694700623
transform 1 0 30728 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1042_
timestamp 1694700623
transform -1 0 32660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 1694700623
transform -1 0 33488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1044_
timestamp 1694700623
transform -1 0 31188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1045_
timestamp 1694700623
transform 1 0 21436 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1046_
timestamp 1694700623
transform 1 0 30268 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1694700623
transform -1 0 29808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1048_
timestamp 1694700623
transform -1 0 31372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1049_
timestamp 1694700623
transform 1 0 29532 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1050_
timestamp 1694700623
transform 1 0 29624 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1051_
timestamp 1694700623
transform 1 0 29440 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1694700623
transform 1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1053_
timestamp 1694700623
transform 1 0 31372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1694700623
transform 1 0 31188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1055_
timestamp 1694700623
transform -1 0 32752 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1056_
timestamp 1694700623
transform -1 0 20792 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1057_
timestamp 1694700623
transform 1 0 20332 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1058_
timestamp 1694700623
transform 1 0 25208 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1059_
timestamp 1694700623
transform 1 0 27600 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1060_
timestamp 1694700623
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1061_
timestamp 1694700623
transform -1 0 21252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 1694700623
transform 1 0 27048 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1063_
timestamp 1694700623
transform -1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1064_
timestamp 1694700623
transform 1 0 26956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1694700623
transform 1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1694700623
transform -1 0 30912 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1067_
timestamp 1694700623
transform 1 0 28704 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1068_
timestamp 1694700623
transform -1 0 30452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 1694700623
transform 1 0 29624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1694700623
transform -1 0 29624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1071_
timestamp 1694700623
transform -1 0 27876 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1072_
timestamp 1694700623
transform -1 0 27968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1073_
timestamp 1694700623
transform 1 0 29164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 29348 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1075_
timestamp 1694700623
transform 1 0 28796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1076_
timestamp 1694700623
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1077_
timestamp 1694700623
transform -1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1078_
timestamp 1694700623
transform 1 0 29808 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1079_
timestamp 1694700623
transform -1 0 29808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1080_
timestamp 1694700623
transform 1 0 27048 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1081_
timestamp 1694700623
transform 1 0 25300 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1082_
timestamp 1694700623
transform 1 0 25760 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1083_
timestamp 1694700623
transform 1 0 26128 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1084_
timestamp 1694700623
transform -1 0 27600 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1085_
timestamp 1694700623
transform 1 0 26680 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1086_
timestamp 1694700623
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1694700623
transform -1 0 25668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp 1694700623
transform -1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1694700623
transform 1 0 24748 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1090_
timestamp 1694700623
transform 1 0 25392 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 1694700623
transform 1 0 25760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1092_
timestamp 1694700623
transform -1 0 25760 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1694700623
transform 1 0 24380 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1694700623
transform 1 0 23184 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1095_
timestamp 1694700623
transform 1 0 22632 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1096_
timestamp 1694700623
transform -1 0 26496 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1097_
timestamp 1694700623
transform -1 0 23920 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1098_
timestamp 1694700623
transform 1 0 22264 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1099_
timestamp 1694700623
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1100_
timestamp 1694700623
transform -1 0 15640 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1101_
timestamp 1694700623
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1102_
timestamp 1694700623
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1103_
timestamp 1694700623
transform 1 0 20148 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1104_
timestamp 1694700623
transform 1 0 21988 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1105_
timestamp 1694700623
transform 1 0 20792 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1106_
timestamp 1694700623
transform -1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1107_
timestamp 1694700623
transform -1 0 23368 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1108_
timestamp 1694700623
transform -1 0 23368 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1694700623
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1110_
timestamp 1694700623
transform -1 0 23644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1111_
timestamp 1694700623
transform 1 0 21436 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1112_
timestamp 1694700623
transform 1 0 20516 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1113_
timestamp 1694700623
transform -1 0 23092 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1114_
timestamp 1694700623
transform 1 0 21620 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1115_
timestamp 1694700623
transform -1 0 21712 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1116_
timestamp 1694700623
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1117_
timestamp 1694700623
transform 1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1118_
timestamp 1694700623
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1119_
timestamp 1694700623
transform -1 0 18216 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1120_
timestamp 1694700623
transform 1 0 21068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1121_
timestamp 1694700623
transform -1 0 21160 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1122_
timestamp 1694700623
transform 1 0 18216 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1123_
timestamp 1694700623
transform -1 0 16836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1124_
timestamp 1694700623
transform 1 0 16836 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1694700623
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1126_
timestamp 1694700623
transform -1 0 20332 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1127_
timestamp 1694700623
transform 1 0 18584 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1128_
timestamp 1694700623
transform -1 0 20056 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1129_
timestamp 1694700623
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1130_
timestamp 1694700623
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1694700623
transform -1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1132_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 14904 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 1694700623
transform -1 0 15824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1134_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16744 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1135_
timestamp 1694700623
transform 1 0 18768 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1136_
timestamp 1694700623
transform 1 0 15088 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1694700623
transform 1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1138_
timestamp 1694700623
transform 1 0 18492 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1139_
timestamp 1694700623
transform 1 0 19504 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1140_
timestamp 1694700623
transform -1 0 20332 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1694700623
transform 1 0 19964 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1694700623
transform 1 0 16376 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1143_
timestamp 1694700623
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1144_
timestamp 1694700623
transform 1 0 15824 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1145_
timestamp 1694700623
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1146_
timestamp 1694700623
transform 1 0 16192 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1147_
timestamp 1694700623
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1694700623
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1149_
timestamp 1694700623
transform -1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1150_
timestamp 1694700623
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1151_
timestamp 1694700623
transform -1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1694700623
transform 1 0 15548 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1153_
timestamp 1694700623
transform -1 0 14996 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1154_
timestamp 1694700623
transform 1 0 13432 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1694700623
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1156_
timestamp 1694700623
transform 1 0 11960 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1157_
timestamp 1694700623
transform 1 0 12052 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1158_
timestamp 1694700623
transform -1 0 13156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1159_
timestamp 1694700623
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1694700623
transform 1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1162_
timestamp 1694700623
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1163_
timestamp 1694700623
transform -1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1164_
timestamp 1694700623
transform 1 0 14536 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1165_
timestamp 1694700623
transform -1 0 12328 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1166_
timestamp 1694700623
transform 1 0 12512 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1167_
timestamp 1694700623
transform 1 0 13064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 1694700623
transform 1 0 9384 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1694700623
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1170_
timestamp 1694700623
transform 1 0 11868 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1694700623
transform 1 0 11776 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1172_
timestamp 1694700623
transform -1 0 14352 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1173_
timestamp 1694700623
transform -1 0 13248 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1174_
timestamp 1694700623
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1694700623
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1176_
timestamp 1694700623
transform 1 0 13340 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1177_
timestamp 1694700623
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1178_
timestamp 1694700623
transform 1 0 13800 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 1694700623
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1180_
timestamp 1694700623
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1181_
timestamp 1694700623
transform 1 0 12236 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1182_
timestamp 1694700623
transform -1 0 14996 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1183_
timestamp 1694700623
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1694700623
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1185_
timestamp 1694700623
transform -1 0 15364 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1186_
timestamp 1694700623
transform 1 0 12052 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1187_
timestamp 1694700623
transform -1 0 14720 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1188_
timestamp 1694700623
transform 1 0 9568 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1189_
timestamp 1694700623
transform 1 0 9016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1190_
timestamp 1694700623
transform 1 0 14720 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 1694700623
transform 1 0 14720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1192_
timestamp 1694700623
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1193_
timestamp 1694700623
transform -1 0 15732 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1194_
timestamp 1694700623
transform -1 0 14904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1195_
timestamp 1694700623
transform 1 0 14904 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1196_
timestamp 1694700623
transform -1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1197_
timestamp 1694700623
transform 1 0 11960 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1694700623
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1199_
timestamp 1694700623
transform 1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1694700623
transform -1 0 16192 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1201_
timestamp 1694700623
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1202_
timestamp 1694700623
transform 1 0 15364 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1203_
timestamp 1694700623
transform 1 0 15364 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1204_
timestamp 1694700623
transform 1 0 12144 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1694700623
transform -1 0 11868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1694700623
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1207_
timestamp 1694700623
transform -1 0 18400 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1208_
timestamp 1694700623
transform 1 0 16652 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1209_
timestamp 1694700623
transform -1 0 18032 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1210_
timestamp 1694700623
transform 1 0 16928 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1694700623
transform -1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1212_
timestamp 1694700623
transform -1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1694700623
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1214_
timestamp 1694700623
transform 1 0 20148 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1694700623
transform -1 0 9936 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1217_
timestamp 1694700623
transform 1 0 8464 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1218_
timestamp 1694700623
transform -1 0 9568 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1219_
timestamp 1694700623
transform -1 0 5152 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1220_
timestamp 1694700623
transform 1 0 2852 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3404 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1694700623
transform 1 0 5980 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _1223_
timestamp 1694700623
transform 1 0 5520 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7728 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 9660 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 9752 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8648 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1228_
timestamp 1694700623
transform 1 0 8004 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1229_
timestamp 1694700623
transform -1 0 8372 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  _1230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6992 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1231_
timestamp 1694700623
transform -1 0 23368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp 1694700623
transform -1 0 23000 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1233_
timestamp 1694700623
transform 1 0 20240 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1234_
timestamp 1694700623
transform -1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1235_
timestamp 1694700623
transform -1 0 20700 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1694700623
transform -1 0 20148 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1237_
timestamp 1694700623
transform 1 0 21988 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1694700623
transform -1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1239_
timestamp 1694700623
transform 1 0 21804 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1240_
timestamp 1694700623
transform -1 0 22448 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1241_
timestamp 1694700623
transform -1 0 20240 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1242_
timestamp 1694700623
transform 1 0 18860 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 1694700623
transform 1 0 16744 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1244_
timestamp 1694700623
transform 1 0 14996 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1245_
timestamp 1694700623
transform -1 0 14628 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1246_
timestamp 1694700623
transform -1 0 13984 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 24104 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1248_
timestamp 1694700623
transform 1 0 18584 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1694700623
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1250_
timestamp 1694700623
transform -1 0 18032 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1694700623
transform 1 0 11960 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1694700623
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1694700623
transform 1 0 9384 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1254_
timestamp 1694700623
transform -1 0 9844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1694700623
transform -1 0 8832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1694700623
transform 1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1257_
timestamp 1694700623
transform -1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1258_
timestamp 1694700623
transform 1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1259_
timestamp 1694700623
transform -1 0 24380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1694700623
transform -1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1694700623
transform -1 0 21528 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1694700623
transform -1 0 16468 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1263_
timestamp 1694700623
transform -1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1694700623
transform -1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1694700623
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1266_
timestamp 1694700623
transform 1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1694700623
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1268_
timestamp 1694700623
transform 1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1269_
timestamp 1694700623
transform 1 0 29992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1270_
timestamp 1694700623
transform 1 0 24380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 1694700623
transform 1 0 30176 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1694700623
transform -1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1694700623
transform 1 0 28612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1694700623
transform 1 0 30728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1275_
timestamp 1694700623
transform 1 0 30176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1694700623
transform 1 0 31556 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1694700623
transform 1 0 30452 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1694700623
transform 1 0 26312 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1694700623
transform 1 0 25392 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1694700623
transform -1 0 28428 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1281_
timestamp 1694700623
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1694700623
transform 1 0 22632 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 1694700623
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1694700623
transform -1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1694700623
transform -1 0 17480 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1694700623
transform 1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1694700623
transform -1 0 12604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1694700623
transform -1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1694700623
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1694700623
transform -1 0 21528 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1694700623
transform 1 0 19964 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1292_
timestamp 1694700623
transform 1 0 10856 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1293_
timestamp 1694700623
transform 1 0 12144 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1694700623
transform 1 0 21252 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1694700623
transform 1 0 23368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1296_
timestamp 1694700623
transform 1 0 22172 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1297_
timestamp 1694700623
transform 1 0 22816 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1694700623
transform -1 0 22816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1299_
timestamp 1694700623
transform 1 0 10304 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1694700623
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1694700623
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1302_
timestamp 1694700623
transform 1 0 2668 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1303_
timestamp 1694700623
transform 1 0 4968 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1304_
timestamp 1694700623
transform 1 0 5060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1305_
timestamp 1694700623
transform -1 0 5704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1694700623
transform -1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1694700623
transform 1 0 7176 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1694700623
transform -1 0 8556 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1694700623
transform 1 0 7820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1694700623
transform -1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1311_
timestamp 1694700623
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1312_
timestamp 1694700623
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1694700623
transform 1 0 9752 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_
timestamp 1694700623
transform 1 0 9568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1315_
timestamp 1694700623
transform -1 0 8740 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1316_
timestamp 1694700623
transform 1 0 7636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1317_
timestamp 1694700623
transform 1 0 7544 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1318_
timestamp 1694700623
transform 1 0 9384 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1319_
timestamp 1694700623
transform -1 0 11316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1320_
timestamp 1694700623
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1321_
timestamp 1694700623
transform -1 0 6164 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1322_
timestamp 1694700623
transform -1 0 5704 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1323_
timestamp 1694700623
transform 1 0 5060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1324_
timestamp 1694700623
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1325_
timestamp 1694700623
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1326_
timestamp 1694700623
transform -1 0 4324 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1694700623
transform -1 0 3680 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1694700623
transform -1 0 2852 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp 1694700623
transform -1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1330_
timestamp 1694700623
transform -1 0 2300 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1331_
timestamp 1694700623
transform 1 0 1380 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1332_
timestamp 1694700623
transform -1 0 4692 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1333_
timestamp 1694700623
transform -1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1694700623
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1335_
timestamp 1694700623
transform -1 0 5980 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1336_
timestamp 1694700623
transform 1 0 5060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1337_
timestamp 1694700623
transform -1 0 5520 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1338_
timestamp 1694700623
transform 1 0 6348 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1339_
timestamp 1694700623
transform 1 0 7084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1340_
timestamp 1694700623
transform 1 0 6808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1341_
timestamp 1694700623
transform 1 0 4968 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1342_
timestamp 1694700623
transform -1 0 6256 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1343_
timestamp 1694700623
transform -1 0 6992 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1344_
timestamp 1694700623
transform 1 0 7084 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1345_
timestamp 1694700623
transform 1 0 8188 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1694700623
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1694700623
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1348_
timestamp 1694700623
transform 1 0 9752 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1349_
timestamp 1694700623
transform 1 0 10580 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1694700623
transform -1 0 10488 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8924 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__o21ai_1  _1352_
timestamp 1694700623
transform -1 0 11408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1353_
timestamp 1694700623
transform -1 0 7636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1694700623
transform -1 0 7360 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1694700623
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1694700623
transform 1 0 17572 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1694700623
transform -1 0 15824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1694700623
transform -1 0 12696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1694700623
transform 1 0 13248 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1360_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 21068 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 1694700623
transform 1 0 16652 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 11500 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1363_
timestamp 1694700623
transform 1 0 8924 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1364_
timestamp 1694700623
transform 1 0 8464 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1365_
timestamp 1694700623
transform 1 0 7728 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1366_
timestamp 1694700623
transform 1 0 7728 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1367_
timestamp 1694700623
transform 1 0 8924 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1368_
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1369_
timestamp 1694700623
transform 1 0 11592 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1370_
timestamp 1694700623
transform 1 0 15548 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 1694700623
transform 1 0 19412 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1694700623
transform 1 0 14996 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1373_
timestamp 1694700623
transform 1 0 15732 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1374_
timestamp 1694700623
transform 1 0 21804 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1375_
timestamp 1694700623
transform -1 0 25576 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1376_
timestamp 1694700623
transform 1 0 21160 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1377_
timestamp 1694700623
transform 1 0 22540 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 1694700623
transform 1 0 26220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1379_
timestamp 1694700623
transform 1 0 29532 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1380_
timestamp 1694700623
transform 1 0 29532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1381_
timestamp 1694700623
transform 1 0 25024 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1382_
timestamp 1694700623
transform 1 0 27600 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1383_
timestamp 1694700623
transform 1 0 29808 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1384_
timestamp 1694700623
transform 1 0 29256 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 1694700623
transform 1 0 30728 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 1694700623
transform 1 0 29440 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1387_
timestamp 1694700623
transform 1 0 25392 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 1694700623
transform 1 0 24380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1389_
timestamp 1694700623
transform 1 0 26312 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1694700623
transform 1 0 20792 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1391_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 21528 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1392_
timestamp 1694700623
transform 1 0 17296 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1393_
timestamp 1694700623
transform 1 0 15364 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1394_
timestamp 1694700623
transform 1 0 13432 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1395_
timestamp 1694700623
transform 1 0 11500 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1396_
timestamp 1694700623
transform 1 0 11040 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1397_
timestamp 1694700623
transform 1 0 17572 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1398_
timestamp 1694700623
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1399_
timestamp 1694700623
transform 1 0 18952 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1400_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 12880 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1401_
timestamp 1694700623
transform 1 0 20240 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1694700623
transform -1 0 24104 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1694700623
transform 1 0 24104 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1694700623
transform -1 0 24104 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1694700623
transform 1 0 19320 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1694700623
transform 1 0 10580 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1407_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3680 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1694700623
transform 1 0 3312 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1694700623
transform 1 0 4324 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1694700623
transform -1 0 7268 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1694700623
transform 1 0 7268 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1694700623
transform -1 0 11132 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1694700623
transform -1 0 10396 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1694700623
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1694700623
transform 1 0 9108 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1694700623
transform -1 0 11040 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1694700623
transform 1 0 4416 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1694700623
transform -1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1694700623
transform 1 0 3772 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1694700623
transform 1 0 1656 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1694700623
transform -1 0 3128 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1694700623
transform -1 0 3680 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1423_
timestamp 1694700623
transform 1 0 4600 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1424_
timestamp 1694700623
transform 1 0 3772 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1425_
timestamp 1694700623
transform 1 0 6348 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1426_
timestamp 1694700623
transform -1 0 6256 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1427_
timestamp 1694700623
transform -1 0 7728 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1428_
timestamp 1694700623
transform -1 0 8924 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1429_
timestamp 1694700623
transform 1 0 8280 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1430_
timestamp 1694700623
transform -1 0 11132 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1431_
timestamp 1694700623
transform 1 0 8372 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1432_
timestamp 1694700623
transform 1 0 6532 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1433_
timestamp 1694700623
transform 1 0 9752 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_2  _1434_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 17756 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1435_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16376 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1436_
timestamp 1694700623
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1437_
timestamp 1694700623
transform 1 0 10764 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1438_
timestamp 1694700623
transform 1 0 10488 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1439_
timestamp 1694700623
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1440_
timestamp 1694700623
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1441_
timestamp 1694700623
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1442_
timestamp 1694700623
transform 1 0 10488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1443_
timestamp 1694700623
transform 1 0 14168 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1444_
timestamp 1694700623
transform -1 0 19044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1445_
timestamp 1694700623
transform -1 0 22172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1446_
timestamp 1694700623
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1447_
timestamp 1694700623
transform 1 0 18584 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1448_
timestamp 1694700623
transform -1 0 23736 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_2  _1449_
timestamp 1694700623
transform -1 0 25576 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1450_
timestamp 1694700623
transform 1 0 23000 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1451_
timestamp 1694700623
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1452_
timestamp 1694700623
transform -1 0 29716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1453_
timestamp 1694700623
transform -1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1454_
timestamp 1694700623
transform -1 0 34224 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1455_
timestamp 1694700623
transform -1 0 28244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1456_
timestamp 1694700623
transform -1 0 34868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1457_
timestamp 1694700623
transform 1 0 33304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1458_
timestamp 1694700623
transform 1 0 33304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1459_
timestamp 1694700623
transform -1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1460_
timestamp 1694700623
transform -1 0 29440 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1461_
timestamp 1694700623
transform -1 0 28336 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1462_
timestamp 1694700623
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1463_
timestamp 1694700623
transform -1 0 26036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1464_
timestamp 1694700623
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1465_
timestamp 1694700623
transform 1 0 23552 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 19044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1467_
timestamp 1694700623
transform -1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1468_
timestamp 1694700623
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1469_
timestamp 1694700623
transform -1 0 10948 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1470_
timestamp 1694700623
transform -1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1471_
timestamp 1694700623
transform -1 0 10212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1472_
timestamp 1694700623
transform -1 0 10120 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1473_
timestamp 1694700623
transform -1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1474_
timestamp 1694700623
transform 1 0 9844 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1475_
timestamp 1694700623
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1476_
timestamp 1694700623
transform 1 0 17296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1477_
timestamp 1694700623
transform 1 0 20608 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1478_
timestamp 1694700623
transform 1 0 16928 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1479_
timestamp 1694700623
transform 1 0 17756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1480_
timestamp 1694700623
transform 1 0 21988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1481_
timestamp 1694700623
transform 1 0 23828 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1482_
timestamp 1694700623
transform -1 0 24104 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1483_
timestamp 1694700623
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1484_
timestamp 1694700623
transform 1 0 28060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1485_
timestamp 1694700623
transform 1 0 30820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1486_
timestamp 1694700623
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1487_
timestamp 1694700623
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1488_
timestamp 1694700623
transform 1 0 32660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1489_
timestamp 1694700623
transform 1 0 32200 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1490_
timestamp 1694700623
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1491_
timestamp 1694700623
transform 1 0 32568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1492_
timestamp 1694700623
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1493_
timestamp 1694700623
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1494_
timestamp 1694700623
transform 1 0 24932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1495_
timestamp 1694700623
transform 1 0 24564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1496_
timestamp 1694700623
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1497_
timestamp 1694700623
transform 1 0 22448 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1498_
timestamp 1694700623
transform 1 0 20792 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1499_
timestamp 1694700623
transform 1 0 20332 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1500_
timestamp 1694700623
transform 1 0 18216 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1501_
timestamp 1694700623
transform 1 0 16560 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1502_
timestamp 1694700623
transform 1 0 14444 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1503_
timestamp 1694700623
transform -1 0 12420 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1504_
timestamp 1694700623
transform 1 0 12328 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clock
timestamp 1694700623
transform -1 0 10488 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clock
timestamp 1694700623
transform 1 0 11868 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clock
timestamp 1694700623
transform -1 0 10028 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clock
timestamp 1694700623
transform -1 0 12696 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clock
timestamp 1694700623
transform -1 0 23736 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clock
timestamp 1694700623
transform 1 0 25208 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clock
timestamp 1694700623
transform 1 0 18676 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clock
timestamp 1694700623
transform 1 0 23184 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  fanout9
timestamp 1694700623
transform -1 0 9568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout10
timestamp 1694700623
transform -1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1694700623
transform -1 0 18860 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1694700623
transform -1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout13
timestamp 1694700623
transform -1 0 24748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1694700623
transform 1 0 25024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1694700623
transform 1 0 25024 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1694700623
transform 1 0 22816 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1694700623
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1694700623
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1694700623
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1694700623
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1694700623
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1694700623
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1694700623
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1694700623
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1694700623
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1694700623
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1694700623
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1694700623
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1694700623
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1694700623
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1694700623
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1694700623
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1694700623
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1694700623
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1694700623
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1694700623
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1694700623
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1694700623
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1694700623
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1694700623
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1694700623
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1694700623
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1694700623
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1694700623
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1694700623
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1694700623
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1694700623
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1694700623
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1694700623
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1694700623
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1694700623
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1694700623
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1694700623
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1694700623
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_405 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1694700623
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1694700623
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1694700623
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1694700623
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1694700623
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1694700623
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1694700623
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1694700623
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1694700623
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1694700623
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1694700623
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1694700623
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1694700623
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1694700623
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1694700623
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1694700623
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1694700623
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1694700623
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1694700623
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1694700623
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1694700623
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1694700623
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1694700623
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1694700623
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1694700623
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1694700623
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1694700623
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1694700623
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1694700623
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1694700623
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1694700623
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1694700623
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1694700623
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1694700623
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1694700623
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1694700623
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1694700623
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1694700623
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1694700623
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_405
timestamp 1694700623
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1694700623
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1694700623
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1694700623
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1694700623
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1694700623
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1694700623
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1694700623
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1694700623
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1694700623
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1694700623
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1694700623
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1694700623
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1694700623
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1694700623
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1694700623
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1694700623
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1694700623
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1694700623
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1694700623
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1694700623
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1694700623
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1694700623
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1694700623
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1694700623
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1694700623
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1694700623
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1694700623
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1694700623
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1694700623
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1694700623
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1694700623
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1694700623
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1694700623
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1694700623
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1694700623
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1694700623
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1694700623
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1694700623
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1694700623
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_401
timestamp 1694700623
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1694700623
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1694700623
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1694700623
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1694700623
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1694700623
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1694700623
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1694700623
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1694700623
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1694700623
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1694700623
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1694700623
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1694700623
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1694700623
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1694700623
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1694700623
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1694700623
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1694700623
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1694700623
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1694700623
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1694700623
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1694700623
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1694700623
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1694700623
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1694700623
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1694700623
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1694700623
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1694700623
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1694700623
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1694700623
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1694700623
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1694700623
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1694700623
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1694700623
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1694700623
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1694700623
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1694700623
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1694700623
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1694700623
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1694700623
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1694700623
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_405
timestamp 1694700623
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1694700623
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1694700623
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1694700623
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1694700623
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1694700623
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1694700623
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1694700623
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1694700623
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1694700623
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1694700623
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1694700623
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1694700623
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1694700623
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1694700623
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1694700623
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1694700623
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1694700623
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1694700623
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1694700623
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1694700623
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1694700623
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1694700623
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1694700623
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1694700623
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1694700623
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1694700623
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1694700623
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1694700623
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1694700623
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1694700623
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1694700623
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1694700623
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1694700623
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1694700623
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1694700623
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1694700623
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1694700623
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1694700623
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1694700623
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_401
timestamp 1694700623
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1694700623
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1694700623
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1694700623
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1694700623
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1694700623
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1694700623
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1694700623
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1694700623
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1694700623
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1694700623
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1694700623
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1694700623
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1694700623
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1694700623
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1694700623
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1694700623
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1694700623
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1694700623
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1694700623
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1694700623
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1694700623
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1694700623
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1694700623
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1694700623
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1694700623
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1694700623
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1694700623
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1694700623
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1694700623
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1694700623
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1694700623
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1694700623
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1694700623
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1694700623
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1694700623
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1694700623
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1694700623
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1694700623
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1694700623
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1694700623
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1694700623
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 1694700623
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1694700623
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1694700623
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1694700623
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1694700623
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1694700623
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1694700623
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1694700623
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1694700623
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1694700623
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1694700623
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1694700623
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1694700623
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1694700623
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1694700623
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1694700623
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1694700623
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1694700623
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1694700623
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1694700623
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1694700623
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1694700623
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1694700623
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1694700623
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1694700623
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1694700623
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1694700623
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1694700623
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1694700623
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1694700623
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1694700623
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1694700623
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1694700623
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1694700623
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1694700623
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1694700623
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1694700623
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1694700623
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1694700623
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1694700623
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_401
timestamp 1694700623
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1694700623
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1694700623
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1694700623
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1694700623
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1694700623
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1694700623
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1694700623
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1694700623
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1694700623
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1694700623
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1694700623
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1694700623
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1694700623
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1694700623
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1694700623
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1694700623
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1694700623
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1694700623
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1694700623
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1694700623
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1694700623
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1694700623
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1694700623
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1694700623
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1694700623
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1694700623
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1694700623
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1694700623
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1694700623
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1694700623
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1694700623
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1694700623
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1694700623
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1694700623
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1694700623
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1694700623
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1694700623
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1694700623
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1694700623
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1694700623
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1694700623
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_405
timestamp 1694700623
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1694700623
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1694700623
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1694700623
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1694700623
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1694700623
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1694700623
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1694700623
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1694700623
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1694700623
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1694700623
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1694700623
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1694700623
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1694700623
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1694700623
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1694700623
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1694700623
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1694700623
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1694700623
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1694700623
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1694700623
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1694700623
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1694700623
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1694700623
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1694700623
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1694700623
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1694700623
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1694700623
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1694700623
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1694700623
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1694700623
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1694700623
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1694700623
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1694700623
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1694700623
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1694700623
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1694700623
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1694700623
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1694700623
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1694700623
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_401
timestamp 1694700623
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1694700623
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1694700623
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1694700623
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1694700623
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1694700623
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1694700623
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1694700623
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1694700623
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1694700623
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1694700623
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1694700623
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1694700623
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1694700623
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1694700623
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_161
timestamp 1694700623
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1694700623
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 1694700623
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp 1694700623
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_188
timestamp 1694700623
transform 1 0 18400 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_200
timestamp 1694700623
transform 1 0 19504 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_212
timestamp 1694700623
transform 1 0 20608 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1694700623
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1694700623
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1694700623
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1694700623
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1694700623
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1694700623
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_281
timestamp 1694700623
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_287
timestamp 1694700623
transform 1 0 27508 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_299
timestamp 1694700623
transform 1 0 28612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_311
timestamp 1694700623
transform 1 0 29716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_323
timestamp 1694700623
transform 1 0 30820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1694700623
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1694700623
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1694700623
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1694700623
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1694700623
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1694700623
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1694700623
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1694700623
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_405
timestamp 1694700623
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1694700623
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1694700623
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1694700623
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1694700623
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1694700623
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1694700623
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1694700623
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1694700623
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1694700623
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1694700623
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_127
timestamp 1694700623
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1694700623
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_154
timestamp 1694700623
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_180
timestamp 1694700623
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1694700623
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_197 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_208
timestamp 1694700623
transform 1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_224
timestamp 1694700623
transform 1 0 21712 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_236
timestamp 1694700623
transform 1 0 22816 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_242
timestamp 1694700623
transform 1 0 23368 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_246
timestamp 1694700623
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1694700623
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_265
timestamp 1694700623
transform 1 0 25484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_305
timestamp 1694700623
transform 1 0 29164 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1694700623
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1694700623
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1694700623
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1694700623
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1694700623
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1694700623
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1694700623
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1694700623
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1694700623
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_401
timestamp 1694700623
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1694700623
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1694700623
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1694700623
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1694700623
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1694700623
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1694700623
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1694700623
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1694700623
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1694700623
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1694700623
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1694700623
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1694700623
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1694700623
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_178
timestamp 1694700623
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_193
timestamp 1694700623
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1694700623
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1694700623
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_281
timestamp 1694700623
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_292
timestamp 1694700623
transform 1 0 27968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_298
timestamp 1694700623
transform 1 0 28520 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_311
timestamp 1694700623
transform 1 0 29716 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1694700623
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1694700623
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1694700623
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1694700623
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1694700623
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1694700623
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1694700623
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1694700623
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1694700623
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1694700623
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_401
timestamp 1694700623
transform 1 0 37996 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1694700623
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1694700623
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1694700623
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1694700623
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1694700623
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1694700623
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_97
timestamp 1694700623
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_101
timestamp 1694700623
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_114
timestamp 1694700623
transform 1 0 11592 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_126
timestamp 1694700623
transform 1 0 12696 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1694700623
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1694700623
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_149
timestamp 1694700623
transform 1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_162
timestamp 1694700623
transform 1 0 16008 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_177
timestamp 1694700623
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 1694700623
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_209
timestamp 1694700623
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_229
timestamp 1694700623
transform 1 0 22172 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_237
timestamp 1694700623
transform 1 0 22908 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_243
timestamp 1694700623
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1694700623
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_275
timestamp 1694700623
transform 1 0 26404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_287
timestamp 1694700623
transform 1 0 27508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_299
timestamp 1694700623
transform 1 0 28612 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_329
timestamp 1694700623
transform 1 0 31372 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_341
timestamp 1694700623
transform 1 0 32476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_353
timestamp 1694700623
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_361
timestamp 1694700623
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1694700623
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1694700623
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1694700623
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_401
timestamp 1694700623
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1694700623
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1694700623
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1694700623
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1694700623
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1694700623
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1694700623
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1694700623
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_81
timestamp 1694700623
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_92
timestamp 1694700623
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 1694700623
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1694700623
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_113
timestamp 1694700623
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_117
timestamp 1694700623
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1694700623
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_137
timestamp 1694700623
transform 1 0 13708 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_143
timestamp 1694700623
transform 1 0 14260 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_151
timestamp 1694700623
transform 1 0 14996 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_163
timestamp 1694700623
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1694700623
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1694700623
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1694700623
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_193
timestamp 1694700623
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_199
timestamp 1694700623
transform 1 0 19412 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_207
timestamp 1694700623
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 1694700623
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1694700623
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 1694700623
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_231
timestamp 1694700623
transform 1 0 22356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_237
timestamp 1694700623
transform 1 0 22908 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_250
timestamp 1694700623
transform 1 0 24104 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_262
timestamp 1694700623
transform 1 0 25208 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_269
timestamp 1694700623
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1694700623
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 1694700623
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_289
timestamp 1694700623
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_295
timestamp 1694700623
transform 1 0 28244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_307
timestamp 1694700623
transform 1 0 29348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_321
timestamp 1694700623
transform 1 0 30636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1694700623
transform 1 0 31740 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1694700623
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1694700623
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1694700623
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1694700623
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1694700623
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1694700623
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1694700623
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_405
timestamp 1694700623
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1694700623
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1694700623
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1694700623
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1694700623
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1694700623
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1694700623
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1694700623
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1694700623
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_118
timestamp 1694700623
transform 1 0 11960 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_131
timestamp 1694700623
transform 1 0 13156 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_146
timestamp 1694700623
transform 1 0 14536 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_158
timestamp 1694700623
transform 1 0 15640 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_171
timestamp 1694700623
transform 1 0 16836 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_179
timestamp 1694700623
transform 1 0 17572 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_185
timestamp 1694700623
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1694700623
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1694700623
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_205
timestamp 1694700623
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1694700623
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_253
timestamp 1694700623
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_271
timestamp 1694700623
transform 1 0 26036 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_279
timestamp 1694700623
transform 1 0 26772 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_288
timestamp 1694700623
transform 1 0 27600 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_300
timestamp 1694700623
transform 1 0 28704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1694700623
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_309
timestamp 1694700623
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_315
timestamp 1694700623
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_319
timestamp 1694700623
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_335
timestamp 1694700623
transform 1 0 31924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_347
timestamp 1694700623
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_359
timestamp 1694700623
transform 1 0 34132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1694700623
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1694700623
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1694700623
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1694700623
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_401
timestamp 1694700623
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1694700623
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1694700623
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1694700623
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1694700623
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1694700623
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1694700623
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1694700623
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1694700623
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1694700623
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1694700623
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1694700623
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1694700623
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_117
timestamp 1694700623
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_126
timestamp 1694700623
transform 1 0 12696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_134
timestamp 1694700623
transform 1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_148
timestamp 1694700623
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_169
timestamp 1694700623
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_191
timestamp 1694700623
transform 1 0 18676 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_199
timestamp 1694700623
transform 1 0 19412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_211
timestamp 1694700623
transform 1 0 20516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1694700623
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_228
timestamp 1694700623
transform 1 0 22080 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_240
timestamp 1694700623
transform 1 0 23184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_250
timestamp 1694700623
transform 1 0 24104 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_259
timestamp 1694700623
transform 1 0 24932 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_271
timestamp 1694700623
transform 1 0 26036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1694700623
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_281
timestamp 1694700623
transform 1 0 26956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1694700623
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1694700623
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1694700623
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1694700623
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1694700623
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1694700623
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1694700623
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1694700623
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_405
timestamp 1694700623
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1694700623
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1694700623
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1694700623
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1694700623
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1694700623
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1694700623
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1694700623
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1694700623
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1694700623
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1694700623
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1694700623
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 1694700623
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_126
timestamp 1694700623
transform 1 0 12696 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_132
timestamp 1694700623
transform 1 0 13248 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_149
timestamp 1694700623
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_164
timestamp 1694700623
transform 1 0 16192 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_176
timestamp 1694700623
transform 1 0 17296 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_187
timestamp 1694700623
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1694700623
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1694700623
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1694700623
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_221
timestamp 1694700623
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_229
timestamp 1694700623
transform 1 0 22172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_239
timestamp 1694700623
transform 1 0 23092 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 1694700623
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_256
timestamp 1694700623
transform 1 0 24656 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_270
timestamp 1694700623
transform 1 0 25944 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_282
timestamp 1694700623
transform 1 0 27048 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_288
timestamp 1694700623
transform 1 0 27600 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_301
timestamp 1694700623
transform 1 0 28796 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1694700623
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_320
timestamp 1694700623
transform 1 0 30544 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_332
timestamp 1694700623
transform 1 0 31648 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_344
timestamp 1694700623
transform 1 0 32752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_356
timestamp 1694700623
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1694700623
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1694700623
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1694700623
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_401
timestamp 1694700623
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1694700623
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1694700623
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1694700623
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1694700623
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1694700623
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1694700623
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1694700623
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1694700623
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_81
timestamp 1694700623
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1694700623
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1694700623
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1694700623
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1694700623
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_161
timestamp 1694700623
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1694700623
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_178
timestamp 1694700623
transform 1 0 17480 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_190
timestamp 1694700623
transform 1 0 18584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_198
timestamp 1694700623
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_206
timestamp 1694700623
transform 1 0 20056 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 1694700623
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1694700623
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1694700623
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1694700623
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1694700623
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_261
timestamp 1694700623
transform 1 0 25116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_274
timestamp 1694700623
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_293
timestamp 1694700623
transform 1 0 28060 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_304
timestamp 1694700623
transform 1 0 29072 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_316
timestamp 1694700623
transform 1 0 30176 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1694700623
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_343
timestamp 1694700623
transform 1 0 32660 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_355
timestamp 1694700623
transform 1 0 33764 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_367
timestamp 1694700623
transform 1 0 34868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_379
timestamp 1694700623
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1694700623
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1694700623
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_405
timestamp 1694700623
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1694700623
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1694700623
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1694700623
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1694700623
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1694700623
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1694700623
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1694700623
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_77
timestamp 1694700623
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_106
timestamp 1694700623
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_114
timestamp 1694700623
transform 1 0 11592 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_123
timestamp 1694700623
transform 1 0 12420 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1694700623
transform 1 0 13064 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1694700623
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 1694700623
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1694700623
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_171
timestamp 1694700623
transform 1 0 16836 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1694700623
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1694700623
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_228
timestamp 1694700623
transform 1 0 22080 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1694700623
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_253
timestamp 1694700623
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_264
timestamp 1694700623
transform 1 0 25392 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_273
timestamp 1694700623
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_285
timestamp 1694700623
transform 1 0 27324 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_291
timestamp 1694700623
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_303
timestamp 1694700623
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1694700623
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1694700623
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_321
timestamp 1694700623
transform 1 0 30636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_360
timestamp 1694700623
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1694700623
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1694700623
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1694700623
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_401
timestamp 1694700623
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1694700623
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1694700623
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1694700623
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1694700623
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1694700623
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1694700623
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1694700623
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1694700623
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_81
timestamp 1694700623
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_89
timestamp 1694700623
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 1694700623
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1694700623
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1694700623
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_129
timestamp 1694700623
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_138
timestamp 1694700623
transform 1 0 13800 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_150
timestamp 1694700623
transform 1 0 14904 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_159
timestamp 1694700623
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1694700623
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_182
timestamp 1694700623
transform 1 0 17848 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_197
timestamp 1694700623
transform 1 0 19228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_209
timestamp 1694700623
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_221
timestamp 1694700623
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_225
timestamp 1694700623
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1694700623
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_249
timestamp 1694700623
transform 1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_268
timestamp 1694700623
transform 1 0 25760 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_276
timestamp 1694700623
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 1694700623
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_297
timestamp 1694700623
transform 1 0 28428 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_324
timestamp 1694700623
transform 1 0 30912 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_342
timestamp 1694700623
transform 1 0 32568 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_354
timestamp 1694700623
transform 1 0 33672 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_366
timestamp 1694700623
transform 1 0 34776 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_378
timestamp 1694700623
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_390
timestamp 1694700623
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1694700623
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_405
timestamp 1694700623
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1694700623
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1694700623
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1694700623
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1694700623
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1694700623
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1694700623
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1694700623
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_77
timestamp 1694700623
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1694700623
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_98
timestamp 1694700623
transform 1 0 10120 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_112
timestamp 1694700623
transform 1 0 11408 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_120
timestamp 1694700623
transform 1 0 12144 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_125
timestamp 1694700623
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_129
timestamp 1694700623
transform 1 0 12972 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1694700623
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1694700623
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_177
timestamp 1694700623
transform 1 0 17388 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_188
timestamp 1694700623
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1694700623
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1694700623
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_228
timestamp 1694700623
transform 1 0 22080 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_242
timestamp 1694700623
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1694700623
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1694700623
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_268
timestamp 1694700623
transform 1 0 25760 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_280
timestamp 1694700623
transform 1 0 26864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_286
timestamp 1694700623
transform 1 0 27416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_291
timestamp 1694700623
transform 1 0 27876 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_296
timestamp 1694700623
transform 1 0 28336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_332
timestamp 1694700623
transform 1 0 31648 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_339
timestamp 1694700623
transform 1 0 32292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_351
timestamp 1694700623
transform 1 0 33396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1694700623
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1694700623
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1694700623
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1694700623
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_401
timestamp 1694700623
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1694700623
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1694700623
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1694700623
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1694700623
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1694700623
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1694700623
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1694700623
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_69
timestamp 1694700623
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_92
timestamp 1694700623
transform 1 0 9568 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1694700623
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_123
timestamp 1694700623
transform 1 0 12420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_135
timestamp 1694700623
transform 1 0 13524 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_156
timestamp 1694700623
transform 1 0 15456 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1694700623
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_177
timestamp 1694700623
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_182
timestamp 1694700623
transform 1 0 17848 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_193
timestamp 1694700623
transform 1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_197
timestamp 1694700623
transform 1 0 19228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_204
timestamp 1694700623
transform 1 0 19872 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_212
timestamp 1694700623
transform 1 0 20608 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 1694700623
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1694700623
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_234
timestamp 1694700623
transform 1 0 22632 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_245
timestamp 1694700623
transform 1 0 23644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_257
timestamp 1694700623
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_261
timestamp 1694700623
transform 1 0 25116 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_267
timestamp 1694700623
transform 1 0 25668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1694700623
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1694700623
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1694700623
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_305
timestamp 1694700623
transform 1 0 29164 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_319
timestamp 1694700623
transform 1 0 30452 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_344
timestamp 1694700623
transform 1 0 32752 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_356
timestamp 1694700623
transform 1 0 33856 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_368
timestamp 1694700623
transform 1 0 34960 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_380
timestamp 1694700623
transform 1 0 36064 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1694700623
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_405
timestamp 1694700623
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1694700623
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1694700623
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1694700623
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1694700623
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1694700623
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1694700623
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1694700623
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_77
timestamp 1694700623
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1694700623
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_94
timestamp 1694700623
transform 1 0 9752 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_106
timestamp 1694700623
transform 1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_122
timestamp 1694700623
transform 1 0 12328 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_132
timestamp 1694700623
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_147
timestamp 1694700623
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_151
timestamp 1694700623
transform 1 0 14996 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_165
timestamp 1694700623
transform 1 0 16284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_169
timestamp 1694700623
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_178
timestamp 1694700623
transform 1 0 17480 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_183
timestamp 1694700623
transform 1 0 17940 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_200
timestamp 1694700623
transform 1 0 19504 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_208
timestamp 1694700623
transform 1 0 20240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_220
timestamp 1694700623
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_224
timestamp 1694700623
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_239
timestamp 1694700623
transform 1 0 23092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1694700623
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_266
timestamp 1694700623
transform 1 0 25576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_278
timestamp 1694700623
transform 1 0 26680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_285
timestamp 1694700623
transform 1 0 27324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_293
timestamp 1694700623
transform 1 0 28060 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_304
timestamp 1694700623
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1694700623
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1694700623
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_319
timestamp 1694700623
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_323
timestamp 1694700623
transform 1 0 30820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_333
timestamp 1694700623
transform 1 0 31740 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_348
timestamp 1694700623
transform 1 0 33120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_360
timestamp 1694700623
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1694700623
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1694700623
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1694700623
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 1694700623
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1694700623
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1694700623
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1694700623
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1694700623
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1694700623
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1694700623
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1694700623
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1694700623
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1694700623
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1694700623
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1694700623
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1694700623
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_118
timestamp 1694700623
transform 1 0 11960 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_130
timestamp 1694700623
transform 1 0 13064 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_136
timestamp 1694700623
transform 1 0 13616 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1694700623
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1694700623
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1694700623
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 1694700623
transform 1 0 17388 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_190
timestamp 1694700623
transform 1 0 18584 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_202
timestamp 1694700623
transform 1 0 19688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1694700623
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1694700623
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_272
timestamp 1694700623
transform 1 0 26128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1694700623
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_290
timestamp 1694700623
transform 1 0 27784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_298
timestamp 1694700623
transform 1 0 28520 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_304
timestamp 1694700623
transform 1 0 29072 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_312
timestamp 1694700623
transform 1 0 29808 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_316
timestamp 1694700623
transform 1 0 30176 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_328
timestamp 1694700623
transform 1 0 31280 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1694700623
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1694700623
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 1694700623
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 1694700623
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 1694700623
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1694700623
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1694700623
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_405
timestamp 1694700623
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1694700623
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1694700623
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1694700623
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1694700623
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1694700623
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1694700623
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1694700623
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_77
timestamp 1694700623
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1694700623
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1694700623
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_99
timestamp 1694700623
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_103
timestamp 1694700623
transform 1 0 10580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_110
timestamp 1694700623
transform 1 0 11224 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1694700623
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_122
timestamp 1694700623
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_141
timestamp 1694700623
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_151
timestamp 1694700623
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_163
timestamp 1694700623
transform 1 0 16100 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_167
timestamp 1694700623
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_175
timestamp 1694700623
transform 1 0 17204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_187
timestamp 1694700623
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1694700623
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_197
timestamp 1694700623
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_205
timestamp 1694700623
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_217
timestamp 1694700623
transform 1 0 21068 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_229
timestamp 1694700623
transform 1 0 22172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_248
timestamp 1694700623
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_253
timestamp 1694700623
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_261
timestamp 1694700623
transform 1 0 25116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_282
timestamp 1694700623
transform 1 0 27048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1694700623
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1694700623
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_317
timestamp 1694700623
transform 1 0 30268 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_329
timestamp 1694700623
transform 1 0 31372 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_341
timestamp 1694700623
transform 1 0 32476 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_353
timestamp 1694700623
transform 1 0 33580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_361
timestamp 1694700623
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1694700623
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1694700623
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1694700623
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_401
timestamp 1694700623
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1694700623
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1694700623
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1694700623
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1694700623
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1694700623
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1694700623
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1694700623
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_69
timestamp 1694700623
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_107
timestamp 1694700623
transform 1 0 10948 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1694700623
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_119
timestamp 1694700623
transform 1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_126
timestamp 1694700623
transform 1 0 12696 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_132
timestamp 1694700623
transform 1 0 13248 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_136
timestamp 1694700623
transform 1 0 13616 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_151
timestamp 1694700623
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_163
timestamp 1694700623
transform 1 0 16100 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1694700623
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_180
timestamp 1694700623
transform 1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_188
timestamp 1694700623
transform 1 0 18400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_195
timestamp 1694700623
transform 1 0 19044 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_203
timestamp 1694700623
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_208
timestamp 1694700623
transform 1 0 20240 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_214
timestamp 1694700623
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1694700623
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1694700623
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_237
timestamp 1694700623
transform 1 0 22908 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_259
timestamp 1694700623
transform 1 0 24932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_293
timestamp 1694700623
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_299
timestamp 1694700623
transform 1 0 28612 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_307
timestamp 1694700623
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_319
timestamp 1694700623
transform 1 0 30452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_334
timestamp 1694700623
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_367
timestamp 1694700623
transform 1 0 34868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_379
timestamp 1694700623
transform 1 0 35972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1694700623
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1694700623
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_405
timestamp 1694700623
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1694700623
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1694700623
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1694700623
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1694700623
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1694700623
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1694700623
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1694700623
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1694700623
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1694700623
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1694700623
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_126
timestamp 1694700623
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_148
timestamp 1694700623
transform 1 0 14720 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_156
timestamp 1694700623
transform 1 0 15456 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_179
timestamp 1694700623
transform 1 0 17572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1694700623
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_197
timestamp 1694700623
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_214
timestamp 1694700623
transform 1 0 20792 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_222
timestamp 1694700623
transform 1 0 21528 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_232
timestamp 1694700623
transform 1 0 22448 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_246
timestamp 1694700623
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_257
timestamp 1694700623
transform 1 0 24748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_269
timestamp 1694700623
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1694700623
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_288
timestamp 1694700623
transform 1 0 27600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_297
timestamp 1694700623
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_305
timestamp 1694700623
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_309
timestamp 1694700623
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_318
timestamp 1694700623
transform 1 0 30360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_333
timestamp 1694700623
transform 1 0 31740 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_339
timestamp 1694700623
transform 1 0 32292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1694700623
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1694700623
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1694700623
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1694700623
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1694700623
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_401
timestamp 1694700623
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1694700623
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1694700623
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1694700623
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1694700623
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1694700623
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1694700623
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1694700623
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1694700623
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_81
timestamp 1694700623
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_102
timestamp 1694700623
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1694700623
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_116
timestamp 1694700623
transform 1 0 11776 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_128
timestamp 1694700623
transform 1 0 12880 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_136
timestamp 1694700623
transform 1 0 13616 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1694700623
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1694700623
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1694700623
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1694700623
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_182
timestamp 1694700623
transform 1 0 17848 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_202
timestamp 1694700623
transform 1 0 19688 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_214
timestamp 1694700623
transform 1 0 20792 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_220
timestamp 1694700623
transform 1 0 21344 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_245
timestamp 1694700623
transform 1 0 23644 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_271
timestamp 1694700623
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1694700623
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_281
timestamp 1694700623
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_287
timestamp 1694700623
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_317
timestamp 1694700623
transform 1 0 30268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_327
timestamp 1694700623
transform 1 0 31188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1694700623
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_337
timestamp 1694700623
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_352
timestamp 1694700623
transform 1 0 33488 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_364
timestamp 1694700623
transform 1 0 34592 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_376
timestamp 1694700623
transform 1 0 35696 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_388
timestamp 1694700623
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1694700623
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_401
timestamp 1694700623
transform 1 0 37996 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1694700623
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1694700623
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1694700623
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1694700623
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1694700623
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1694700623
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1694700623
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1694700623
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1694700623
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp 1694700623
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 1694700623
transform 1 0 9292 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_93
timestamp 1694700623
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_107
timestamp 1694700623
transform 1 0 10948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_123
timestamp 1694700623
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_128
timestamp 1694700623
transform 1 0 12880 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_155
timestamp 1694700623
transform 1 0 15364 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_163
timestamp 1694700623
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_171
timestamp 1694700623
transform 1 0 16836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_183
timestamp 1694700623
transform 1 0 17940 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_189
timestamp 1694700623
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1694700623
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1694700623
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_210
timestamp 1694700623
transform 1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_219
timestamp 1694700623
transform 1 0 21252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_242
timestamp 1694700623
transform 1 0 23368 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1694700623
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1694700623
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_267
timestamp 1694700623
transform 1 0 25668 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_273
timestamp 1694700623
transform 1 0 26220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_297
timestamp 1694700623
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_302
timestamp 1694700623
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_316
timestamp 1694700623
transform 1 0 30176 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_326
timestamp 1694700623
transform 1 0 31096 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_338
timestamp 1694700623
transform 1 0 32200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_342
timestamp 1694700623
transform 1 0 32568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_355
timestamp 1694700623
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1694700623
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1694700623
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1694700623
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1694700623
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 1694700623
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1694700623
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1694700623
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1694700623
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1694700623
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1694700623
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1694700623
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1694700623
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_69
timestamp 1694700623
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_77
timestamp 1694700623
transform 1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_101
timestamp 1694700623
transform 1 0 10396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1694700623
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1694700623
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_134
timestamp 1694700623
transform 1 0 13432 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_146
timestamp 1694700623
transform 1 0 14536 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1694700623
transform 1 0 15088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_162
timestamp 1694700623
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_175
timestamp 1694700623
transform 1 0 17204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_188
timestamp 1694700623
transform 1 0 18400 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_197
timestamp 1694700623
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_220
timestamp 1694700623
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1694700623
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_237
timestamp 1694700623
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_248
timestamp 1694700623
transform 1 0 23920 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_256
timestamp 1694700623
transform 1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_265
timestamp 1694700623
transform 1 0 25484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_273
timestamp 1694700623
transform 1 0 26220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_281
timestamp 1694700623
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_291
timestamp 1694700623
transform 1 0 27876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_303
timestamp 1694700623
transform 1 0 28980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_332
timestamp 1694700623
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_337
timestamp 1694700623
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_362
timestamp 1694700623
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_374
timestamp 1694700623
transform 1 0 35512 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_386
timestamp 1694700623
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1694700623
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_405
timestamp 1694700623
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1694700623
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1694700623
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1694700623
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1694700623
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1694700623
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1694700623
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1694700623
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1694700623
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1694700623
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1694700623
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_97
timestamp 1694700623
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1694700623
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_115
timestamp 1694700623
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 1694700623
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 1694700623
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_167
timestamp 1694700623
transform 1 0 16468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_192
timestamp 1694700623
transform 1 0 18768 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_238
timestamp 1694700623
transform 1 0 23000 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1694700623
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_253
timestamp 1694700623
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1694700623
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_277
timestamp 1694700623
transform 1 0 26588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_288
timestamp 1694700623
transform 1 0 27600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_296
timestamp 1694700623
transform 1 0 28336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_304
timestamp 1694700623
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_309
timestamp 1694700623
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_315
timestamp 1694700623
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_319
timestamp 1694700623
transform 1 0 30452 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_325
timestamp 1694700623
transform 1 0 31004 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_337
timestamp 1694700623
transform 1 0 32108 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_349
timestamp 1694700623
transform 1 0 33212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_361
timestamp 1694700623
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1694700623
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1694700623
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1694700623
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_401
timestamp 1694700623
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1694700623
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1694700623
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1694700623
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1694700623
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1694700623
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1694700623
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1694700623
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1694700623
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1694700623
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_93
timestamp 1694700623
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1694700623
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1694700623
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp 1694700623
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_144
timestamp 1694700623
transform 1 0 14352 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_154
timestamp 1694700623
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_158
timestamp 1694700623
transform 1 0 15640 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1694700623
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_192
timestamp 1694700623
transform 1 0 18768 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_200
timestamp 1694700623
transform 1 0 19504 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_207
timestamp 1694700623
transform 1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_219
timestamp 1694700623
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1694700623
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_237
timestamp 1694700623
transform 1 0 22908 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_255
timestamp 1694700623
transform 1 0 24564 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_268
timestamp 1694700623
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_281
timestamp 1694700623
transform 1 0 26956 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_289
timestamp 1694700623
transform 1 0 27692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_301
timestamp 1694700623
transform 1 0 28796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_305
timestamp 1694700623
transform 1 0 29164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_326
timestamp 1694700623
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1694700623
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_337
timestamp 1694700623
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_349
timestamp 1694700623
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_362
timestamp 1694700623
transform 1 0 34408 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_374
timestamp 1694700623
transform 1 0 35512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_386
timestamp 1694700623
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1694700623
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_405
timestamp 1694700623
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1694700623
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1694700623
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1694700623
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1694700623
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1694700623
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1694700623
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1694700623
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1694700623
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1694700623
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_151
timestamp 1694700623
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_163
timestamp 1694700623
transform 1 0 16100 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_175
timestamp 1694700623
transform 1 0 17204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1694700623
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1694700623
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1694700623
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1694700623
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_233
timestamp 1694700623
transform 1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_242
timestamp 1694700623
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1694700623
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_253
timestamp 1694700623
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_262
timestamp 1694700623
transform 1 0 25208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_266
timestamp 1694700623
transform 1 0 25576 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_291
timestamp 1694700623
transform 1 0 27876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_303
timestamp 1694700623
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1694700623
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_314
timestamp 1694700623
transform 1 0 29992 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_324
timestamp 1694700623
transform 1 0 30912 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_328
timestamp 1694700623
transform 1 0 31280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_359
timestamp 1694700623
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1694700623
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1694700623
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1694700623
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1694700623
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_401
timestamp 1694700623
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1694700623
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1694700623
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1694700623
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1694700623
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1694700623
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1694700623
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1694700623
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1694700623
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_81
timestamp 1694700623
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_89
timestamp 1694700623
transform 1 0 9292 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1694700623
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1694700623
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1694700623
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_137
timestamp 1694700623
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1694700623
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1694700623
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1694700623
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1694700623
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_214
timestamp 1694700623
transform 1 0 20792 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1694700623
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_234
timestamp 1694700623
transform 1 0 22632 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_242
timestamp 1694700623
transform 1 0 23368 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_262
timestamp 1694700623
transform 1 0 25208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_276
timestamp 1694700623
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_287
timestamp 1694700623
transform 1 0 27508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_297
timestamp 1694700623
transform 1 0 28428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_307
timestamp 1694700623
transform 1 0 29348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_314
timestamp 1694700623
transform 1 0 29992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_320
timestamp 1694700623
transform 1 0 30544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1694700623
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_337
timestamp 1694700623
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_341
timestamp 1694700623
transform 1 0 32476 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1694700623
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1694700623
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1694700623
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1694700623
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1694700623
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1694700623
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_405
timestamp 1694700623
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1694700623
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1694700623
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1694700623
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1694700623
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_41
timestamp 1694700623
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_50
timestamp 1694700623
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_62
timestamp 1694700623
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_74
timestamp 1694700623
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1694700623
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_92
timestamp 1694700623
transform 1 0 9568 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_104
timestamp 1694700623
transform 1 0 10672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_112
timestamp 1694700623
transform 1 0 11408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_117
timestamp 1694700623
transform 1 0 11868 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1694700623
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1694700623
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1694700623
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 1694700623
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_154
timestamp 1694700623
transform 1 0 15272 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_160
timestamp 1694700623
transform 1 0 15824 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1694700623
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_197
timestamp 1694700623
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_203
timestamp 1694700623
transform 1 0 19780 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_208
timestamp 1694700623
transform 1 0 20240 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_237
timestamp 1694700623
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1694700623
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_253
timestamp 1694700623
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_261
timestamp 1694700623
transform 1 0 25116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_269
timestamp 1694700623
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_276
timestamp 1694700623
transform 1 0 26496 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_284
timestamp 1694700623
transform 1 0 27232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_306
timestamp 1694700623
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1694700623
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_320
timestamp 1694700623
transform 1 0 30544 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1694700623
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_345
timestamp 1694700623
transform 1 0 32844 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_350
timestamp 1694700623
transform 1 0 33304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_362
timestamp 1694700623
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1694700623
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1694700623
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1694700623
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_401
timestamp 1694700623
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1694700623
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_15
timestamp 1694700623
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_21
timestamp 1694700623
transform 1 0 3036 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_30
timestamp 1694700623
transform 1 0 3864 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_38
timestamp 1694700623
transform 1 0 4600 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_69
timestamp 1694700623
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_101
timestamp 1694700623
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1694700623
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_134
timestamp 1694700623
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_142
timestamp 1694700623
transform 1 0 14168 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_163
timestamp 1694700623
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1694700623
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_184
timestamp 1694700623
transform 1 0 18032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_196
timestamp 1694700623
transform 1 0 19136 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_231
timestamp 1694700623
transform 1 0 22356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_239
timestamp 1694700623
transform 1 0 23092 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_245
timestamp 1694700623
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_259
timestamp 1694700623
transform 1 0 24932 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_267
timestamp 1694700623
transform 1 0 25668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1694700623
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1694700623
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1694700623
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1694700623
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1694700623
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_329
timestamp 1694700623
transform 1 0 31372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_344
timestamp 1694700623
transform 1 0 32752 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_351
timestamp 1694700623
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_363
timestamp 1694700623
transform 1 0 34500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_375
timestamp 1694700623
transform 1 0 35604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_387
timestamp 1694700623
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1694700623
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1694700623
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_405
timestamp 1694700623
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1694700623
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_32
timestamp 1694700623
transform 1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1694700623
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1694700623
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_121
timestamp 1694700623
transform 1 0 12236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_125
timestamp 1694700623
transform 1 0 12604 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_160
timestamp 1694700623
transform 1 0 15824 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_182
timestamp 1694700623
transform 1 0 17848 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1694700623
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1694700623
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_209
timestamp 1694700623
transform 1 0 20332 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_218
timestamp 1694700623
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_226
timestamp 1694700623
transform 1 0 21896 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_231
timestamp 1694700623
transform 1 0 22356 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_239
timestamp 1694700623
transform 1 0 23092 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_249
timestamp 1694700623
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1694700623
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_265
timestamp 1694700623
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_276
timestamp 1694700623
transform 1 0 26496 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_288
timestamp 1694700623
transform 1 0 27600 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_296
timestamp 1694700623
transform 1 0 28336 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1694700623
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_324
timestamp 1694700623
transform 1 0 30912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_332
timestamp 1694700623
transform 1 0 31648 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_337
timestamp 1694700623
transform 1 0 32108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_345
timestamp 1694700623
transform 1 0 32844 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1694700623
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1694700623
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1694700623
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1694700623
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1694700623
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_401
timestamp 1694700623
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1694700623
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_15
timestamp 1694700623
transform 1 0 2484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_40
timestamp 1694700623
transform 1 0 4784 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1694700623
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_60
timestamp 1694700623
transform 1 0 6624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_89
timestamp 1694700623
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_106
timestamp 1694700623
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_133
timestamp 1694700623
transform 1 0 13340 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_154
timestamp 1694700623
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1694700623
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1694700623
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_177
timestamp 1694700623
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_218
timestamp 1694700623
transform 1 0 21160 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_231
timestamp 1694700623
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_251
timestamp 1694700623
transform 1 0 24196 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_284
timestamp 1694700623
transform 1 0 27232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_288
timestamp 1694700623
transform 1 0 27600 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_293
timestamp 1694700623
transform 1 0 28060 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_324
timestamp 1694700623
transform 1 0 30912 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_337
timestamp 1694700623
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_354
timestamp 1694700623
transform 1 0 33672 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_366
timestamp 1694700623
transform 1 0 34776 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_378
timestamp 1694700623
transform 1 0 35880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_390
timestamp 1694700623
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1694700623
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_405
timestamp 1694700623
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1694700623
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_15
timestamp 1694700623
transform 1 0 2484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_24
timestamp 1694700623
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_29
timestamp 1694700623
transform 1 0 3772 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_38
timestamp 1694700623
transform 1 0 4600 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_50
timestamp 1694700623
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_64
timestamp 1694700623
transform 1 0 6992 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_76
timestamp 1694700623
transform 1 0 8096 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1694700623
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1694700623
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_109
timestamp 1694700623
transform 1 0 11132 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_118
timestamp 1694700623
transform 1 0 11960 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1694700623
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1694700623
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_147
timestamp 1694700623
transform 1 0 14628 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_178
timestamp 1694700623
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_182
timestamp 1694700623
transform 1 0 17848 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_192
timestamp 1694700623
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 1694700623
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1694700623
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1694700623
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_253
timestamp 1694700623
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_259
timestamp 1694700623
transform 1 0 24932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_264
timestamp 1694700623
transform 1 0 25392 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_277
timestamp 1694700623
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1694700623
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1694700623
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_324
timestamp 1694700623
transform 1 0 30912 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_336
timestamp 1694700623
transform 1 0 32016 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_344
timestamp 1694700623
transform 1 0 32752 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_351
timestamp 1694700623
transform 1 0 33396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1694700623
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1694700623
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1694700623
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 1694700623
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_401
timestamp 1694700623
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_3
timestamp 1694700623
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_9
timestamp 1694700623
transform 1 0 1932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_13
timestamp 1694700623
transform 1 0 2300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_17
timestamp 1694700623
transform 1 0 2668 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_26
timestamp 1694700623
transform 1 0 3496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_52
timestamp 1694700623
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1694700623
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_69
timestamp 1694700623
transform 1 0 7452 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_77
timestamp 1694700623
transform 1 0 8188 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_95
timestamp 1694700623
transform 1 0 9844 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_107
timestamp 1694700623
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1694700623
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_113
timestamp 1694700623
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_117
timestamp 1694700623
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_124
timestamp 1694700623
transform 1 0 12512 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_138
timestamp 1694700623
transform 1 0 13800 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_159
timestamp 1694700623
transform 1 0 15732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_163
timestamp 1694700623
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1694700623
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_198
timestamp 1694700623
transform 1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_204
timestamp 1694700623
transform 1 0 19872 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_216
timestamp 1694700623
transform 1 0 20976 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1694700623
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_225
timestamp 1694700623
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_231
timestamp 1694700623
transform 1 0 22356 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1694700623
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_293
timestamp 1694700623
transform 1 0 28060 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_302
timestamp 1694700623
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_314
timestamp 1694700623
transform 1 0 29992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_318
timestamp 1694700623
transform 1 0 30360 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_325
timestamp 1694700623
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_333
timestamp 1694700623
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_337
timestamp 1694700623
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_360
timestamp 1694700623
transform 1 0 34224 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_372
timestamp 1694700623
transform 1 0 35328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_384
timestamp 1694700623
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 1694700623
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_405
timestamp 1694700623
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_3
timestamp 1694700623
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 1694700623
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_85
timestamp 1694700623
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_91
timestamp 1694700623
transform 1 0 9476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1694700623
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1694700623
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1694700623
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_165
timestamp 1694700623
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_173
timestamp 1694700623
transform 1 0 17020 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_205
timestamp 1694700623
transform 1 0 19964 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_217
timestamp 1694700623
transform 1 0 21068 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_222
timestamp 1694700623
transform 1 0 21528 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_230
timestamp 1694700623
transform 1 0 22264 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_240
timestamp 1694700623
transform 1 0 23184 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_273
timestamp 1694700623
transform 1 0 26220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_286
timestamp 1694700623
transform 1 0 27416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 1694700623
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_309
timestamp 1694700623
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_318
timestamp 1694700623
transform 1 0 30360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_354
timestamp 1694700623
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1694700623
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1694700623
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1694700623
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1694700623
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_401
timestamp 1694700623
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_19
timestamp 1694700623
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 1694700623
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1694700623
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_75
timestamp 1694700623
transform 1 0 8004 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1694700623
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_117
timestamp 1694700623
transform 1 0 11868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_129
timestamp 1694700623
transform 1 0 12972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_147
timestamp 1694700623
transform 1 0 14628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_158
timestamp 1694700623
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1694700623
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_169
timestamp 1694700623
transform 1 0 16652 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_177
timestamp 1694700623
transform 1 0 17388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_189
timestamp 1694700623
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_200
timestamp 1694700623
transform 1 0 19504 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_209
timestamp 1694700623
transform 1 0 20332 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1694700623
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_232
timestamp 1694700623
transform 1 0 22448 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_267
timestamp 1694700623
transform 1 0 25668 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_273
timestamp 1694700623
transform 1 0 26220 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 1694700623
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_281
timestamp 1694700623
transform 1 0 26956 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_302
timestamp 1694700623
transform 1 0 28888 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_319
timestamp 1694700623
transform 1 0 30452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_327
timestamp 1694700623
transform 1 0 31188 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_334
timestamp 1694700623
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_346
timestamp 1694700623
transform 1 0 32936 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_358
timestamp 1694700623
transform 1 0 34040 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_370
timestamp 1694700623
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_382
timestamp 1694700623
transform 1 0 36248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_390
timestamp 1694700623
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 1694700623
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_405
timestamp 1694700623
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_3
timestamp 1694700623
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_17
timestamp 1694700623
transform 1 0 2668 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_32
timestamp 1694700623
transform 1 0 4048 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_40
timestamp 1694700623
transform 1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_49
timestamp 1694700623
transform 1 0 5612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_61
timestamp 1694700623
transform 1 0 6716 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_69
timestamp 1694700623
transform 1 0 7452 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1694700623
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1694700623
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1694700623
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_103
timestamp 1694700623
transform 1 0 10580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_112
timestamp 1694700623
transform 1 0 11408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_121
timestamp 1694700623
transform 1 0 12236 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_129
timestamp 1694700623
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1694700623
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_141
timestamp 1694700623
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_164
timestamp 1694700623
transform 1 0 16192 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_168
timestamp 1694700623
transform 1 0 16560 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_180
timestamp 1694700623
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_192
timestamp 1694700623
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_197
timestamp 1694700623
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_221
timestamp 1694700623
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_243
timestamp 1694700623
transform 1 0 23460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1694700623
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_253
timestamp 1694700623
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_261
timestamp 1694700623
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_296
timestamp 1694700623
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_312
timestamp 1694700623
transform 1 0 29808 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_318
timestamp 1694700623
transform 1 0 30360 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_322
timestamp 1694700623
transform 1 0 30728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_334
timestamp 1694700623
transform 1 0 31832 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_346
timestamp 1694700623
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_358
timestamp 1694700623
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1694700623
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 1694700623
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 1694700623
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_401
timestamp 1694700623
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_3
timestamp 1694700623
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_22
timestamp 1694700623
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_34
timestamp 1694700623
transform 1 0 4232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_39
timestamp 1694700623
transform 1 0 4692 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_49
timestamp 1694700623
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1694700623
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_57
timestamp 1694700623
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_63
timestamp 1694700623
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1694700623
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_81
timestamp 1694700623
transform 1 0 8556 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_96
timestamp 1694700623
transform 1 0 9936 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_104
timestamp 1694700623
transform 1 0 10672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_126
timestamp 1694700623
transform 1 0 12696 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_139
timestamp 1694700623
transform 1 0 13892 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_151
timestamp 1694700623
transform 1 0 14996 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_169
timestamp 1694700623
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_186
timestamp 1694700623
transform 1 0 18216 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_190
timestamp 1694700623
transform 1 0 18584 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_214
timestamp 1694700623
transform 1 0 20792 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_218
timestamp 1694700623
transform 1 0 21160 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1694700623
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_232
timestamp 1694700623
transform 1 0 22448 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_266
timestamp 1694700623
transform 1 0 25576 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 1694700623
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1694700623
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_293
timestamp 1694700623
transform 1 0 28060 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_328
timestamp 1694700623
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1694700623
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1694700623
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1694700623
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1694700623
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1694700623
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1694700623
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1694700623
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_405
timestamp 1694700623
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_3
timestamp 1694700623
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_11
timestamp 1694700623
transform 1 0 2116 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_29
timestamp 1694700623
transform 1 0 3772 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_54
timestamp 1694700623
transform 1 0 6072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_58
timestamp 1694700623
transform 1 0 6440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_80
timestamp 1694700623
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_104
timestamp 1694700623
transform 1 0 10672 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_126
timestamp 1694700623
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1694700623
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1694700623
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_158
timestamp 1694700623
transform 1 0 15640 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_164
timestamp 1694700623
transform 1 0 16192 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_173
timestamp 1694700623
transform 1 0 17020 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_185
timestamp 1694700623
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1694700623
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_210
timestamp 1694700623
transform 1 0 20424 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_222
timestamp 1694700623
transform 1 0 21528 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_233
timestamp 1694700623
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1694700623
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1694700623
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1694700623
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1694700623
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1694700623
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_289
timestamp 1694700623
transform 1 0 27692 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_293
timestamp 1694700623
transform 1 0 28060 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_306
timestamp 1694700623
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1694700623
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1694700623
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1694700623
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1694700623
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1694700623
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1694700623
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 1694700623
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 1694700623
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 1694700623
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_401
timestamp 1694700623
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1694700623
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_15
timestamp 1694700623
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_23
timestamp 1694700623
transform 1 0 3220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_32
timestamp 1694700623
transform 1 0 4048 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_68
timestamp 1694700623
transform 1 0 7360 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_113
timestamp 1694700623
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_130
timestamp 1694700623
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_147
timestamp 1694700623
transform 1 0 14628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_164
timestamp 1694700623
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_181
timestamp 1694700623
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_198
timestamp 1694700623
transform 1 0 19320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_206
timestamp 1694700623
transform 1 0 20056 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_218
timestamp 1694700623
transform 1 0 21160 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_222
timestamp 1694700623
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_241
timestamp 1694700623
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_253
timestamp 1694700623
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_265
timestamp 1694700623
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_277
timestamp 1694700623
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1694700623
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1694700623
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1694700623
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1694700623
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1694700623
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1694700623
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1694700623
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1694700623
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1694700623
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 1694700623
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 1694700623
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 1694700623
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1694700623
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_405
timestamp 1694700623
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1694700623
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1694700623
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1694700623
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_58
timestamp 1694700623
transform 1 0 6440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_66
timestamp 1694700623
transform 1 0 7176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_71
timestamp 1694700623
transform 1 0 7636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_80
timestamp 1694700623
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_109
timestamp 1694700623
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_117
timestamp 1694700623
transform 1 0 11868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_148
timestamp 1694700623
transform 1 0 14720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_159
timestamp 1694700623
transform 1 0 15732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_167
timestamp 1694700623
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_176
timestamp 1694700623
transform 1 0 17296 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_184
timestamp 1694700623
transform 1 0 18032 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1694700623
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_203
timestamp 1694700623
transform 1 0 19780 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_207
timestamp 1694700623
transform 1 0 20148 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_228
timestamp 1694700623
transform 1 0 22080 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_250
timestamp 1694700623
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1694700623
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1694700623
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1694700623
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1694700623
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1694700623
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1694700623
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1694700623
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1694700623
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1694700623
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1694700623
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1694700623
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1694700623
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1694700623
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1694700623
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1694700623
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_401
timestamp 1694700623
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1694700623
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1694700623
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1694700623
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1694700623
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1694700623
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1694700623
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_66
timestamp 1694700623
transform 1 0 7176 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_74
timestamp 1694700623
transform 1 0 7912 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_82
timestamp 1694700623
transform 1 0 8648 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_102
timestamp 1694700623
transform 1 0 10488 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1694700623
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1694700623
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_125
timestamp 1694700623
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_135
timestamp 1694700623
transform 1 0 13524 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_143
timestamp 1694700623
transform 1 0 14260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_152
timestamp 1694700623
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_156
timestamp 1694700623
transform 1 0 15456 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1694700623
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_181
timestamp 1694700623
transform 1 0 17756 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_187
timestamp 1694700623
transform 1 0 18308 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_194
timestamp 1694700623
transform 1 0 18952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_204
timestamp 1694700623
transform 1 0 19872 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_210
timestamp 1694700623
transform 1 0 20424 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1694700623
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1694700623
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_225
timestamp 1694700623
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_241
timestamp 1694700623
transform 1 0 23276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_253
timestamp 1694700623
transform 1 0 24380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_265
timestamp 1694700623
transform 1 0 25484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_277
timestamp 1694700623
transform 1 0 26588 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1694700623
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1694700623
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1694700623
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1694700623
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1694700623
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1694700623
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1694700623
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1694700623
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1694700623
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1694700623
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1694700623
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1694700623
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 1694700623
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_405
timestamp 1694700623
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1694700623
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1694700623
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1694700623
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1694700623
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_41
timestamp 1694700623
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_73
timestamp 1694700623
transform 1 0 7820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_126
timestamp 1694700623
transform 1 0 12696 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_134
timestamp 1694700623
transform 1 0 13432 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1694700623
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_153
timestamp 1694700623
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_161
timestamp 1694700623
transform 1 0 15916 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_170
timestamp 1694700623
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_182
timestamp 1694700623
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1694700623
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_200
timestamp 1694700623
transform 1 0 19504 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_208
timestamp 1694700623
transform 1 0 20240 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_225
timestamp 1694700623
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_237
timestamp 1694700623
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1694700623
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1694700623
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1694700623
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1694700623
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1694700623
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1694700623
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1694700623
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1694700623
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1694700623
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1694700623
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1694700623
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1694700623
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1694700623
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1694700623
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 1694700623
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 1694700623
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_401
timestamp 1694700623
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1694700623
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1694700623
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1694700623
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_39
timestamp 1694700623
transform 1 0 4692 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_77
timestamp 1694700623
transform 1 0 8188 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_110
timestamp 1694700623
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_113
timestamp 1694700623
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_121
timestamp 1694700623
transform 1 0 12236 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_158
timestamp 1694700623
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1694700623
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_169
timestamp 1694700623
transform 1 0 16652 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_177
timestamp 1694700623
transform 1 0 17388 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_182
timestamp 1694700623
transform 1 0 17848 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_209
timestamp 1694700623
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1694700623
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1694700623
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1694700623
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1694700623
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1694700623
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1694700623
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1694700623
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1694700623
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1694700623
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1694700623
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1694700623
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1694700623
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1694700623
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1694700623
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1694700623
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1694700623
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1694700623
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1694700623
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1694700623
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 1694700623
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_405
timestamp 1694700623
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1694700623
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1694700623
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1694700623
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1694700623
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_41
timestamp 1694700623
transform 1 0 4876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1694700623
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_88
timestamp 1694700623
transform 1 0 9200 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_100
timestamp 1694700623
transform 1 0 10304 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_119
timestamp 1694700623
transform 1 0 12052 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_127
timestamp 1694700623
transform 1 0 12788 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_131
timestamp 1694700623
transform 1 0 13156 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_135
timestamp 1694700623
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1694700623
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_141
timestamp 1694700623
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_191
timestamp 1694700623
transform 1 0 18676 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1694700623
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_197
timestamp 1694700623
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_203
timestamp 1694700623
transform 1 0 19780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_213
timestamp 1694700623
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_230
timestamp 1694700623
transform 1 0 22264 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_242
timestamp 1694700623
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 1694700623
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1694700623
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1694700623
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1694700623
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1694700623
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1694700623
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1694700623
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1694700623
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1694700623
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1694700623
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1694700623
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1694700623
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1694700623
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1694700623
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1694700623
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1694700623
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_401
timestamp 1694700623
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1694700623
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1694700623
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1694700623
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1694700623
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1694700623
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1694700623
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_57
timestamp 1694700623
transform 1 0 6348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_67
timestamp 1694700623
transform 1 0 7268 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_85
timestamp 1694700623
transform 1 0 8924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_97
timestamp 1694700623
transform 1 0 10028 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 1694700623
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_125
timestamp 1694700623
transform 1 0 12604 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_144
timestamp 1694700623
transform 1 0 14352 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_156
timestamp 1694700623
transform 1 0 15456 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_160
timestamp 1694700623
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1694700623
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1694700623
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_193
timestamp 1694700623
transform 1 0 18860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_197
timestamp 1694700623
transform 1 0 19228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_214
timestamp 1694700623
transform 1 0 20792 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1694700623
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1694700623
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1694700623
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1694700623
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1694700623
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1694700623
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1694700623
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1694700623
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1694700623
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1694700623
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1694700623
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1694700623
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1694700623
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1694700623
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1694700623
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1694700623
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1694700623
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1694700623
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1694700623
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1694700623
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_405
timestamp 1694700623
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1694700623
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1694700623
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1694700623
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1694700623
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1694700623
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_53
timestamp 1694700623
transform 1 0 5980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_64
timestamp 1694700623
transform 1 0 6992 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_80
timestamp 1694700623
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1694700623
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_97
timestamp 1694700623
transform 1 0 10028 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_106
timestamp 1694700623
transform 1 0 10856 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_118
timestamp 1694700623
transform 1 0 11960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_129
timestamp 1694700623
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_137
timestamp 1694700623
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1694700623
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1694700623
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_165
timestamp 1694700623
transform 1 0 16284 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_171
timestamp 1694700623
transform 1 0 16836 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_180
timestamp 1694700623
transform 1 0 17664 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_192
timestamp 1694700623
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1694700623
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1694700623
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1694700623
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1694700623
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1694700623
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1694700623
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1694700623
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1694700623
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1694700623
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1694700623
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1694700623
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1694700623
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1694700623
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1694700623
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1694700623
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1694700623
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1694700623
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1694700623
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1694700623
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1694700623
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1694700623
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_401
timestamp 1694700623
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1694700623
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1694700623
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1694700623
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1694700623
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1694700623
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1694700623
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1694700623
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_69
timestamp 1694700623
transform 1 0 7452 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_78
timestamp 1694700623
transform 1 0 8280 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_90
timestamp 1694700623
transform 1 0 9384 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_102
timestamp 1694700623
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 1694700623
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1694700623
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1694700623
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1694700623
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1694700623
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1694700623
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1694700623
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1694700623
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1694700623
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1694700623
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1694700623
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1694700623
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1694700623
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1694700623
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1694700623
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1694700623
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1694700623
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1694700623
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1694700623
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1694700623
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1694700623
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1694700623
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1694700623
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1694700623
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1694700623
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1694700623
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1694700623
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1694700623
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1694700623
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 1694700623
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 1694700623
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 1694700623
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_405
timestamp 1694700623
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1694700623
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1694700623
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1694700623
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1694700623
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1694700623
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1694700623
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1694700623
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1694700623
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1694700623
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1694700623
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1694700623
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1694700623
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1694700623
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1694700623
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1694700623
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1694700623
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1694700623
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1694700623
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1694700623
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1694700623
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1694700623
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1694700623
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1694700623
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1694700623
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1694700623
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1694700623
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1694700623
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1694700623
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1694700623
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1694700623
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1694700623
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1694700623
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1694700623
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1694700623
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1694700623
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1694700623
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1694700623
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1694700623
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1694700623
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1694700623
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1694700623
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 1694700623
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_401
timestamp 1694700623
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1694700623
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1694700623
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1694700623
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1694700623
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1694700623
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1694700623
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1694700623
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1694700623
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1694700623
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1694700623
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1694700623
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1694700623
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1694700623
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1694700623
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1694700623
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1694700623
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1694700623
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1694700623
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1694700623
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1694700623
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1694700623
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1694700623
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1694700623
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1694700623
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1694700623
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1694700623
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1694700623
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1694700623
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1694700623
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1694700623
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1694700623
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1694700623
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1694700623
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1694700623
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1694700623
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1694700623
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1694700623
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1694700623
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1694700623
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1694700623
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1694700623
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1694700623
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1694700623
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_405
timestamp 1694700623
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1694700623
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1694700623
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1694700623
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1694700623
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1694700623
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1694700623
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1694700623
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1694700623
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1694700623
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1694700623
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1694700623
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1694700623
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1694700623
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1694700623
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1694700623
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1694700623
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1694700623
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1694700623
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1694700623
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1694700623
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1694700623
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1694700623
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1694700623
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1694700623
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1694700623
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1694700623
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1694700623
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1694700623
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1694700623
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1694700623
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1694700623
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1694700623
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1694700623
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1694700623
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1694700623
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1694700623
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1694700623
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1694700623
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1694700623
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1694700623
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1694700623
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1694700623
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_401
timestamp 1694700623
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1694700623
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1694700623
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1694700623
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1694700623
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1694700623
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1694700623
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1694700623
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1694700623
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1694700623
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1694700623
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1694700623
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1694700623
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1694700623
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1694700623
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1694700623
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1694700623
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1694700623
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1694700623
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1694700623
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1694700623
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1694700623
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1694700623
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1694700623
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1694700623
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1694700623
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1694700623
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1694700623
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1694700623
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1694700623
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1694700623
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1694700623
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1694700623
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1694700623
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1694700623
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1694700623
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1694700623
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1694700623
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1694700623
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1694700623
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1694700623
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1694700623
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1694700623
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1694700623
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_405
timestamp 1694700623
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1694700623
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1694700623
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1694700623
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1694700623
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1694700623
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1694700623
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1694700623
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1694700623
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1694700623
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1694700623
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1694700623
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1694700623
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1694700623
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1694700623
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1694700623
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1694700623
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1694700623
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1694700623
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1694700623
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1694700623
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1694700623
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1694700623
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1694700623
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1694700623
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1694700623
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1694700623
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1694700623
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1694700623
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1694700623
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1694700623
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1694700623
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1694700623
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1694700623
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1694700623
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1694700623
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1694700623
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1694700623
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1694700623
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1694700623
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1694700623
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1694700623
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1694700623
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_401
timestamp 1694700623
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1694700623
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1694700623
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1694700623
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1694700623
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1694700623
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1694700623
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1694700623
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1694700623
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1694700623
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1694700623
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1694700623
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1694700623
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1694700623
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1694700623
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1694700623
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1694700623
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1694700623
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1694700623
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1694700623
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1694700623
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1694700623
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1694700623
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1694700623
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1694700623
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1694700623
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1694700623
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1694700623
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1694700623
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1694700623
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1694700623
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1694700623
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1694700623
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1694700623
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1694700623
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1694700623
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1694700623
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1694700623
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1694700623
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1694700623
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1694700623
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1694700623
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1694700623
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1694700623
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_405
timestamp 1694700623
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1694700623
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1694700623
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1694700623
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1694700623
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1694700623
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1694700623
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1694700623
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1694700623
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1694700623
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1694700623
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1694700623
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1694700623
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1694700623
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1694700623
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1694700623
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1694700623
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1694700623
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1694700623
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1694700623
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1694700623
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1694700623
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1694700623
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1694700623
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1694700623
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1694700623
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1694700623
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1694700623
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1694700623
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1694700623
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1694700623
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1694700623
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1694700623
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1694700623
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1694700623
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1694700623
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1694700623
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1694700623
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1694700623
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1694700623
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1694700623
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1694700623
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1694700623
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_401
timestamp 1694700623
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1694700623
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1694700623
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1694700623
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1694700623
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1694700623
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1694700623
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1694700623
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1694700623
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1694700623
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1694700623
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1694700623
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1694700623
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1694700623
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1694700623
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1694700623
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1694700623
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1694700623
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1694700623
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1694700623
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1694700623
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1694700623
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1694700623
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1694700623
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1694700623
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1694700623
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1694700623
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1694700623
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1694700623
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1694700623
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1694700623
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1694700623
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1694700623
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1694700623
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1694700623
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1694700623
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1694700623
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1694700623
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1694700623
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1694700623
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1694700623
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1694700623
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1694700623
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1694700623
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_405
timestamp 1694700623
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1694700623
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1694700623
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1694700623
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1694700623
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1694700623
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1694700623
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1694700623
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1694700623
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1694700623
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1694700623
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1694700623
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1694700623
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1694700623
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1694700623
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1694700623
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1694700623
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1694700623
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1694700623
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1694700623
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1694700623
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1694700623
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1694700623
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1694700623
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1694700623
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1694700623
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1694700623
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1694700623
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1694700623
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1694700623
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1694700623
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1694700623
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1694700623
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1694700623
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1694700623
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1694700623
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1694700623
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1694700623
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1694700623
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1694700623
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1694700623
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1694700623
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1694700623
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_401
timestamp 1694700623
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1694700623
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1694700623
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1694700623
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1694700623
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1694700623
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1694700623
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1694700623
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1694700623
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1694700623
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1694700623
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1694700623
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1694700623
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1694700623
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1694700623
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1694700623
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1694700623
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1694700623
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1694700623
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1694700623
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1694700623
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1694700623
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1694700623
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1694700623
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1694700623
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1694700623
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1694700623
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1694700623
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1694700623
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1694700623
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1694700623
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1694700623
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1694700623
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1694700623
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1694700623
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1694700623
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1694700623
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1694700623
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1694700623
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1694700623
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1694700623
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1694700623
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1694700623
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1694700623
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_405
timestamp 1694700623
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1694700623
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1694700623
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1694700623
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1694700623
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1694700623
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 1694700623
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1694700623
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1694700623
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 1694700623
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1694700623
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1694700623
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 1694700623
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1694700623
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1694700623
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1694700623
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1694700623
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_153
timestamp 1694700623
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_163
timestamp 1694700623
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_167
timestamp 1694700623
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_169
timestamp 1694700623
transform 1 0 16652 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_177
timestamp 1694700623
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_184
timestamp 1694700623
transform 1 0 18032 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_197
timestamp 1694700623
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_205
timestamp 1694700623
transform 1 0 19964 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_217
timestamp 1694700623
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_223
timestamp 1694700623
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_225
timestamp 1694700623
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1694700623
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1694700623
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1694700623
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1694700623
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1694700623
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 1694700623
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 1694700623
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 1694700623
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 1694700623
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1694700623
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1694700623
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 1694700623
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1694700623
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1694700623
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 1694700623
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1694700623
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1694700623
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 1694700623
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1694700623
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_405
timestamp 1694700623
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 20884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1694700623
transform 1 0 16928 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1694700623
transform 1 0 3128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1694700623
transform 1 0 7452 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1694700623
transform 1 0 7544 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1694700623
transform 1 0 6256 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1694700623
transform -1 0 7452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1694700623
transform 1 0 9016 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1694700623
transform 1 0 9384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1694700623
transform -1 0 5888 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1694700623
transform -1 0 4416 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1694700623
transform -1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1694700623
transform 1 0 3312 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1694700623
transform -1 0 4600 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1694700623
transform -1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1694700623
transform -1 0 4876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1694700623
transform -1 0 5980 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1694700623
transform -1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1694700623
transform -1 0 8464 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1694700623
transform -1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1694700623
transform -1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1694700623
transform -1 0 6256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1694700623
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1694700623
transform -1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1694700623
transform -1 0 3496 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1694700623
transform 1 0 10028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1694700623
transform 1 0 10672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1694700623
transform 1 0 6532 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1694700623
transform 1 0 10120 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1694700623
transform -1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1694700623
transform 1 0 12236 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1694700623
transform 1 0 1932 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1694700623
transform -1 0 10672 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1694700623
transform -1 0 22540 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1694700623
transform -1 0 4600 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1694700623
transform -1 0 8188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1694700623
transform -1 0 11960 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1694700623
transform 1 0 6992 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1694700623
transform 1 0 8648 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1694700623
transform -1 0 14996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1694700623
transform 1 0 19412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1694700623
transform -1 0 19964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1694700623
transform -1 0 18216 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1694700623
transform -1 0 13800 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1694700623
transform -1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1694700623
transform -1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1694700623
transform -1 0 13708 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1694700623
transform -1 0 9660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1694700623
transform -1 0 10580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 38548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output2
timestamp 1694700623
transform 1 0 19412 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 1694700623
transform 1 0 17480 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1694700623
transform 1 0 15548 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1694700623
transform -1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1694700623
transform -1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1694700623
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1694700623
transform -1 0 22540 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 1694700623
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1694700623
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 1694700623
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1694700623
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 1694700623
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1694700623
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 1694700623
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1694700623
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 1694700623
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1694700623
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 1694700623
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1694700623
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 1694700623
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1694700623
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 1694700623
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1694700623
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 1694700623
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1694700623
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 1694700623
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1694700623
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 1694700623
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1694700623
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 1694700623
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1694700623
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 1694700623
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1694700623
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 1694700623
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1694700623
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 1694700623
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1694700623
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 1694700623
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1694700623
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 1694700623
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1694700623
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 1694700623
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1694700623
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 1694700623
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1694700623
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 1694700623
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1694700623
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 1694700623
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1694700623
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 1694700623
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1694700623
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 1694700623
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1694700623
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 1694700623
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1694700623
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 1694700623
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1694700623
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 1694700623
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1694700623
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 1694700623
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1694700623
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 1694700623
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1694700623
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 1694700623
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1694700623
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 1694700623
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1694700623
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 1694700623
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1694700623
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 1694700623
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1694700623
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 1694700623
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1694700623
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 1694700623
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1694700623
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 1694700623
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1694700623
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 1694700623
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1694700623
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 1694700623
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1694700623
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 1694700623
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1694700623
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 1694700623
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1694700623
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 1694700623
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1694700623
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 1694700623
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1694700623
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 1694700623
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1694700623
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 1694700623
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1694700623
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 1694700623
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1694700623
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 1694700623
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1694700623
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 1694700623
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1694700623
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 1694700623
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1694700623
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 1694700623
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1694700623
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 1694700623
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1694700623
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 1694700623
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1694700623
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 3312 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 1694700623
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 1694700623
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 1694700623
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 1694700623
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 1694700623
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 1694700623
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 1694700623
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 1694700623
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 1694700623
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 1694700623
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 1694700623
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 1694700623
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 1694700623
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 1694700623
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 1694700623
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_149
timestamp 1694700623
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_150
timestamp 1694700623
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 1694700623
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 1694700623
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 1694700623
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_156
timestamp 1694700623
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_157
timestamp 1694700623
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 1694700623
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 1694700623
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 1694700623
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_162
timestamp 1694700623
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_163
timestamp 1694700623
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_164
timestamp 1694700623
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 1694700623
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 1694700623
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_169
timestamp 1694700623
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_170
timestamp 1694700623
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_171
timestamp 1694700623
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 1694700623
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 1694700623
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_175
timestamp 1694700623
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_176
timestamp 1694700623
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_177
timestamp 1694700623
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_178
timestamp 1694700623
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 1694700623
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_182
timestamp 1694700623
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_183
timestamp 1694700623
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_184
timestamp 1694700623
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_185
timestamp 1694700623
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 1694700623
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_188
timestamp 1694700623
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_189
timestamp 1694700623
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_190
timestamp 1694700623
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_191
timestamp 1694700623
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_192
timestamp 1694700623
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_195
timestamp 1694700623
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_196
timestamp 1694700623
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_197
timestamp 1694700623
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_198
timestamp 1694700623
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_199
timestamp 1694700623
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_201
timestamp 1694700623
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_202
timestamp 1694700623
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_203
timestamp 1694700623
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_204
timestamp 1694700623
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_205
timestamp 1694700623
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_206
timestamp 1694700623
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_208
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_209
timestamp 1694700623
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_210
timestamp 1694700623
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_211
timestamp 1694700623
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_212
timestamp 1694700623
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_213
timestamp 1694700623
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_214
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_215
timestamp 1694700623
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_216
timestamp 1694700623
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_217
timestamp 1694700623
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_218
timestamp 1694700623
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_219
timestamp 1694700623
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_220
timestamp 1694700623
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_221
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_222
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_223
timestamp 1694700623
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_224
timestamp 1694700623
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_225
timestamp 1694700623
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_226
timestamp 1694700623
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_227
timestamp 1694700623
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_228
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_229
timestamp 1694700623
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_230
timestamp 1694700623
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_231
timestamp 1694700623
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_232
timestamp 1694700623
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_233
timestamp 1694700623
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_234
timestamp 1694700623
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_235
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_236
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_237
timestamp 1694700623
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_238
timestamp 1694700623
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_239
timestamp 1694700623
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_240
timestamp 1694700623
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_241
timestamp 1694700623
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_242
timestamp 1694700623
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_243
timestamp 1694700623
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_244
timestamp 1694700623
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_245
timestamp 1694700623
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_246
timestamp 1694700623
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_247
timestamp 1694700623
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_248
timestamp 1694700623
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_249
timestamp 1694700623
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_250
timestamp 1694700623
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_251
timestamp 1694700623
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_252
timestamp 1694700623
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_253
timestamp 1694700623
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_254
timestamp 1694700623
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_255
timestamp 1694700623
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_256
timestamp 1694700623
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_257
timestamp 1694700623
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_258
timestamp 1694700623
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_259
timestamp 1694700623
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_260
timestamp 1694700623
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_261
timestamp 1694700623
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_262
timestamp 1694700623
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_263
timestamp 1694700623
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_264
timestamp 1694700623
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_265
timestamp 1694700623
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_266
timestamp 1694700623
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_267
timestamp 1694700623
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_268
timestamp 1694700623
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_269
timestamp 1694700623
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_270
timestamp 1694700623
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_271
timestamp 1694700623
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_272
timestamp 1694700623
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_273
timestamp 1694700623
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_274
timestamp 1694700623
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_275
timestamp 1694700623
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_276
timestamp 1694700623
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_277
timestamp 1694700623
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_278
timestamp 1694700623
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_279
timestamp 1694700623
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_280
timestamp 1694700623
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_281
timestamp 1694700623
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_282
timestamp 1694700623
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_283
timestamp 1694700623
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_284
timestamp 1694700623
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_285
timestamp 1694700623
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_286
timestamp 1694700623
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_287
timestamp 1694700623
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_288
timestamp 1694700623
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_289
timestamp 1694700623
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_290
timestamp 1694700623
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_291
timestamp 1694700623
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_292
timestamp 1694700623
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_293
timestamp 1694700623
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_294
timestamp 1694700623
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_295
timestamp 1694700623
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_296
timestamp 1694700623
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_297
timestamp 1694700623
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_298
timestamp 1694700623
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_299
timestamp 1694700623
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_300
timestamp 1694700623
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_301
timestamp 1694700623
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_302
timestamp 1694700623
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_303
timestamp 1694700623
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_304
timestamp 1694700623
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_305
timestamp 1694700623
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_306
timestamp 1694700623
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_307
timestamp 1694700623
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_308
timestamp 1694700623
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_309
timestamp 1694700623
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_310
timestamp 1694700623
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_311
timestamp 1694700623
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_312
timestamp 1694700623
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_313
timestamp 1694700623
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_314
timestamp 1694700623
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_315
timestamp 1694700623
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_316
timestamp 1694700623
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_317
timestamp 1694700623
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_318
timestamp 1694700623
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_319
timestamp 1694700623
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_320
timestamp 1694700623
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_321
timestamp 1694700623
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_322
timestamp 1694700623
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_323
timestamp 1694700623
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_324
timestamp 1694700623
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_325
timestamp 1694700623
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_326
timestamp 1694700623
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_327
timestamp 1694700623
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_328
timestamp 1694700623
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_329
timestamp 1694700623
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_330
timestamp 1694700623
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_331
timestamp 1694700623
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_332
timestamp 1694700623
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_333
timestamp 1694700623
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_334
timestamp 1694700623
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_335
timestamp 1694700623
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_336
timestamp 1694700623
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_337
timestamp 1694700623
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_338
timestamp 1694700623
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_339
timestamp 1694700623
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_340
timestamp 1694700623
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_341
timestamp 1694700623
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_342
timestamp 1694700623
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_343
timestamp 1694700623
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_344
timestamp 1694700623
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_345
timestamp 1694700623
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_346
timestamp 1694700623
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_347
timestamp 1694700623
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_348
timestamp 1694700623
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_349
timestamp 1694700623
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_350
timestamp 1694700623
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_351
timestamp 1694700623
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_352
timestamp 1694700623
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_353
timestamp 1694700623
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_354
timestamp 1694700623
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_355
timestamp 1694700623
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_356
timestamp 1694700623
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_357
timestamp 1694700623
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_358
timestamp 1694700623
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_359
timestamp 1694700623
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_360
timestamp 1694700623
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_361
timestamp 1694700623
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_362
timestamp 1694700623
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_363
timestamp 1694700623
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_364
timestamp 1694700623
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_365
timestamp 1694700623
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_366
timestamp 1694700623
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_367
timestamp 1694700623
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_368
timestamp 1694700623
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_369
timestamp 1694700623
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_370
timestamp 1694700623
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_371
timestamp 1694700623
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_372
timestamp 1694700623
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_373
timestamp 1694700623
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_374
timestamp 1694700623
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_375
timestamp 1694700623
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_376
timestamp 1694700623
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_377
timestamp 1694700623
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_378
timestamp 1694700623
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_379
timestamp 1694700623
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_380
timestamp 1694700623
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_381
timestamp 1694700623
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_382
timestamp 1694700623
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_383
timestamp 1694700623
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_384
timestamp 1694700623
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_385
timestamp 1694700623
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_386
timestamp 1694700623
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_387
timestamp 1694700623
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_388
timestamp 1694700623
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_389
timestamp 1694700623
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_390
timestamp 1694700623
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_391
timestamp 1694700623
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_392
timestamp 1694700623
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_393
timestamp 1694700623
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_394
timestamp 1694700623
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_395
timestamp 1694700623
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_396
timestamp 1694700623
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_397
timestamp 1694700623
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_398
timestamp 1694700623
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_399
timestamp 1694700623
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_400
timestamp 1694700623
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_401
timestamp 1694700623
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_402
timestamp 1694700623
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_403
timestamp 1694700623
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_404
timestamp 1694700623
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_405
timestamp 1694700623
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_406
timestamp 1694700623
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_407
timestamp 1694700623
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_408
timestamp 1694700623
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_409
timestamp 1694700623
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_410
timestamp 1694700623
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_411
timestamp 1694700623
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_412
timestamp 1694700623
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_413
timestamp 1694700623
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_414
timestamp 1694700623
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_415
timestamp 1694700623
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_416
timestamp 1694700623
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_417
timestamp 1694700623
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_418
timestamp 1694700623
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_419
timestamp 1694700623
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_420
timestamp 1694700623
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_421
timestamp 1694700623
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_422
timestamp 1694700623
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_423
timestamp 1694700623
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_424
timestamp 1694700623
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_425
timestamp 1694700623
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_426
timestamp 1694700623
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_427
timestamp 1694700623
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_428
timestamp 1694700623
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_429
timestamp 1694700623
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_430
timestamp 1694700623
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_431
timestamp 1694700623
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_432
timestamp 1694700623
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_433
timestamp 1694700623
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_434
timestamp 1694700623
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_435
timestamp 1694700623
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_436
timestamp 1694700623
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_437
timestamp 1694700623
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_438
timestamp 1694700623
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_439
timestamp 1694700623
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_440
timestamp 1694700623
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_441
timestamp 1694700623
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_442
timestamp 1694700623
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_443
timestamp 1694700623
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_444
timestamp 1694700623
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_445
timestamp 1694700623
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_446
timestamp 1694700623
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_447
timestamp 1694700623
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_448
timestamp 1694700623
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_449
timestamp 1694700623
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_450
timestamp 1694700623
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_451
timestamp 1694700623
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_452
timestamp 1694700623
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_453
timestamp 1694700623
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_454
timestamp 1694700623
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_455
timestamp 1694700623
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_456
timestamp 1694700623
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_457
timestamp 1694700623
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_458
timestamp 1694700623
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_459
timestamp 1694700623
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_460
timestamp 1694700623
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_461
timestamp 1694700623
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_462
timestamp 1694700623
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_463
timestamp 1694700623
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_464
timestamp 1694700623
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_465
timestamp 1694700623
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_466
timestamp 1694700623
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_467
timestamp 1694700623
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_468
timestamp 1694700623
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_469
timestamp 1694700623
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_470
timestamp 1694700623
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_471
timestamp 1694700623
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_472
timestamp 1694700623
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_473
timestamp 1694700623
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_474
timestamp 1694700623
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_475
timestamp 1694700623
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_476
timestamp 1694700623
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_477
timestamp 1694700623
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_478
timestamp 1694700623
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_479
timestamp 1694700623
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_480
timestamp 1694700623
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_481
timestamp 1694700623
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_482
timestamp 1694700623
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_483
timestamp 1694700623
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_484
timestamp 1694700623
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_485
timestamp 1694700623
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_486
timestamp 1694700623
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_487
timestamp 1694700623
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_488
timestamp 1694700623
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_489
timestamp 1694700623
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_490
timestamp 1694700623
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_491
timestamp 1694700623
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_492
timestamp 1694700623
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_493
timestamp 1694700623
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_494
timestamp 1694700623
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_495
timestamp 1694700623
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_496
timestamp 1694700623
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_497
timestamp 1694700623
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_498
timestamp 1694700623
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_499
timestamp 1694700623
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_500
timestamp 1694700623
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_501
timestamp 1694700623
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_502
timestamp 1694700623
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_503
timestamp 1694700623
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_504
timestamp 1694700623
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_505
timestamp 1694700623
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_506
timestamp 1694700623
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_507
timestamp 1694700623
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_508
timestamp 1694700623
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_509
timestamp 1694700623
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_510
timestamp 1694700623
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_511
timestamp 1694700623
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_512
timestamp 1694700623
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_513
timestamp 1694700623
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_514
timestamp 1694700623
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_515
timestamp 1694700623
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_516
timestamp 1694700623
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_517
timestamp 1694700623
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_518
timestamp 1694700623
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_519
timestamp 1694700623
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_520
timestamp 1694700623
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_521
timestamp 1694700623
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_522
timestamp 1694700623
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_523
timestamp 1694700623
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_524
timestamp 1694700623
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_525
timestamp 1694700623
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_526
timestamp 1694700623
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_527
timestamp 1694700623
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_528
timestamp 1694700623
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_529
timestamp 1694700623
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_530
timestamp 1694700623
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_531
timestamp 1694700623
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_532
timestamp 1694700623
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_533
timestamp 1694700623
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_534
timestamp 1694700623
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_535
timestamp 1694700623
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_536
timestamp 1694700623
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_537
timestamp 1694700623
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_538
timestamp 1694700623
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_539
timestamp 1694700623
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_540
timestamp 1694700623
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_541
timestamp 1694700623
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_542
timestamp 1694700623
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_543
timestamp 1694700623
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_544
timestamp 1694700623
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_545
timestamp 1694700623
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_546
timestamp 1694700623
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_547
timestamp 1694700623
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_548
timestamp 1694700623
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_549
timestamp 1694700623
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_550
timestamp 1694700623
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_551
timestamp 1694700623
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_552
timestamp 1694700623
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_553
timestamp 1694700623
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_554
timestamp 1694700623
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_555
timestamp 1694700623
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_556
timestamp 1694700623
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_557
timestamp 1694700623
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_558
timestamp 1694700623
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_559
timestamp 1694700623
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_560
timestamp 1694700623
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_561
timestamp 1694700623
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_562
timestamp 1694700623
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_563
timestamp 1694700623
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_564
timestamp 1694700623
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_565
timestamp 1694700623
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_566
timestamp 1694700623
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_567
timestamp 1694700623
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_568
timestamp 1694700623
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_569
timestamp 1694700623
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_570
timestamp 1694700623
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_571
timestamp 1694700623
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_572
timestamp 1694700623
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_573
timestamp 1694700623
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_574
timestamp 1694700623
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_575
timestamp 1694700623
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_576
timestamp 1694700623
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_577
timestamp 1694700623
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_578
timestamp 1694700623
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_579
timestamp 1694700623
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_580
timestamp 1694700623
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_581
timestamp 1694700623
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_582
timestamp 1694700623
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_583
timestamp 1694700623
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_584
timestamp 1694700623
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_585
timestamp 1694700623
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_586
timestamp 1694700623
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_587
timestamp 1694700623
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_588
timestamp 1694700623
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_589
timestamp 1694700623
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_590
timestamp 1694700623
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_591
timestamp 1694700623
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_592
timestamp 1694700623
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_593
timestamp 1694700623
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_594
timestamp 1694700623
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_595
timestamp 1694700623
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_596
timestamp 1694700623
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_597
timestamp 1694700623
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_598
timestamp 1694700623
transform 1 0 37168 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6006 38872 6326 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 36642 38872 36962 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5346 38872 5666 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 35982 38872 36302 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 clock
port 2 nsew signal input
flabel metal2 s 19338 39200 19394 40000 0 FreeSans 224 90 0 0 ram_addr_o[0]
port 3 nsew signal tristate
flabel metal2 s 17406 39200 17462 40000 0 FreeSans 224 90 0 0 ram_addr_o[1]
port 4 nsew signal tristate
flabel metal2 s 15474 39200 15530 40000 0 FreeSans 224 90 0 0 ram_addr_o[2]
port 5 nsew signal tristate
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 ram_addr_o[3]
port 6 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 ram_addr_o[4]
port 7 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 ram_data_io[0]
port 8 nsew signal bidirectional
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 ram_data_io[10]
port 9 nsew signal bidirectional
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 ram_data_io[11]
port 10 nsew signal bidirectional
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 ram_data_io[12]
port 11 nsew signal bidirectional
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 ram_data_io[13]
port 12 nsew signal bidirectional
flabel metal3 s 39200 16328 40000 16448 0 FreeSans 480 0 0 0 ram_data_io[14]
port 13 nsew signal bidirectional
flabel metal3 s 39200 14288 40000 14408 0 FreeSans 480 0 0 0 ram_data_io[15]
port 14 nsew signal bidirectional
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 ram_data_io[16]
port 15 nsew signal bidirectional
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 ram_data_io[17]
port 16 nsew signal bidirectional
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 ram_data_io[18]
port 17 nsew signal bidirectional
flabel metal3 s 39200 10208 40000 10328 0 FreeSans 480 0 0 0 ram_data_io[19]
port 18 nsew signal bidirectional
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 ram_data_io[1]
port 19 nsew signal bidirectional
flabel metal3 s 39200 12248 40000 12368 0 FreeSans 480 0 0 0 ram_data_io[20]
port 20 nsew signal bidirectional
flabel metal3 s 39200 14968 40000 15088 0 FreeSans 480 0 0 0 ram_data_io[21]
port 21 nsew signal bidirectional
flabel metal3 s 39200 15648 40000 15768 0 FreeSans 480 0 0 0 ram_data_io[22]
port 22 nsew signal bidirectional
flabel metal3 s 39200 18368 40000 18488 0 FreeSans 480 0 0 0 ram_data_io[23]
port 23 nsew signal bidirectional
flabel metal3 s 39200 19728 40000 19848 0 FreeSans 480 0 0 0 ram_data_io[24]
port 24 nsew signal bidirectional
flabel metal3 s 39200 24488 40000 24608 0 FreeSans 480 0 0 0 ram_data_io[25]
port 25 nsew signal bidirectional
flabel metal3 s 39200 25848 40000 25968 0 FreeSans 480 0 0 0 ram_data_io[26]
port 26 nsew signal bidirectional
flabel metal3 s 39200 25168 40000 25288 0 FreeSans 480 0 0 0 ram_data_io[27]
port 27 nsew signal bidirectional
flabel metal3 s 39200 23128 40000 23248 0 FreeSans 480 0 0 0 ram_data_io[28]
port 28 nsew signal bidirectional
flabel metal3 s 39200 17688 40000 17808 0 FreeSans 480 0 0 0 ram_data_io[29]
port 29 nsew signal bidirectional
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 ram_data_io[2]
port 30 nsew signal bidirectional
flabel metal3 s 39200 19048 40000 19168 0 FreeSans 480 0 0 0 ram_data_io[30]
port 31 nsew signal bidirectional
flabel metal2 s 23202 39200 23258 40000 0 FreeSans 224 90 0 0 ram_data_io[31]
port 32 nsew signal bidirectional
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 ram_data_io[3]
port 33 nsew signal bidirectional
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 ram_data_io[4]
port 34 nsew signal bidirectional
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 ram_data_io[5]
port 35 nsew signal bidirectional
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 ram_data_io[6]
port 36 nsew signal bidirectional
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ram_data_io[7]
port 37 nsew signal bidirectional
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 ram_data_io[8]
port 38 nsew signal bidirectional
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 ram_data_io[9]
port 39 nsew signal bidirectional
flabel metal3 s 39200 8168 40000 8288 0 FreeSans 480 0 0 0 ram_rw_en_o
port 40 nsew signal tristate
flabel metal3 s 39200 17008 40000 17128 0 FreeSans 480 0 0 0 reset_i
port 41 nsew signal input
flabel metal2 s 21914 39200 21970 40000 0 FreeSans 224 90 0 0 stop_lamp_o
port 42 nsew signal tristate
rlabel metal1 19964 36992 19964 36992 0 VGND
rlabel metal1 19964 37536 19964 37536 0 VPWR
rlabel metal1 20552 28526 20552 28526 0 _0000_
rlabel metal1 19267 18666 19267 18666 0 _0001_
rlabel metal1 18025 20910 18025 20910 0 _0002_
rlabel metal2 12098 21352 12098 21352 0 _0003_
rlabel metal2 9890 19992 9890 19992 0 _0004_
rlabel metal1 9660 17850 9660 17850 0 _0005_
rlabel metal1 9483 16150 9483 16150 0 _0006_
rlabel metal2 8694 13736 8694 13736 0 _0007_
rlabel metal1 9384 11866 9384 11866 0 _0008_
rlabel metal1 10495 10030 10495 10030 0 _0009_
rlabel metal2 12650 8296 12650 8296 0 _0010_
rlabel metal1 17303 7786 17303 7786 0 _0011_
rlabel metal1 21167 8534 21167 8534 0 _0012_
rlabel metal2 16330 12002 16330 12002 0 _0013_
rlabel metal1 17441 16558 17441 16558 0 _0014_
rlabel metal2 23230 17340 23230 17340 0 _0015_
rlabel metal1 25261 15062 25261 15062 0 _0016_
rlabel metal2 22218 9826 22218 9826 0 _0017_
rlabel metal2 23598 8296 23598 8296 0 _0018_
rlabel metal1 27324 7514 27324 7514 0 _0019_
rlabel metal2 30130 8738 30130 8738 0 _0020_
rlabel metal1 30360 14246 30360 14246 0 _0021_
rlabel metal2 26450 15606 26450 15606 0 _0022_
rlabel metal2 28658 17374 28658 17374 0 _0023_
rlabel metal2 30866 18462 30866 18462 0 _0024_
rlabel metal1 30452 18938 30452 18938 0 _0025_
rlabel metal2 31694 24344 31694 24344 0 _0026_
rlabel metal1 30544 25466 30544 25466 0 _0027_
rlabel metal2 26450 25058 26450 25058 0 _0028_
rlabel metal1 25484 24582 25484 24582 0 _0029_
rlabel metal1 28067 17578 28067 17578 0 _0030_
rlabel metal1 22547 20842 22547 20842 0 _0031_
rlabel metal2 22310 22882 22310 22882 0 _0032_
rlabel metal1 19044 23698 19044 23698 0 _0033_
rlabel metal1 17119 23018 17119 23018 0 _0034_
rlabel metal2 14490 22814 14490 22814 0 _0035_
rlabel metal2 12466 22440 12466 22440 0 _0036_
rlabel metal2 12374 23970 12374 23970 0 _0037_
rlabel metal2 18630 22814 18630 22814 0 _0038_
rlabel metal1 21167 23018 21167 23018 0 _0039_
rlabel metal2 20010 20638 20010 20638 0 _0040_
rlabel metal1 21344 27098 21344 27098 0 _0041_
rlabel metal1 19458 28730 19458 28730 0 _0042_
rlabel metal1 17664 29274 17664 29274 0 _0043_
rlabel metal1 15817 29614 15817 29614 0 _0044_
rlabel metal1 11691 28458 11691 28458 0 _0045_
rlabel metal2 13386 29342 13386 29342 0 _0046_
rlabel metal1 20608 18054 20608 18054 0 _0047_
rlabel metal1 16974 20808 16974 20808 0 _0048_
rlabel metal2 11822 21284 11822 21284 0 _0049_
rlabel metal1 9292 19890 9292 19890 0 _0050_
rlabel metal1 8924 17850 8924 17850 0 _0051_
rlabel metal1 8234 15674 8234 15674 0 _0052_
rlabel metal1 8188 13974 8188 13974 0 _0053_
rlabel metal1 9016 12138 9016 12138 0 _0054_
rlabel metal1 9292 9690 9292 9690 0 _0055_
rlabel metal1 12098 8058 12098 8058 0 _0056_
rlabel metal1 15962 7514 15962 7514 0 _0057_
rlabel metal1 19872 8058 19872 8058 0 _0058_
rlabel metal2 15410 12308 15410 12308 0 _0059_
rlabel metal1 16192 16218 16192 16218 0 _0060_
rlabel metal1 21666 17272 21666 17272 0 _0061_
rlabel metal2 23598 14484 23598 14484 0 _0062_
rlabel metal1 21567 10234 21567 10234 0 _0063_
rlabel metal1 23046 8534 23046 8534 0 _0064_
rlabel metal1 26588 7922 26588 7922 0 _0065_
rlabel metal1 29762 9010 29762 9010 0 _0066_
rlabel metal1 29716 12954 29716 12954 0 _0067_
rlabel metal2 25898 15572 25898 15572 0 _0068_
rlabel metal1 28060 16762 28060 16762 0 _0069_
rlabel metal1 29946 18326 29946 18326 0 _0070_
rlabel metal1 29578 19448 29578 19448 0 _0071_
rlabel metal1 31096 24242 31096 24242 0 _0072_
rlabel metal2 29762 25636 29762 25636 0 _0073_
rlabel metal1 25852 24922 25852 24922 0 _0074_
rlabel metal2 24702 23970 24702 23970 0 _0075_
rlabel metal2 26634 17816 26634 17816 0 _0076_
rlabel metal1 21252 20570 21252 20570 0 _0077_
rlabel metal2 22126 22610 22126 22610 0 _0078_
rlabel metal1 18124 23290 18124 23290 0 _0079_
rlabel metal1 15732 23018 15732 23018 0 _0080_
rlabel metal1 13754 22712 13754 22712 0 _0081_
rlabel metal2 11822 22746 11822 22746 0 _0082_
rlabel metal2 11638 23970 11638 23970 0 _0083_
rlabel metal1 17894 22712 17894 22712 0 _0084_
rlabel metal1 19780 23154 19780 23154 0 _0085_
rlabel metal1 19412 20502 19412 20502 0 _0086_
rlabel metal1 12696 29818 12696 29818 0 _0087_
rlabel metal1 20516 27098 20516 27098 0 _0088_
rlabel metal2 22586 25670 22586 25670 0 _0089_
rlabel metal1 23996 25942 23996 25942 0 _0090_
rlabel metal1 23648 27438 23648 27438 0 _0091_
rlabel viali 10897 29614 10897 29614 0 _0092_
rlabel metal1 3649 21930 3649 21930 0 _0093_
rlabel via1 3629 22610 3629 22610 0 _0094_
rlabel metal2 5566 21284 5566 21284 0 _0095_
rlabel metal2 7314 22100 7314 22100 0 _0096_
rlabel via1 7585 21930 7585 21930 0 _0097_
rlabel metal1 9798 21114 9798 21114 0 _0098_
rlabel metal1 9706 22610 9706 22610 0 _0099_
rlabel metal2 7682 23970 7682 23970 0 _0100_
rlabel via1 9425 25194 9425 25194 0 _0101_
rlabel metal1 11009 24106 11009 24106 0 _0102_
rlabel metal1 4779 24854 4779 24854 0 _0103_
rlabel metal1 6956 24174 6956 24174 0 _0104_
rlabel metal1 3802 24106 3802 24106 0 _0105_
rlabel metal2 2070 23970 2070 23970 0 _0106_
rlabel metal2 1978 25092 1978 25092 0 _0107_
rlabel metal1 3772 25466 3772 25466 0 _0108_
rlabel metal1 4968 26010 4968 26010 0 _0109_
rlabel metal1 4876 26894 4876 26894 0 _0110_
rlabel metal1 6762 27914 6762 27914 0 _0111_
rlabel metal1 5990 29138 5990 29138 0 _0112_
rlabel metal1 6486 30226 6486 30226 0 _0113_
rlabel metal1 8514 30294 8514 30294 0 _0114_
rlabel metal1 9108 28594 9108 28594 0 _0115_
rlabel metal1 10630 27438 10630 27438 0 _0116_
rlabel metal1 10580 26758 10580 26758 0 _0117_
rlabel metal1 7033 26350 7033 26350 0 _0118_
rlabel metal2 18262 28832 18262 28832 0 _0119_
rlabel metal1 16836 29274 16836 29274 0 _0120_
rlabel metal1 14904 29274 14904 29274 0 _0121_
rlabel metal2 12098 28322 12098 28322 0 _0122_
rlabel metal1 12742 28730 12742 28730 0 _0123_
rlabel metal1 20930 26554 20930 26554 0 _0124_
rlabel metal1 19826 26282 19826 26282 0 _0125_
rlabel metal1 20332 27030 20332 27030 0 _0126_
rlabel metal1 20010 26010 20010 26010 0 _0127_
rlabel metal2 21298 25330 21298 25330 0 _0128_
rlabel metal1 19458 27472 19458 27472 0 _0129_
rlabel metal1 20194 28186 20194 28186 0 _0130_
rlabel metal1 18446 28458 18446 28458 0 _0131_
rlabel metal1 13662 18768 13662 18768 0 _0132_
rlabel metal1 14674 24922 14674 24922 0 _0133_
rlabel metal1 16836 18734 16836 18734 0 _0134_
rlabel metal1 17480 25874 17480 25874 0 _0135_
rlabel metal1 17941 26962 17941 26962 0 _0136_
rlabel metal1 17802 25704 17802 25704 0 _0137_
rlabel metal1 17618 25364 17618 25364 0 _0138_
rlabel metal1 16330 25772 16330 25772 0 _0139_
rlabel metal1 14766 25330 14766 25330 0 _0140_
rlabel metal1 15226 25126 15226 25126 0 _0141_
rlabel metal1 12558 25228 12558 25228 0 _0142_
rlabel metal1 11086 25908 11086 25908 0 _0143_
rlabel metal1 11362 25806 11362 25806 0 _0144_
rlabel metal1 12834 26996 12834 26996 0 _0145_
rlabel metal1 12374 26894 12374 26894 0 _0146_
rlabel metal1 12098 26758 12098 26758 0 _0147_
rlabel metal1 12926 25874 12926 25874 0 _0148_
rlabel metal1 12604 27098 12604 27098 0 _0149_
rlabel metal1 19780 27438 19780 27438 0 _0150_
rlabel metal1 13846 27030 13846 27030 0 _0151_
rlabel metal1 14214 27098 14214 27098 0 _0152_
rlabel metal2 17066 27183 17066 27183 0 _0153_
rlabel metal1 15042 26928 15042 26928 0 _0154_
rlabel metal1 15042 27948 15042 27948 0 _0155_
rlabel metal1 14996 27506 14996 27506 0 _0156_
rlabel metal1 14122 27608 14122 27608 0 _0157_
rlabel metal1 13708 25874 13708 25874 0 _0158_
rlabel metal1 18538 27472 18538 27472 0 _0159_
rlabel metal1 13018 27336 13018 27336 0 _0160_
rlabel metal1 12328 27438 12328 27438 0 _0161_
rlabel metal1 13064 27642 13064 27642 0 _0162_
rlabel metal1 12696 25330 12696 25330 0 _0163_
rlabel metal1 13156 25466 13156 25466 0 _0164_
rlabel metal1 13892 26010 13892 26010 0 _0165_
rlabel metal1 13294 27098 13294 27098 0 _0166_
rlabel metal1 13570 28118 13570 28118 0 _0167_
rlabel metal2 15410 27642 15410 27642 0 _0168_
rlabel metal1 16192 25262 16192 25262 0 _0169_
rlabel metal1 15456 25330 15456 25330 0 _0170_
rlabel metal1 15272 25466 15272 25466 0 _0171_
rlabel metal2 15226 26758 15226 26758 0 _0172_
rlabel metal1 15640 27098 15640 27098 0 _0173_
rlabel metal1 15088 27574 15088 27574 0 _0174_
rlabel metal1 16836 27370 16836 27370 0 _0175_
rlabel metal2 16882 26214 16882 26214 0 _0176_
rlabel metal1 17526 26928 17526 26928 0 _0177_
rlabel metal1 17181 26282 17181 26282 0 _0178_
rlabel metal1 16468 26554 16468 26554 0 _0179_
rlabel metal1 17204 27574 17204 27574 0 _0180_
rlabel metal1 19090 26962 19090 26962 0 _0181_
rlabel metal2 18446 27574 18446 27574 0 _0182_
rlabel metal1 18676 27370 18676 27370 0 _0183_
rlabel metal2 18354 27234 18354 27234 0 _0184_
rlabel metal2 18722 27846 18722 27846 0 _0185_
rlabel metal1 18768 28186 18768 28186 0 _0186_
rlabel metal2 21482 24718 21482 24718 0 _0187_
rlabel metal1 21298 25942 21298 25942 0 _0188_
rlabel metal1 21666 24174 21666 24174 0 _0189_
rlabel metal1 20194 21386 20194 21386 0 _0190_
rlabel metal1 19734 21012 19734 21012 0 _0191_
rlabel metal1 19550 22746 19550 22746 0 _0192_
rlabel metal1 18124 22202 18124 22202 0 _0193_
rlabel metal1 12926 23800 12926 23800 0 _0194_
rlabel metal1 12052 23086 12052 23086 0 _0195_
rlabel metal1 14168 23698 14168 23698 0 _0196_
rlabel metal1 16376 23698 16376 23698 0 _0197_
rlabel metal1 18354 23086 18354 23086 0 _0198_
rlabel metal1 25208 18938 25208 18938 0 _0199_
rlabel metal1 23644 20434 23644 20434 0 _0200_
rlabel metal1 23414 20026 23414 20026 0 _0201_
rlabel metal2 24886 20196 24886 20196 0 _0202_
rlabel metal1 24656 20230 24656 20230 0 _0203_
rlabel metal1 25760 21114 25760 21114 0 _0204_
rlabel metal1 25392 18394 25392 18394 0 _0205_
rlabel metal1 25668 20434 25668 20434 0 _0206_
rlabel metal1 27462 20298 27462 20298 0 _0207_
rlabel metal1 27554 20978 27554 20978 0 _0208_
rlabel metal1 27830 20910 27830 20910 0 _0209_
rlabel metal1 26910 19856 26910 19856 0 _0210_
rlabel metal1 13570 13328 13570 13328 0 _0211_
rlabel viali 13479 13272 13479 13272 0 _0212_
rlabel metal1 14306 13940 14306 13940 0 _0213_
rlabel metal1 11454 15062 11454 15062 0 _0214_
rlabel metal2 11546 14722 11546 14722 0 _0215_
rlabel metal1 14122 14892 14122 14892 0 _0216_
rlabel metal2 12006 16762 12006 16762 0 _0217_
rlabel metal1 11914 16592 11914 16592 0 _0218_
rlabel metal1 12972 16558 12972 16558 0 _0219_
rlabel metal2 12558 17918 12558 17918 0 _0220_
rlabel metal1 14214 19312 14214 19312 0 _0221_
rlabel metal1 13294 17306 13294 17306 0 _0222_
rlabel metal1 13340 16490 13340 16490 0 _0223_
rlabel metal1 13892 15470 13892 15470 0 _0224_
rlabel metal1 13110 13226 13110 13226 0 _0225_
rlabel metal1 13984 13498 13984 13498 0 _0226_
rlabel metal1 14490 13430 14490 13430 0 _0227_
rlabel metal2 15226 14450 15226 14450 0 _0228_
rlabel metal2 14766 15300 14766 15300 0 _0229_
rlabel metal1 13261 20502 13261 20502 0 _0230_
rlabel metal1 13386 18632 13386 18632 0 _0231_
rlabel metal1 19228 18802 19228 18802 0 _0232_
rlabel metal1 16514 18394 16514 18394 0 _0233_
rlabel metal1 18078 18326 18078 18326 0 _0234_
rlabel metal1 18354 18938 18354 18938 0 _0235_
rlabel metal2 15410 19006 15410 19006 0 _0236_
rlabel metal1 15732 19278 15732 19278 0 _0237_
rlabel metal1 13432 18938 13432 18938 0 _0238_
rlabel metal2 14766 20060 14766 20060 0 _0239_
rlabel metal1 15778 18190 15778 18190 0 _0240_
rlabel metal1 14444 18734 14444 18734 0 _0241_
rlabel metal1 14628 17170 14628 17170 0 _0242_
rlabel metal2 14306 17680 14306 17680 0 _0243_
rlabel metal2 13754 16184 13754 16184 0 _0244_
rlabel metal1 15042 14382 15042 14382 0 _0245_
rlabel metal1 19274 10030 19274 10030 0 _0246_
rlabel metal1 17664 8942 17664 8942 0 _0247_
rlabel metal1 17940 10642 17940 10642 0 _0248_
rlabel metal1 18078 8602 18078 8602 0 _0249_
rlabel metal1 17434 10030 17434 10030 0 _0250_
rlabel metal1 17066 10098 17066 10098 0 _0251_
rlabel metal1 17480 10234 17480 10234 0 _0252_
rlabel metal2 14306 9146 14306 9146 0 _0253_
rlabel metal1 13754 9962 13754 9962 0 _0254_
rlabel metal1 14674 10676 14674 10676 0 _0255_
rlabel metal1 13754 10540 13754 10540 0 _0256_
rlabel metal1 14076 10438 14076 10438 0 _0257_
rlabel metal2 12466 10914 12466 10914 0 _0258_
rlabel metal2 11730 10948 11730 10948 0 _0259_
rlabel metal1 11868 11050 11868 11050 0 _0260_
rlabel metal1 14260 10642 14260 10642 0 _0261_
rlabel metal1 14306 11220 14306 11220 0 _0262_
rlabel metal1 15594 14382 15594 14382 0 _0263_
rlabel metal1 20930 15504 20930 15504 0 _0264_
rlabel metal2 21574 14722 21574 14722 0 _0265_
rlabel metal1 19964 14450 19964 14450 0 _0266_
rlabel metal1 20148 16422 20148 16422 0 _0267_
rlabel metal1 19228 16558 19228 16558 0 _0268_
rlabel metal1 20470 16082 20470 16082 0 _0269_
rlabel metal1 19826 16082 19826 16082 0 _0270_
rlabel metal1 20148 15470 20148 15470 0 _0271_
rlabel metal1 16882 15470 16882 15470 0 _0272_
rlabel metal1 17112 14382 17112 14382 0 _0273_
rlabel metal2 17802 15130 17802 15130 0 _0274_
rlabel metal1 17618 13294 17618 13294 0 _0275_
rlabel metal1 18078 13328 18078 13328 0 _0276_
rlabel metal1 18262 14416 18262 14416 0 _0277_
rlabel metal1 19780 14314 19780 14314 0 _0278_
rlabel metal1 17940 14518 17940 14518 0 _0279_
rlabel metal1 19918 13906 19918 13906 0 _0280_
rlabel metal1 16054 10472 16054 10472 0 _0281_
rlabel metal1 17710 10676 17710 10676 0 _0282_
rlabel metal1 17526 10710 17526 10710 0 _0283_
rlabel metal1 19458 13872 19458 13872 0 _0284_
rlabel metal1 16744 14586 16744 14586 0 _0285_
rlabel metal2 18630 14722 18630 14722 0 _0286_
rlabel metal1 20286 14960 20286 14960 0 _0287_
rlabel metal1 20470 15028 20470 15028 0 _0288_
rlabel metal1 19642 13974 19642 13974 0 _0289_
rlabel metal1 20953 13770 20953 13770 0 _0290_
rlabel metal1 33166 16422 33166 16422 0 _0291_
rlabel metal1 32844 19346 32844 19346 0 _0292_
rlabel via1 33710 16422 33710 16422 0 _0293_
rlabel metal1 33028 15878 33028 15878 0 _0294_
rlabel metal1 32108 16082 32108 16082 0 _0295_
rlabel metal1 31924 16490 31924 16490 0 _0296_
rlabel metal1 29486 15470 29486 15470 0 _0297_
rlabel metal2 29026 15164 29026 15164 0 _0298_
rlabel metal2 29946 15164 29946 15164 0 _0299_
rlabel metal1 30130 15062 30130 15062 0 _0300_
rlabel metal2 30682 15198 30682 15198 0 _0301_
rlabel metal1 31050 16082 31050 16082 0 _0302_
rlabel metal1 28658 14994 28658 14994 0 _0303_
rlabel metal1 32108 14382 32108 14382 0 _0304_
rlabel metal1 32476 12818 32476 12818 0 _0305_
rlabel metal1 32384 13906 32384 13906 0 _0306_
rlabel metal1 32062 12410 32062 12410 0 _0307_
rlabel metal1 31878 12240 31878 12240 0 _0308_
rlabel metal1 29854 10982 29854 10982 0 _0309_
rlabel metal1 30866 10676 30866 10676 0 _0310_
rlabel metal1 31924 11594 31924 11594 0 _0311_
rlabel metal2 31878 13940 31878 13940 0 _0312_
rlabel metal1 28842 14382 28842 14382 0 _0313_
rlabel metal1 30682 10506 30682 10506 0 _0314_
rlabel metal2 29854 9690 29854 9690 0 _0315_
rlabel metal1 29670 10540 29670 10540 0 _0316_
rlabel metal2 28106 10744 28106 10744 0 _0317_
rlabel metal1 28106 8840 28106 8840 0 _0318_
rlabel metal1 27140 8874 27140 8874 0 _0319_
rlabel metal1 28014 9520 28014 9520 0 _0320_
rlabel metal1 28336 9146 28336 9146 0 _0321_
rlabel metal1 27876 10642 27876 10642 0 _0322_
rlabel metal1 28290 10778 28290 10778 0 _0323_
rlabel metal1 25162 11118 25162 11118 0 _0324_
rlabel metal1 25070 10642 25070 10642 0 _0325_
rlabel metal2 25898 11492 25898 11492 0 _0326_
rlabel metal1 24794 11254 24794 11254 0 _0327_
rlabel metal1 26174 12240 26174 12240 0 _0328_
rlabel metal1 25116 13294 25116 13294 0 _0329_
rlabel metal2 24794 13124 24794 13124 0 _0330_
rlabel metal1 24426 11152 24426 11152 0 _0331_
rlabel metal1 24564 13362 24564 13362 0 _0332_
rlabel metal1 25254 12784 25254 12784 0 _0333_
rlabel metal2 28014 12619 28014 12619 0 _0334_
rlabel metal1 28060 13498 28060 13498 0 _0335_
rlabel metal1 29624 19754 29624 19754 0 _0336_
rlabel metal1 32890 14314 32890 14314 0 _0337_
rlabel metal1 33074 14008 33074 14008 0 _0338_
rlabel metal1 31142 15368 31142 15368 0 _0339_
rlabel metal1 29762 19992 29762 19992 0 _0340_
rlabel metal1 25484 12886 25484 12886 0 _0341_
rlabel metal1 27140 10642 27140 10642 0 _0342_
rlabel metal1 28014 11152 28014 11152 0 _0343_
rlabel metal1 28520 13362 28520 13362 0 _0344_
rlabel metal1 29448 19686 29448 19686 0 _0345_
rlabel metal1 33258 21862 33258 21862 0 _0346_
rlabel metal1 32890 23562 32890 23562 0 _0347_
rlabel metal1 33534 23222 33534 23222 0 _0348_
rlabel metal1 33166 22100 33166 22100 0 _0349_
rlabel metal1 32844 21862 32844 21862 0 _0350_
rlabel metal1 32890 21590 32890 21590 0 _0351_
rlabel metal1 33350 21556 33350 21556 0 _0352_
rlabel metal1 32614 21522 32614 21522 0 _0353_
rlabel metal1 33626 19822 33626 19822 0 _0354_
rlabel metal1 33166 19380 33166 19380 0 _0355_
rlabel metal1 31878 19788 31878 19788 0 _0356_
rlabel metal1 32292 19482 32292 19482 0 _0357_
rlabel metal1 31809 19686 31809 19686 0 _0358_
rlabel metal1 30728 20910 30728 20910 0 _0359_
rlabel metal1 28716 24242 28716 24242 0 _0360_
rlabel metal1 28290 23732 28290 23732 0 _0361_
rlabel metal1 28796 23086 28796 23086 0 _0362_
rlabel metal2 28704 21998 28704 21998 0 _0363_
rlabel metal1 29348 23154 29348 23154 0 _0364_
rlabel metal1 30406 23698 30406 23698 0 _0365_
rlabel metal2 30682 23290 30682 23290 0 _0366_
rlabel metal1 30728 22610 30728 22610 0 _0367_
rlabel metal1 30866 22678 30866 22678 0 _0368_
rlabel metal1 30682 21998 30682 21998 0 _0369_
rlabel metal1 29440 21862 29440 21862 0 _0370_
rlabel metal1 28704 20570 28704 20570 0 _0371_
rlabel metal1 31602 21930 31602 21930 0 _0372_
rlabel metal2 29302 22039 29302 22039 0 _0373_
rlabel metal1 28106 20944 28106 20944 0 _0374_
rlabel metal1 27922 20502 27922 20502 0 _0375_
rlabel metal1 28474 20842 28474 20842 0 _0376_
rlabel metal2 28474 21012 28474 21012 0 _0377_
rlabel metal2 26358 20128 26358 20128 0 _0378_
rlabel metal1 25024 19822 25024 19822 0 _0379_
rlabel metal1 25714 19822 25714 19822 0 _0380_
rlabel metal2 24150 20128 24150 20128 0 _0381_
rlabel metal1 23736 22066 23736 22066 0 _0382_
rlabel metal1 24058 21522 24058 21522 0 _0383_
rlabel metal1 23694 21522 23694 21522 0 _0384_
rlabel metal1 21528 23766 21528 23766 0 _0385_
rlabel metal1 17710 14892 17710 14892 0 _0386_
rlabel metal1 23736 21318 23736 21318 0 _0387_
rlabel metal1 21022 21522 21022 21522 0 _0388_
rlabel metal2 21758 18122 21758 18122 0 _0389_
rlabel metal1 24150 19482 24150 19482 0 _0390_
rlabel metal1 15870 21590 15870 21590 0 _0391_
rlabel metal2 12466 12886 12466 12886 0 _0392_
rlabel metal1 12742 12784 12742 12784 0 _0393_
rlabel metal2 12926 13090 12926 13090 0 _0394_
rlabel metal1 14912 8806 14912 8806 0 _0395_
rlabel metal1 20516 11730 20516 11730 0 _0396_
rlabel metal1 21160 12206 21160 12206 0 _0397_
rlabel metal1 21528 12138 21528 12138 0 _0398_
rlabel metal1 26634 12954 26634 12954 0 _0399_
rlabel metal2 27554 12206 27554 12206 0 _0400_
rlabel metal1 27784 13838 27784 13838 0 _0401_
rlabel metal2 33074 17085 33074 17085 0 _0402_
rlabel metal1 32798 22644 32798 22644 0 _0403_
rlabel metal1 26680 22066 26680 22066 0 _0404_
rlabel metal1 26036 22202 26036 22202 0 _0405_
rlabel metal2 25898 19601 25898 19601 0 _0406_
rlabel metal1 23690 18088 23690 18088 0 _0407_
rlabel metal1 23322 18326 23322 18326 0 _0408_
rlabel metal1 23782 18394 23782 18394 0 _0409_
rlabel metal1 23092 21658 23092 21658 0 _0410_
rlabel metal1 21528 21862 21528 21862 0 _0411_
rlabel metal2 17618 19346 17618 19346 0 _0412_
rlabel metal1 21390 18666 21390 18666 0 _0413_
rlabel metal1 20286 19346 20286 19346 0 _0414_
rlabel metal1 22402 21998 22402 21998 0 _0415_
rlabel metal1 17250 9622 17250 9622 0 _0416_
rlabel metal1 25852 20570 25852 20570 0 _0417_
rlabel viali 24241 20456 24241 20456 0 _0418_
rlabel metal1 23736 18870 23736 18870 0 _0419_
rlabel metal1 23828 18938 23828 18938 0 _0420_
rlabel metal1 32522 17034 32522 17034 0 _0421_
rlabel metal1 23322 20570 23322 20570 0 _0422_
rlabel metal1 21712 20434 21712 20434 0 _0423_
rlabel metal2 19642 19516 19642 19516 0 _0424_
rlabel metal1 27140 19346 27140 19346 0 _0425_
rlabel metal1 27554 19278 27554 19278 0 _0426_
rlabel metal1 27462 18734 27462 18734 0 _0427_
rlabel metal2 26174 18530 26174 18530 0 _0428_
rlabel metal1 15042 16082 15042 16082 0 _0429_
rlabel metal1 27508 18394 27508 18394 0 _0430_
rlabel metal1 26956 18258 26956 18258 0 _0431_
rlabel metal1 26496 22406 26496 22406 0 _0432_
rlabel metal1 25576 22610 25576 22610 0 _0433_
rlabel metal1 27278 21114 27278 21114 0 _0434_
rlabel metal1 25990 22746 25990 22746 0 _0435_
rlabel metal1 24886 23732 24886 23732 0 _0436_
rlabel metal1 31050 19788 31050 19788 0 _0437_
rlabel metal2 30406 21488 30406 21488 0 _0438_
rlabel metal1 29210 22644 29210 22644 0 _0439_
rlabel metal1 28753 22746 28753 22746 0 _0440_
rlabel metal1 28336 22746 28336 22746 0 _0441_
rlabel metal1 27830 22678 27830 22678 0 _0442_
rlabel metal1 28106 22746 28106 22746 0 _0443_
rlabel metal1 28244 23290 28244 23290 0 _0444_
rlabel metal1 26404 24378 26404 24378 0 _0445_
rlabel metal1 30498 22202 30498 22202 0 _0446_
rlabel metal1 29854 22712 29854 22712 0 _0447_
rlabel metal2 30590 23800 30590 23800 0 _0448_
rlabel metal1 29624 24922 29624 24922 0 _0449_
rlabel metal1 32154 21522 32154 21522 0 _0450_
rlabel via1 31789 21658 31789 21658 0 _0451_
rlabel metal2 32154 21828 32154 21828 0 _0452_
rlabel metal1 33028 22474 33028 22474 0 _0453_
rlabel metal1 32338 22066 32338 22066 0 _0454_
rlabel metal1 32154 21862 32154 21862 0 _0455_
rlabel metal1 32154 24684 32154 24684 0 _0456_
rlabel metal1 31004 20026 31004 20026 0 _0457_
rlabel metal1 32614 20536 32614 20536 0 _0458_
rlabel metal2 30498 20026 30498 20026 0 _0459_
rlabel metal1 30038 20026 30038 20026 0 _0460_
rlabel metal1 28014 13260 28014 13260 0 _0461_
rlabel metal2 30866 13158 30866 13158 0 _0462_
rlabel metal1 31464 15402 31464 15402 0 _0463_
rlabel metal1 30958 16524 30958 16524 0 _0464_
rlabel viali 31142 17172 31142 17172 0 _0465_
rlabel metal1 30912 16762 30912 16762 0 _0466_
rlabel metal1 32982 17034 32982 17034 0 _0467_
rlabel metal1 30866 17068 30866 17068 0 _0468_
rlabel metal1 30774 17306 30774 17306 0 _0469_
rlabel metal1 30176 17102 30176 17102 0 _0470_
rlabel metal1 29946 17850 29946 17850 0 _0471_
rlabel metal1 29854 16490 29854 16490 0 _0472_
rlabel via1 30143 16558 30143 16558 0 _0473_
rlabel metal1 29762 16762 29762 16762 0 _0474_
rlabel metal1 28842 16558 28842 16558 0 _0475_
rlabel metal1 31234 13940 31234 13940 0 _0476_
rlabel metal1 31878 13838 31878 13838 0 _0477_
rlabel metal1 31234 13804 31234 13804 0 _0478_
rlabel metal2 20746 12308 20746 12308 0 _0479_
rlabel metal1 20930 11832 20930 11832 0 _0480_
rlabel metal1 27792 11798 27792 11798 0 _0481_
rlabel metal1 28336 12750 28336 12750 0 _0482_
rlabel metal1 27554 13702 27554 13702 0 _0483_
rlabel metal1 22540 14314 22540 14314 0 _0484_
rlabel metal2 27094 14212 27094 14212 0 _0485_
rlabel metal1 27324 14586 27324 14586 0 _0486_
rlabel metal1 26082 15028 26082 15028 0 _0487_
rlabel metal1 30544 12750 30544 12750 0 _0488_
rlabel metal2 29302 13430 29302 13430 0 _0489_
rlabel metal1 30268 12954 30268 12954 0 _0490_
rlabel metal1 29532 12818 29532 12818 0 _0491_
rlabel metal1 27462 10710 27462 10710 0 _0492_
rlabel metal2 27922 10200 27922 10200 0 _0493_
rlabel metal1 29026 10710 29026 10710 0 _0494_
rlabel metal2 28934 10438 28934 10438 0 _0495_
rlabel metal1 29394 11152 29394 11152 0 _0496_
rlabel metal1 28632 10744 28632 10744 0 _0497_
rlabel metal1 29670 9690 29670 9690 0 _0498_
rlabel metal1 29716 9554 29716 9554 0 _0499_
rlabel metal2 27370 10234 27370 10234 0 _0500_
rlabel metal1 25576 10438 25576 10438 0 _0501_
rlabel metal1 25990 10064 25990 10064 0 _0502_
rlabel metal1 26887 9962 26887 9962 0 _0503_
rlabel metal1 27324 8942 27324 8942 0 _0504_
rlabel metal1 26772 8466 26772 8466 0 _0505_
rlabel metal1 25438 12818 25438 12818 0 _0506_
rlabel metal2 25070 12444 25070 12444 0 _0507_
rlabel metal2 25346 11152 25346 11152 0 _0508_
rlabel metal2 25806 9860 25806 9860 0 _0509_
rlabel metal1 25714 9962 25714 9962 0 _0510_
rlabel metal1 24978 8942 24978 8942 0 _0511_
rlabel metal1 23920 8942 23920 8942 0 _0512_
rlabel metal1 23368 12206 23368 12206 0 _0513_
rlabel metal1 24794 12138 24794 12138 0 _0514_
rlabel metal1 22678 11220 22678 11220 0 _0515_
rlabel metal2 22310 10812 22310 10812 0 _0516_
rlabel metal1 17848 14246 17848 14246 0 _0517_
rlabel metal1 18906 14042 18906 14042 0 _0518_
rlabel metal1 20792 14926 20792 14926 0 _0519_
rlabel metal2 21298 14620 21298 14620 0 _0520_
rlabel metal1 22724 13906 22724 13906 0 _0521_
rlabel metal1 21344 13362 21344 13362 0 _0522_
rlabel metal1 22858 12954 22858 12954 0 _0523_
rlabel metal1 23230 13498 23230 13498 0 _0524_
rlabel metal1 23506 13838 23506 13838 0 _0525_
rlabel metal1 23368 13906 23368 13906 0 _0526_
rlabel metal1 22034 13464 22034 13464 0 _0527_
rlabel metal2 21114 14688 21114 14688 0 _0528_
rlabel metal2 22494 15504 22494 15504 0 _0529_
rlabel metal1 21574 16762 21574 16762 0 _0530_
rlabel metal2 17848 14382 17848 14382 0 _0531_
rlabel metal1 18032 14586 18032 14586 0 _0532_
rlabel metal1 17940 14994 17940 14994 0 _0533_
rlabel metal1 18262 14790 18262 14790 0 _0534_
rlabel metal1 21117 12954 21117 12954 0 _0535_
rlabel metal1 20286 14042 20286 14042 0 _0536_
rlabel metal1 18492 15130 18492 15130 0 _0537_
rlabel metal1 17250 16014 17250 16014 0 _0538_
rlabel metal1 16698 16082 16698 16082 0 _0539_
rlabel metal2 19642 11900 19642 11900 0 _0540_
rlabel metal1 19504 12682 19504 12682 0 _0541_
rlabel metal1 18262 11866 18262 11866 0 _0542_
rlabel metal1 16192 12818 16192 12818 0 _0543_
rlabel metal1 14628 11186 14628 11186 0 _0544_
rlabel metal1 15456 10642 15456 10642 0 _0545_
rlabel metal1 16514 10608 16514 10608 0 _0546_
rlabel metal1 17848 10574 17848 10574 0 _0547_
rlabel metal2 19918 9996 19918 9996 0 _0548_
rlabel metal1 16422 8976 16422 8976 0 _0549_
rlabel metal1 17940 9010 17940 9010 0 _0550_
rlabel metal1 19412 9146 19412 9146 0 _0551_
rlabel metal1 20010 8942 20010 8942 0 _0552_
rlabel metal1 20240 7854 20240 7854 0 _0553_
rlabel metal1 16836 8942 16836 8942 0 _0554_
rlabel metal1 16790 10030 16790 10030 0 _0555_
rlabel metal1 16284 10642 16284 10642 0 _0556_
rlabel metal1 16376 10030 16376 10030 0 _0557_
rlabel metal1 16928 8602 16928 8602 0 _0558_
rlabel metal1 16468 7378 16468 7378 0 _0559_
rlabel metal1 13892 11186 13892 11186 0 _0560_
rlabel metal1 14306 9554 14306 9554 0 _0561_
rlabel metal1 15594 8976 15594 8976 0 _0562_
rlabel metal2 15962 9316 15962 9316 0 _0563_
rlabel metal1 14122 8534 14122 8534 0 _0564_
rlabel viali 12450 7850 12450 7850 0 _0565_
rlabel metal1 12650 9690 12650 9690 0 _0566_
rlabel metal1 12926 10064 12926 10064 0 _0567_
rlabel metal2 12558 10370 12558 10370 0 _0568_
rlabel metal1 9660 9554 9660 9554 0 _0569_
rlabel metal1 13984 14926 13984 14926 0 _0570_
rlabel metal1 14536 13838 14536 13838 0 _0571_
rlabel metal1 13294 12852 13294 12852 0 _0572_
rlabel metal1 13984 12818 13984 12818 0 _0573_
rlabel metal2 12466 12517 12466 12517 0 _0574_
rlabel metal1 13386 12410 13386 12410 0 _0575_
rlabel metal1 13110 12920 13110 12920 0 _0576_
rlabel metal1 9154 12614 9154 12614 0 _0577_
rlabel metal1 12190 15334 12190 15334 0 _0578_
rlabel metal1 12742 14382 12742 14382 0 _0579_
rlabel metal1 13018 14416 13018 14416 0 _0580_
rlabel metal1 12535 14246 12535 14246 0 _0581_
rlabel metal1 8786 14382 8786 14382 0 _0582_
rlabel metal1 13938 16218 13938 16218 0 _0583_
rlabel metal1 14904 17306 14904 17306 0 _0584_
rlabel metal1 14444 16626 14444 16626 0 _0585_
rlabel metal1 14582 16116 14582 16116 0 _0586_
rlabel metal1 11684 15946 11684 15946 0 _0587_
rlabel metal1 14766 16048 14766 16048 0 _0588_
rlabel metal1 14398 16184 14398 16184 0 _0589_
rlabel metal1 8602 15572 8602 15572 0 _0590_
rlabel metal1 14306 17680 14306 17680 0 _0591_
rlabel metal1 14536 17646 14536 17646 0 _0592_
rlabel metal2 14122 16694 14122 16694 0 _0593_
rlabel metal1 9430 16762 9430 16762 0 _0594_
rlabel metal1 14536 19482 14536 19482 0 _0595_
rlabel metal1 14628 19890 14628 19890 0 _0596_
rlabel metal1 14628 20026 14628 20026 0 _0597_
rlabel metal1 15456 20910 15456 20910 0 _0598_
rlabel metal1 14950 21046 14950 21046 0 _0599_
rlabel metal1 14812 20366 14812 20366 0 _0600_
rlabel metal1 13064 19754 13064 19754 0 _0601_
rlabel metal2 12006 20162 12006 20162 0 _0602_
rlabel metal2 16330 19584 16330 19584 0 _0603_
rlabel metal1 15686 19482 15686 19482 0 _0604_
rlabel metal2 15410 20791 15410 20791 0 _0605_
rlabel via1 15883 19822 15883 19822 0 _0606_
rlabel metal1 14720 19958 14720 19958 0 _0607_
rlabel metal1 11914 20298 11914 20298 0 _0608_
rlabel metal1 17940 18666 17940 18666 0 _0609_
rlabel metal1 17848 18394 17848 18394 0 _0610_
rlabel metal1 17365 18666 17365 18666 0 _0611_
rlabel metal2 17986 19686 17986 19686 0 _0612_
rlabel metal1 16790 20570 16790 20570 0 _0613_
rlabel metal1 20562 18326 20562 18326 0 _0614_
rlabel metal1 20332 18258 20332 18258 0 _0615_
rlabel metal1 9752 26010 9752 26010 0 _0616_
rlabel metal1 7866 21454 7866 21454 0 _0617_
rlabel metal2 9706 23868 9706 23868 0 _0618_
rlabel metal1 9844 23834 9844 23834 0 _0619_
rlabel metal1 3450 24106 3450 24106 0 _0620_
rlabel metal2 3542 25670 3542 25670 0 _0621_
rlabel metal2 4094 25568 4094 25568 0 _0622_
rlabel metal1 6440 28050 6440 28050 0 _0623_
rlabel metal1 6026 29580 6026 29580 0 _0624_
rlabel metal1 8970 29580 8970 29580 0 _0625_
rlabel metal2 9246 27302 9246 27302 0 _0626_
rlabel metal1 11040 26962 11040 26962 0 _0627_
rlabel metal1 7590 27472 7590 27472 0 _0628_
rlabel metal1 8326 26554 8326 26554 0 _0629_
rlabel metal1 7590 25874 7590 25874 0 _0630_
rlabel metal1 23046 26214 23046 26214 0 _0631_
rlabel metal1 20390 25194 20390 25194 0 _0632_
rlabel metal2 20930 25670 20930 25670 0 _0633_
rlabel metal1 19918 29648 19918 29648 0 _0634_
rlabel metal1 23046 26996 23046 26996 0 _0635_
rlabel metal1 22402 25398 22402 25398 0 _0636_
rlabel metal2 22126 24990 22126 24990 0 _0637_
rlabel metal2 19090 24956 19090 24956 0 _0638_
rlabel metal2 21942 17697 21942 17697 0 _0639_
rlabel metal1 17986 21556 17986 21556 0 _0640_
rlabel metal1 17618 17170 17618 17170 0 _0641_
rlabel metal1 30222 18768 30222 18768 0 _0642_
rlabel metal1 20010 21012 20010 21012 0 _0643_
rlabel metal1 11822 30362 11822 30362 0 _0644_
rlabel metal1 22724 27642 22724 27642 0 _0645_
rlabel metal1 22586 28016 22586 28016 0 _0646_
rlabel metal1 10718 30362 10718 30362 0 _0647_
rlabel metal1 5980 22474 5980 22474 0 _0648_
rlabel metal1 5336 21114 5336 21114 0 _0649_
rlabel metal2 6394 22916 6394 22916 0 _0650_
rlabel metal1 8418 21318 8418 21318 0 _0651_
rlabel metal1 8234 21658 8234 21658 0 _0652_
rlabel metal2 8970 22644 8970 22644 0 _0653_
rlabel metal1 8096 23698 8096 23698 0 _0654_
rlabel metal1 8188 23494 8188 23494 0 _0655_
rlabel metal1 8372 25466 8372 25466 0 _0656_
rlabel metal2 10810 25092 10810 25092 0 _0657_
rlabel metal1 5796 24922 5796 24922 0 _0658_
rlabel metal1 5382 24378 5382 24378 0 _0659_
rlabel metal1 6992 24650 6992 24650 0 _0660_
rlabel metal2 3910 24276 3910 24276 0 _0661_
rlabel metal1 3082 24922 3082 24922 0 _0662_
rlabel metal1 3312 23698 3312 23698 0 _0663_
rlabel metal1 4416 26010 4416 26010 0 _0664_
rlabel metal1 5382 26860 5382 26860 0 _0665_
rlabel metal1 5520 25874 5520 25874 0 _0666_
rlabel metal1 6900 28186 6900 28186 0 _0667_
rlabel metal1 7222 28050 7222 28050 0 _0668_
rlabel metal1 5980 28730 5980 28730 0 _0669_
rlabel metal1 7452 30906 7452 30906 0 _0670_
rlabel metal1 8648 28526 8648 28526 0 _0671_
rlabel metal1 10396 26962 10396 26962 0 _0672_
rlabel metal1 10626 27098 10626 27098 0 _0673_
rlabel metal1 9798 26248 9798 26248 0 _0674_
rlabel metal1 7360 26962 7360 26962 0 _0675_
rlabel metal1 21022 19176 21022 19176 0 clknet_0_clock
rlabel metal1 7774 13974 7774 13974 0 clknet_3_0__leaf_clock
rlabel metal1 13524 19142 13524 19142 0 clknet_3_1__leaf_clock
rlabel metal1 4002 22066 4002 22066 0 clknet_3_2__leaf_clock
rlabel metal1 15548 29682 15548 29682 0 clknet_3_3__leaf_clock
rlabel metal1 21298 17102 21298 17102 0 clknet_3_4__leaf_clock
rlabel metal1 27002 15368 27002 15368 0 clknet_3_5__leaf_clock
rlabel metal1 16698 20876 16698 20876 0 clknet_3_6__leaf_clock
rlabel metal1 21206 20978 21206 20978 0 clknet_3_7__leaf_clock
rlabel metal3 2062 29988 2062 29988 0 clock
rlabel metal1 4462 21522 4462 21522 0 manchester_baby_instance.BASE_0.s_countReg\[0\]
rlabel metal1 4508 23630 4508 23630 0 manchester_baby_instance.BASE_0.s_countReg\[10\]
rlabel metal1 5980 24378 5980 24378 0 manchester_baby_instance.BASE_0.s_countReg\[11\]
rlabel metal1 5612 23698 5612 23698 0 manchester_baby_instance.BASE_0.s_countReg\[12\]
rlabel metal1 2668 24786 2668 24786 0 manchester_baby_instance.BASE_0.s_countReg\[13\]
rlabel metal1 1656 24786 1656 24786 0 manchester_baby_instance.BASE_0.s_countReg\[14\]
rlabel metal2 3358 26724 3358 26724 0 manchester_baby_instance.BASE_0.s_countReg\[15\]
rlabel metal1 6164 26962 6164 26962 0 manchester_baby_instance.BASE_0.s_countReg\[16\]
rlabel metal1 5520 27506 5520 27506 0 manchester_baby_instance.BASE_0.s_countReg\[17\]
rlabel metal1 7912 28730 7912 28730 0 manchester_baby_instance.BASE_0.s_countReg\[18\]
rlabel metal1 5336 29274 5336 29274 0 manchester_baby_instance.BASE_0.s_countReg\[19\]
rlabel metal1 4968 21114 4968 21114 0 manchester_baby_instance.BASE_0.s_countReg\[1\]
rlabel metal1 7176 29478 7176 29478 0 manchester_baby_instance.BASE_0.s_countReg\[20\]
rlabel metal2 7498 30532 7498 30532 0 manchester_baby_instance.BASE_0.s_countReg\[21\]
rlabel metal2 9706 29444 9706 29444 0 manchester_baby_instance.BASE_0.s_countReg\[22\]
rlabel metal1 10028 27302 10028 27302 0 manchester_baby_instance.BASE_0.s_countReg\[23\]
rlabel metal1 10534 26452 10534 26452 0 manchester_baby_instance.BASE_0.s_countReg\[24\]
rlabel metal1 8326 26282 8326 26282 0 manchester_baby_instance.BASE_0.s_countReg\[25\]
rlabel metal1 5934 21522 5934 21522 0 manchester_baby_instance.BASE_0.s_countReg\[2\]
rlabel metal1 6118 21590 6118 21590 0 manchester_baby_instance.BASE_0.s_countReg\[3\]
rlabel metal1 8694 21896 8694 21896 0 manchester_baby_instance.BASE_0.s_countReg\[4\]
rlabel metal1 9384 21862 9384 21862 0 manchester_baby_instance.BASE_0.s_countReg\[5\]
rlabel metal1 8786 21454 8786 21454 0 manchester_baby_instance.BASE_0.s_countReg\[6\]
rlabel metal1 10350 23698 10350 23698 0 manchester_baby_instance.BASE_0.s_countReg\[7\]
rlabel metal1 9844 25466 9844 25466 0 manchester_baby_instance.BASE_0.s_countReg\[8\]
rlabel metal1 9844 24378 9844 24378 0 manchester_baby_instance.BASE_0.s_countReg\[9\]
rlabel metal1 9614 25772 9614 25772 0 manchester_baby_instance.BASE_0.s_tickNext
rlabel metal1 11362 30226 11362 30226 0 manchester_baby_instance.BASE_0.s_tickReg
rlabel metal1 20838 30158 20838 30158 0 manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
rlabel metal2 12466 29988 12466 29988 0 manchester_baby_instance.BASE_1.s_counterValue
rlabel metal1 14306 30124 14306 30124 0 manchester_baby_instance.BASE_1.s_derivedClock
rlabel metal1 19412 29070 19412 29070 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
rlabel metal2 17066 29308 17066 29308 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
rlabel metal2 16514 28832 16514 28832 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
rlabel metal1 10994 26010 10994 26010 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
rlabel metal1 14490 29070 14490 29070 0 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
rlabel metal1 22402 24616 22402 24616 0 manchester_baby_instance.CIRCUIT_0.Acc.tick
rlabel metal1 22264 27914 22264 27914 0 manchester_baby_instance.CIRCUIT_0.GATES_13.input1
rlabel metal1 24012 27438 24012 27438 0 manchester_baby_instance.CIRCUIT_0.GATES_13.result
rlabel metal1 18998 24378 18998 24378 0 manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
rlabel metal1 18906 21998 18906 21998 0 manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
rlabel metal1 20884 25262 20884 25262 0 manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
rlabel metal1 20838 21862 20838 21862 0 manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
rlabel metal1 16974 23290 16974 23290 0 manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
rlabel metal1 15410 23698 15410 23698 0 manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
rlabel metal1 14122 23154 14122 23154 0 manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
rlabel metal1 13846 23698 13846 23698 0 manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
rlabel metal1 22172 25670 22172 25670 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
rlabel metal2 23322 26180 23322 26180 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
rlabel metal1 21965 26554 21965 26554 0 manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
rlabel metal1 19688 18258 19688 18258 0 manchester_baby_instance.ram_data_i_0
rlabel metal1 17434 21896 17434 21896 0 manchester_baby_instance.ram_data_i_1
rlabel metal1 17342 8874 17342 8874 0 manchester_baby_instance.ram_data_i_10
rlabel metal1 18492 8942 18492 8942 0 manchester_baby_instance.ram_data_i_11
rlabel metal1 20102 12172 20102 12172 0 manchester_baby_instance.ram_data_i_12
rlabel metal2 18906 19584 18906 19584 0 manchester_baby_instance.ram_data_i_13
rlabel metal1 20010 16558 20010 16558 0 manchester_baby_instance.ram_data_i_14
rlabel metal2 20194 21114 20194 21114 0 manchester_baby_instance.ram_data_i_15
rlabel metal1 25438 11662 25438 11662 0 manchester_baby_instance.ram_data_i_16
rlabel metal1 25806 11866 25806 11866 0 manchester_baby_instance.ram_data_i_17
rlabel metal1 27646 11832 27646 11832 0 manchester_baby_instance.ram_data_i_18
rlabel metal2 32154 10914 32154 10914 0 manchester_baby_instance.ram_data_i_19
rlabel metal1 15272 21862 15272 21862 0 manchester_baby_instance.ram_data_i_2
rlabel metal1 32338 11594 32338 11594 0 manchester_baby_instance.ram_data_i_20
rlabel metal1 28290 15062 28290 15062 0 manchester_baby_instance.ram_data_i_21
rlabel metal1 29578 17646 29578 17646 0 manchester_baby_instance.ram_data_i_22
rlabel metal1 33948 17850 33948 17850 0 manchester_baby_instance.ram_data_i_23
rlabel metal1 33672 20434 33672 20434 0 manchester_baby_instance.ram_data_i_24
rlabel metal1 32798 23494 32798 23494 0 manchester_baby_instance.ram_data_i_25
rlabel metal2 28382 24956 28382 24956 0 manchester_baby_instance.ram_data_i_26
rlabel metal1 27876 24922 27876 24922 0 manchester_baby_instance.ram_data_i_27
rlabel metal1 26496 21998 26496 21998 0 manchester_baby_instance.ram_data_i_28
rlabel metal1 24104 19278 24104 19278 0 manchester_baby_instance.ram_data_i_29
rlabel metal1 14398 20910 14398 20910 0 manchester_baby_instance.ram_data_i_3
rlabel metal2 22862 20094 22862 20094 0 manchester_baby_instance.ram_data_i_30
rlabel metal1 24380 22610 24380 22610 0 manchester_baby_instance.ram_data_i_31
rlabel metal1 13294 24106 13294 24106 0 manchester_baby_instance.ram_data_i_4
rlabel metal1 11132 16150 11132 16150 0 manchester_baby_instance.ram_data_i_5
rlabel metal1 11914 12716 11914 12716 0 manchester_baby_instance.ram_data_i_6
rlabel metal1 11822 12784 11822 12784 0 manchester_baby_instance.ram_data_i_7
rlabel metal1 14582 9044 14582 9044 0 manchester_baby_instance.ram_data_i_8
rlabel metal1 15410 9146 15410 9146 0 manchester_baby_instance.ram_data_i_9
rlabel metal2 19550 17918 19550 17918 0 manchester_baby_instance.ram_data_o_0
rlabel metal1 16928 18190 16928 18190 0 manchester_baby_instance.ram_data_o_1
rlabel metal1 17250 8058 17250 8058 0 manchester_baby_instance.ram_data_o_10
rlabel metal1 20470 10064 20470 10064 0 manchester_baby_instance.ram_data_o_11
rlabel metal1 17342 12818 17342 12818 0 manchester_baby_instance.ram_data_o_12
rlabel metal1 17986 16558 17986 16558 0 manchester_baby_instance.ram_data_o_13
rlabel metal2 22034 17102 22034 17102 0 manchester_baby_instance.ram_data_o_14
rlabel metal2 23782 14076 23782 14076 0 manchester_baby_instance.ram_data_o_15
rlabel metal1 22862 10234 22862 10234 0 manchester_baby_instance.ram_data_o_16
rlabel metal1 24518 8466 24518 8466 0 manchester_baby_instance.ram_data_o_17
rlabel metal1 28658 7854 28658 7854 0 manchester_baby_instance.ram_data_o_18
rlabel metal1 30360 9622 30360 9622 0 manchester_baby_instance.ram_data_o_19
rlabel metal1 12873 19822 12873 19822 0 manchester_baby_instance.ram_data_o_2
rlabel metal1 32338 12172 32338 12172 0 manchester_baby_instance.ram_data_o_20
rlabel metal1 27048 16082 27048 16082 0 manchester_baby_instance.ram_data_o_21
rlabel metal2 32982 16354 32982 16354 0 manchester_baby_instance.ram_data_o_22
rlabel metal1 31188 18054 31188 18054 0 manchester_baby_instance.ram_data_o_23
rlabel metal1 32292 19822 32292 19822 0 manchester_baby_instance.ram_data_o_24
rlabel metal1 33028 24174 33028 24174 0 manchester_baby_instance.ram_data_o_25
rlabel metal1 30682 24786 30682 24786 0 manchester_baby_instance.ram_data_o_26
rlabel metal1 27370 24378 27370 24378 0 manchester_baby_instance.ram_data_o_27
rlabel metal1 25714 20978 25714 20978 0 manchester_baby_instance.ram_data_o_28
rlabel metal1 27462 18190 27462 18190 0 manchester_baby_instance.ram_data_o_29
rlabel metal2 13754 19516 13754 19516 0 manchester_baby_instance.ram_data_o_3
rlabel metal1 22218 20366 22218 20366 0 manchester_baby_instance.ram_data_o_30
rlabel metal1 19642 27472 19642 27472 0 manchester_baby_instance.ram_data_o_31
rlabel metal1 10442 17646 10442 17646 0 manchester_baby_instance.ram_data_o_4
rlabel metal1 11178 16558 11178 16558 0 manchester_baby_instance.ram_data_o_5
rlabel metal1 9614 14042 9614 14042 0 manchester_baby_instance.ram_data_o_6
rlabel metal1 9936 11730 9936 11730 0 manchester_baby_instance.ram_data_o_7
rlabel metal1 10626 10234 10626 10234 0 manchester_baby_instance.ram_data_o_8
rlabel metal1 13294 8262 13294 8262 0 manchester_baby_instance.ram_data_o_9
rlabel metal1 35696 17306 35696 17306 0 net1
rlabel metal1 18078 12342 18078 12342 0 net10
rlabel metal1 18538 17170 18538 17170 0 net11
rlabel metal2 18998 18428 18998 18428 0 net12
rlabel via1 25530 14365 25530 14365 0 net13
rlabel metal1 24610 17782 24610 17782 0 net14
rlabel metal2 32798 20985 32798 20985 0 net15
rlabel metal2 18722 20791 18722 20791 0 net16
rlabel metal1 2852 22746 2852 22746 0 net17
rlabel metal1 21339 29614 21339 29614 0 net18
rlabel metal2 17618 30192 17618 30192 0 net19
rlabel metal2 19550 34451 19550 34451 0 net2
rlabel metal1 4462 21318 4462 21318 0 net20
rlabel metal1 7774 30770 7774 30770 0 net21
rlabel metal1 8234 30804 8234 30804 0 net22
rlabel metal1 7084 22950 7084 22950 0 net24
rlabel via1 6950 21998 6950 21998 0 net25
rlabel metal1 9752 23086 9752 23086 0 net27
rlabel via1 10078 21590 10078 21590 0 net28
rlabel metal1 4508 23766 4508 23766 0 net29
rlabel metal1 17480 37162 17480 37162 0 net3
rlabel metal1 3680 24174 3680 24174 0 net30
rlabel metal2 8970 28934 8970 28934 0 net33
rlabel metal1 4370 25874 4370 25874 0 net34
rlabel metal1 3956 25262 3956 25262 0 net35
rlabel metal1 5290 27030 5290 27030 0 net36
rlabel metal2 4186 27234 4186 27234 0 net37
rlabel metal1 5428 28526 5428 28526 0 net38
rlabel metal1 6348 29070 6348 29070 0 net39
rlabel metal2 15686 36521 15686 36521 0 net4
rlabel metal1 7406 27404 7406 27404 0 net40
rlabel metal1 8050 21556 8050 21556 0 net42
rlabel metal1 7728 22610 7728 22610 0 net43
rlabel metal1 5428 21658 5428 21658 0 net44
rlabel metal1 5888 20910 5888 20910 0 net45
rlabel metal2 4830 21794 4830 21794 0 net46
rlabel metal1 2530 23698 2530 23698 0 net48
rlabel metal2 10718 24174 10718 24174 0 net49
rlabel metal1 7314 24616 7314 24616 0 net5
rlabel metal1 11822 24820 11822 24820 0 net50
rlabel via1 7410 29614 7410 29614 0 net52
rlabel via1 10814 21998 10814 21998 0 net54
rlabel metal1 11546 30022 11546 30022 0 net55
rlabel metal2 12926 30124 12926 30124 0 net56
rlabel metal2 2806 25670 2806 25670 0 net58
rlabel metal1 9660 26350 9660 26350 0 net59
rlabel metal1 1886 25194 1886 25194 0 net6
rlabel metal1 20654 26860 20654 26860 0 net60
rlabel metal1 3450 23154 3450 23154 0 net61
rlabel metal2 7498 28390 7498 28390 0 net62
rlabel metal1 10810 30294 10810 30294 0 net63
rlabel metal1 7728 24786 7728 24786 0 net65
rlabel metal1 9384 25874 9384 25874 0 net67
rlabel metal1 13110 28560 13110 28560 0 net68
rlabel metal1 20286 18326 20286 18326 0 net69
rlabel metal1 22448 24174 22448 24174 0 net7
rlabel metal1 18906 23834 18906 23834 0 net70
rlabel metal1 17296 23698 17296 23698 0 net71
rlabel metal1 13202 23834 13202 23834 0 net72
rlabel metal1 14812 23698 14812 23698 0 net73
rlabel metal1 6164 26894 6164 26894 0 net74
rlabel metal1 12788 23018 12788 23018 0 net75
rlabel metal1 9200 27642 9200 27642 0 net76
rlabel metal1 9522 26486 9522 26486 0 net77
rlabel metal2 22034 27132 22034 27132 0 net8
rlabel metal1 12926 7820 12926 7820 0 net9
rlabel metal1 19504 37434 19504 37434 0 ram_addr_o[0]
rlabel metal1 17572 37434 17572 37434 0 ram_addr_o[1]
rlabel metal1 15640 37434 15640 37434 0 ram_addr_o[2]
rlabel metal3 912 24548 912 24548 0 ram_addr_o[3]
rlabel metal3 820 25228 820 25228 0 ram_addr_o[4]
rlabel metal2 4094 20519 4094 20519 0 ram_data_io[0]
rlabel metal1 18216 7174 18216 7174 0 ram_data_io[10]
rlabel metal1 21482 7718 21482 7718 0 ram_data_io[11]
rlabel metal1 18538 12206 18538 12206 0 ram_data_io[12]
rlabel metal1 19044 16694 19044 16694 0 ram_data_io[13]
rlabel metal1 23414 16524 23414 16524 0 ram_data_io[14]
rlabel metal1 32798 14382 32798 14382 0 ram_data_io[15]
rlabel metal2 23230 1761 23230 1761 0 ram_data_io[16]
rlabel metal1 25300 8330 25300 8330 0 ram_data_io[17]
rlabel metal1 29072 7718 29072 7718 0 ram_data_io[18]
rlabel metal1 34132 10642 34132 10642 0 ram_data_io[19]
rlabel metal1 16652 21998 16652 21998 0 ram_data_io[1]
rlabel metal1 33902 12172 33902 12172 0 ram_data_io[20]
rlabel metal2 35466 15351 35466 15351 0 ram_data_io[21]
rlabel metal1 35926 16082 35926 16082 0 ram_data_io[22]
rlabel metal1 34500 18258 34500 18258 0 ram_data_io[23]
rlabel metal1 33810 19720 33810 19720 0 ram_data_io[24]
rlabel metal1 34500 24378 34500 24378 0 ram_data_io[25]
rlabel metal2 35466 25959 35466 25959 0 ram_data_io[26]
rlabel metal2 35466 25313 35466 25313 0 ram_data_io[27]
rlabel metal2 35466 23239 35466 23239 0 ram_data_io[28]
rlabel metal1 25622 17748 25622 17748 0 ram_data_io[29]
rlabel metal2 4002 22355 4002 22355 0 ram_data_io[2]
rlabel metal2 35466 18989 35466 18989 0 ram_data_io[30]
rlabel metal2 23230 37551 23230 37551 0 ram_data_io[31]
rlabel metal1 6992 19482 6992 19482 0 ram_data_io[3]
rlabel metal2 9890 17952 9890 17952 0 ram_data_io[4]
rlabel metal1 5980 15334 5980 15334 0 ram_data_io[5]
rlabel metal1 6578 13430 6578 13430 0 ram_data_io[6]
rlabel metal1 6670 11594 6670 11594 0 ram_data_io[7]
rlabel metal1 10902 8942 10902 8942 0 ram_data_io[8]
rlabel metal1 14076 7718 14076 7718 0 ram_data_io[9]
rlabel metal2 38410 8279 38410 8279 0 ram_rw_en_o
rlabel metal1 38686 17170 38686 17170 0 reset_i
rlabel metal1 22034 37434 22034 37434 0 stop_lamp_o
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
