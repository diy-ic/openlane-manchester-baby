// This is the unpowered netlist.
module manchester_baby (clock,
    clock_o,
    ram_rw_en_o,
    reset_i,
    stop_lamp_o,
    ram_addr_o,
    ram_data_i,
    ram_data_o);
 input clock;
 output clock_o;
 output ram_rw_en_o;
 input reset_i;
 output stop_lamp_o;
 output [4:0] ram_addr_o;
 input [31:0] ram_data_i;
 output [31:0] ram_data_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire clknet_0_clock;
 wire clknet_2_0__leaf_clock;
 wire clknet_2_1__leaf_clock;
 wire clknet_2_2__leaf_clock;
 wire clknet_2_3__leaf_clock;
 wire \manchester_baby_instance.BASE_0.s_countReg[0] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[1] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[2] ;
 wire \manchester_baby_instance.BASE_0.s_tickNext ;
 wire \manchester_baby_instance.BASE_0.s_tickReg ;
 wire \manchester_baby_instance.BASE_1.s_bufferRegs[0] ;
 wire \manchester_baby_instance.BASE_1.s_counterValue ;
 wire \manchester_baby_instance.BASE_1.s_derivedClock ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.Acc.tick ;
 wire \manchester_baby_instance.CIRCUIT_0.GATES_13.result ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[13] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[14] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[15] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__decap_6 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_159 ();
 sky130_fd_sc_hd__inv_2 _0542_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ));
 sky130_fd_sc_hd__and3b_1 _0543_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _0544_ (.A(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .C(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__a31o_1 _0545_ (.A1(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A3(_0102_),
    .B1(net85),
    .X(_0096_));
 sky130_fd_sc_hd__and4b_1 _0546_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .D(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0103_));
 sky130_fd_sc_hd__buf_2 _0547_ (.A(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0548_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .A1(net7),
    .S(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_1 _0549_ (.A(_0105_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0550_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A1(net6),
    .S(_0104_),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0551_ (.A(_0106_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0552_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A1(net5),
    .S(_0104_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0553_ (.A(_0107_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0554_ (.A0(net105),
    .A1(net27),
    .S(_0104_),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0555_ (.A(_0108_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0556_ (.A0(net107),
    .A1(net26),
    .S(_0104_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0557_ (.A(_0109_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _0558_ (.A0(net103),
    .A1(net23),
    .S(_0104_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0559_ (.A(_0110_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0560_ (.A0(net106),
    .A1(net12),
    .S(_0104_),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0111_),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_2 _0562_ (.A(net1),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0563_ (.A0(net100),
    .A1(_0112_),
    .S(_0104_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0564_ (.A(_0113_),
    .X(_0087_));
 sky130_fd_sc_hd__and3b_1 _0565_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .B(_0101_),
    .C(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .X(_0114_));
 sky130_fd_sc_hd__buf_2 _0566_ (.A(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__and4bb_2 _0567_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .C(_0101_),
    .D(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0116_));
 sky130_fd_sc_hd__o21a_2 _0568_ (.A1(_0115_),
    .A2(_0116_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _0569_ (.A(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__or3b_1 _0570_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .C_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .X(_0119_));
 sky130_fd_sc_hd__or4b_1 _0571_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .C(_0119_),
    .D_N(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0120_));
 sky130_fd_sc_hd__or4_4 _0572_ (.A(net26),
    .B(net23),
    .C(net12),
    .D(net1),
    .X(_0121_));
 sky130_fd_sc_hd__or2_1 _0573_ (.A(net27),
    .B(net28),
    .X(_0122_));
 sky130_fd_sc_hd__or2_1 _0574_ (.A(net29),
    .B(net30),
    .X(_0123_));
 sky130_fd_sc_hd__or2_1 _0575_ (.A(net31),
    .B(net32),
    .X(_0124_));
 sky130_fd_sc_hd__or4_4 _0576_ (.A(_0121_),
    .B(_0122_),
    .C(_0123_),
    .D(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _0577_ (.A(net2),
    .B(net3),
    .X(_0126_));
 sky130_fd_sc_hd__or4_4 _0578_ (.A(net5),
    .B(net4),
    .C(_0125_),
    .D(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__or2_1 _0579_ (.A(net7),
    .B(net6),
    .X(_0128_));
 sky130_fd_sc_hd__or4_4 _0580_ (.A(net8),
    .B(net9),
    .C(_0127_),
    .D(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__or2_1 _0581_ (.A(net13),
    .B(net14),
    .X(_0130_));
 sky130_fd_sc_hd__or4_4 _0582_ (.A(net10),
    .B(net11),
    .C(_0129_),
    .D(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__or3_4 _0583_ (.A(net15),
    .B(net16),
    .C(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__or3_4 _0584_ (.A(net17),
    .B(net18),
    .C(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__or3_4 _0585_ (.A(net19),
    .B(net20),
    .C(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__or4_4 _0586_ (.A(net21),
    .B(net22),
    .C(net24),
    .D(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__xnor2_2 _0587_ (.A(net25),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__or2b_1 _0588_ (.A(net24),
    .B_N(net63),
    .X(_0137_));
 sky130_fd_sc_hd__or2b_1 _0589_ (.A(net21),
    .B_N(net60),
    .X(_0138_));
 sky130_fd_sc_hd__or2b_1 _0590_ (.A(net75),
    .B_N(net65),
    .X(_0139_));
 sky130_fd_sc_hd__or2b_1 _0591_ (.A(net23),
    .B_N(net62),
    .X(_0140_));
 sky130_fd_sc_hd__xnor2_1 _0592_ (.A(net23),
    .B(net62),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _0593_ (.A(net12),
    .B(net51),
    .Y(_0142_));
 sky130_fd_sc_hd__or2b_1 _0594_ (.A(net40),
    .B_N(_0112_),
    .X(_0143_));
 sky130_fd_sc_hd__and2b_1 _0595_ (.A_N(net12),
    .B(net51),
    .X(_0144_));
 sky130_fd_sc_hd__a21o_1 _0596_ (.A1(_0142_),
    .A2(_0143_),
    .B1(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_1 _0597_ (.A(_0141_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__and2b_1 _0598_ (.A_N(net67),
    .B(net28),
    .X(_0147_));
 sky130_fd_sc_hd__or2b_1 _0599_ (.A(net28),
    .B_N(net67),
    .X(_0148_));
 sky130_fd_sc_hd__or2b_1 _0600_ (.A(_0147_),
    .B_N(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__or2b_1 _0601_ (.A(net27),
    .B_N(net66),
    .X(_0150_));
 sky130_fd_sc_hd__or2b_1 _0602_ (.A(net66),
    .B_N(net27),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _0603_ (.A(_0150_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__or2_1 _0604_ (.A(_0149_),
    .B(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__and2b_1 _0605_ (.A_N(net65),
    .B(net75),
    .X(_0154_));
 sky130_fd_sc_hd__a311o_1 _0606_ (.A1(_0139_),
    .A2(_0140_),
    .A3(_0146_),
    .B1(_0153_),
    .C1(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(net29),
    .Y(_0156_));
 sky130_fd_sc_hd__or2b_1 _0608_ (.A(net69),
    .B_N(net30),
    .X(_0157_));
 sky130_fd_sc_hd__and2b_1 _0609_ (.A_N(net30),
    .B(net69),
    .X(_0158_));
 sky130_fd_sc_hd__a31o_1 _0610_ (.A1(net68),
    .A2(_0156_),
    .A3(_0157_),
    .B1(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__a21o_1 _0611_ (.A1(_0148_),
    .A2(_0150_),
    .B1(_0147_),
    .X(_0160_));
 sky130_fd_sc_hd__and2b_1 _0612_ (.A_N(_0159_),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__or2_1 _0613_ (.A(net68),
    .B(_0156_),
    .X(_0162_));
 sky130_fd_sc_hd__a21oi_1 _0614_ (.A1(_0157_),
    .A2(_0162_),
    .B1(_0158_),
    .Y(_0163_));
 sky130_fd_sc_hd__xor2_1 _0615_ (.A(net42),
    .B(net3),
    .X(_0164_));
 sky130_fd_sc_hd__xor2_1 _0616_ (.A(net41),
    .B(net2),
    .X(_0165_));
 sky130_fd_sc_hd__or2_1 _0617_ (.A(_0164_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__and2b_1 _0618_ (.A_N(net71),
    .B(net32),
    .X(_0167_));
 sky130_fd_sc_hd__or2b_1 _0619_ (.A(net32),
    .B_N(net71),
    .X(_0168_));
 sky130_fd_sc_hd__or2b_1 _0620_ (.A(_0167_),
    .B_N(_0168_),
    .X(_0169_));
 sky130_fd_sc_hd__or2b_1 _0621_ (.A(net31),
    .B_N(net70),
    .X(_0170_));
 sky130_fd_sc_hd__or2b_1 _0622_ (.A(net70),
    .B_N(net31),
    .X(_0171_));
 sky130_fd_sc_hd__nand2_1 _0623_ (.A(_0170_),
    .B(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__or3_1 _0624_ (.A(_0166_),
    .B(_0169_),
    .C(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__xor2_1 _0625_ (.A(net6),
    .B(net45),
    .X(_0174_));
 sky130_fd_sc_hd__xor2_1 _0626_ (.A(net7),
    .B(net46),
    .X(_0175_));
 sky130_fd_sc_hd__or2b_1 _0627_ (.A(net4),
    .B_N(net43),
    .X(_0176_));
 sky130_fd_sc_hd__or2b_1 _0628_ (.A(net43),
    .B_N(net4),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__and2b_1 _0630_ (.A_N(net5),
    .B(net44),
    .X(_0179_));
 sky130_fd_sc_hd__and2b_1 _0631_ (.A_N(net44),
    .B(net5),
    .X(_0180_));
 sky130_fd_sc_hd__or2_1 _0632_ (.A(_0179_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__or4_1 _0633_ (.A(_0174_),
    .B(_0175_),
    .C(_0178_),
    .D(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__or2_1 _0634_ (.A(_0173_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a211o_1 _0635_ (.A1(_0155_),
    .A2(_0161_),
    .B1(_0163_),
    .C1(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__inv_2 _0636_ (.A(net42),
    .Y(_0185_));
 sky130_fd_sc_hd__a21o_1 _0637_ (.A1(_0168_),
    .A2(_0170_),
    .B1(_0167_),
    .X(_0186_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(net41),
    .Y(_0187_));
 sky130_fd_sc_hd__a211o_1 _0639_ (.A1(_0185_),
    .A2(net3),
    .B1(net2),
    .C1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__o221a_1 _0640_ (.A1(_0185_),
    .A2(net3),
    .B1(_0166_),
    .B2(_0186_),
    .C1(_0188_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(net44),
    .Y(_0190_));
 sky130_fd_sc_hd__o21a_1 _0642_ (.A1(net5),
    .A2(_0190_),
    .B1(_0176_),
    .X(_0191_));
 sky130_fd_sc_hd__or4_1 _0643_ (.A(_0174_),
    .B(_0175_),
    .C(_0180_),
    .D(_0191_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _0644_ (.A(net46),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _0645_ (.A(net45),
    .Y(_0194_));
 sky130_fd_sc_hd__o22a_1 _0646_ (.A1(net7),
    .A2(_0193_),
    .B1(_0194_),
    .B2(net6),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_1 _0647_ (.A1(net7),
    .A2(_0193_),
    .B1(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__o211a_1 _0648_ (.A1(_0182_),
    .A2(_0189_),
    .B1(_0192_),
    .C1(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or2b_1 _0649_ (.A(net54),
    .B_N(net15),
    .X(_0198_));
 sky130_fd_sc_hd__or2b_1 _0650_ (.A(net15),
    .B_N(net54),
    .X(_0199_));
 sky130_fd_sc_hd__nand2_1 _0651_ (.A(_0198_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__and2b_1 _0652_ (.A_N(net16),
    .B(net55),
    .X(_0201_));
 sky130_fd_sc_hd__and2b_1 _0653_ (.A_N(net55),
    .B(net16),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _0654_ (.A(_0201_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _0655_ (.A(_0200_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__or2b_1 _0656_ (.A(net13),
    .B_N(net52),
    .X(_0205_));
 sky130_fd_sc_hd__or2b_1 _0657_ (.A(net52),
    .B_N(net13),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(_0205_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(net53),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _0660_ (.A(_0208_),
    .B(net14),
    .Y(_0209_));
 sky130_fd_sc_hd__and2_1 _0661_ (.A(_0208_),
    .B(net14),
    .X(_0210_));
 sky130_fd_sc_hd__or2_1 _0662_ (.A(_0209_),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__or3_1 _0663_ (.A(_0204_),
    .B(_0207_),
    .C(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__or2b_1 _0664_ (.A(net8),
    .B_N(net47),
    .X(_0213_));
 sky130_fd_sc_hd__or2b_1 _0665_ (.A(net47),
    .B_N(net8),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _0666_ (.A(_0213_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__and2b_1 _0667_ (.A_N(net48),
    .B(net9),
    .X(_0216_));
 sky130_fd_sc_hd__or2b_1 _0668_ (.A(net9),
    .B_N(net48),
    .X(_0217_));
 sky130_fd_sc_hd__or2b_1 _0669_ (.A(_0216_),
    .B_N(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__and2b_1 _0670_ (.A_N(net11),
    .B(net50),
    .X(_0219_));
 sky130_fd_sc_hd__and2b_1 _0671_ (.A_N(net50),
    .B(net11),
    .X(_0220_));
 sky130_fd_sc_hd__and2b_1 _0672_ (.A_N(net10),
    .B(net49),
    .X(_0221_));
 sky130_fd_sc_hd__and2b_1 _0673_ (.A_N(net49),
    .B(net10),
    .X(_0222_));
 sky130_fd_sc_hd__or2_1 _0674_ (.A(_0221_),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__or3_1 _0675_ (.A(_0219_),
    .B(_0220_),
    .C(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__or3_1 _0676_ (.A(_0215_),
    .B(_0218_),
    .C(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__a211o_1 _0677_ (.A1(_0184_),
    .A2(_0197_),
    .B1(_0212_),
    .C1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _0678_ (.A1(_0213_),
    .A2(_0217_),
    .B1(_0216_),
    .X(_0227_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0219_),
    .B(_0221_),
    .Y(_0228_));
 sky130_fd_sc_hd__o22a_1 _0680_ (.A1(_0224_),
    .A2(_0227_),
    .B1(_0228_),
    .B2(_0220_),
    .X(_0229_));
 sky130_fd_sc_hd__o21a_1 _0681_ (.A1(_0208_),
    .A2(net14),
    .B1(_0205_),
    .X(_0230_));
 sky130_fd_sc_hd__or3_1 _0682_ (.A(_0204_),
    .B(_0210_),
    .C(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__o221a_1 _0683_ (.A1(_0199_),
    .A2(_0202_),
    .B1(_0212_),
    .B2(_0229_),
    .C1(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__and2b_1 _0684_ (.A_N(_0201_),
    .B(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__xnor2_1 _0685_ (.A(net59),
    .B(net20),
    .Y(_0234_));
 sky130_fd_sc_hd__and2b_1 _0686_ (.A_N(net19),
    .B(net58),
    .X(_0235_));
 sky130_fd_sc_hd__and2b_1 _0687_ (.A_N(net58),
    .B(net19),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _0688_ (.A(_0235_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _0689_ (.A(_0234_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__and2b_1 _0690_ (.A_N(net18),
    .B(net57),
    .X(_0239_));
 sky130_fd_sc_hd__and2b_1 _0691_ (.A_N(net57),
    .B(net18),
    .X(_0240_));
 sky130_fd_sc_hd__or2_1 _0692_ (.A(_0239_),
    .B(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__or2b_1 _0693_ (.A(net17),
    .B_N(net56),
    .X(_0242_));
 sky130_fd_sc_hd__or2b_1 _0694_ (.A(net56),
    .B_N(net17),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _0695_ (.A(_0242_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__a2111o_1 _0696_ (.A1(_0226_),
    .A2(_0233_),
    .B1(_0238_),
    .C1(_0241_),
    .D1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__and2b_1 _0697_ (.A_N(_0239_),
    .B(_0242_),
    .X(_0246_));
 sky130_fd_sc_hd__or3_1 _0698_ (.A(_0238_),
    .B(_0240_),
    .C(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__inv_2 _0699_ (.A(net20),
    .Y(_0248_));
 sky130_fd_sc_hd__a21o_1 _0700_ (.A1(net59),
    .A2(_0248_),
    .B1(_0235_),
    .X(_0249_));
 sky130_fd_sc_hd__o21ai_1 _0701_ (.A1(net59),
    .A2(_0248_),
    .B1(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__or2b_1 _0702_ (.A(net60),
    .B_N(net21),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _0703_ (.A(_0138_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__a31o_1 _0704_ (.A1(_0245_),
    .A2(_0247_),
    .A3(_0250_),
    .B1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__and2b_1 _0705_ (.A_N(net22),
    .B(net61),
    .X(_0254_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__and2b_1 _0707_ (.A_N(net61),
    .B(net22),
    .X(_0256_));
 sky130_fd_sc_hd__or2b_1 _0708_ (.A(net63),
    .B_N(net24),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _0709_ (.A(_0137_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__a311o_1 _0710_ (.A1(_0138_),
    .A2(_0253_),
    .A3(_0255_),
    .B1(_0256_),
    .C1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__xor2_1 _0711_ (.A(net64),
    .B(net25),
    .X(_0260_));
 sky130_fd_sc_hd__a21oi_1 _0712_ (.A1(_0137_),
    .A2(_0259_),
    .B1(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__or3b_1 _0713_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .B(_0119_),
    .C_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .X(_0262_));
 sky130_fd_sc_hd__a31o_1 _0714_ (.A1(_0137_),
    .A2(_0259_),
    .A3(_0260_),
    .B1(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o22a_1 _0715_ (.A1(_0120_),
    .A2(_0136_),
    .B1(_0261_),
    .B2(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__buf_4 _0716_ (.A(_0117_),
    .X(_0265_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(net64),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21oi_1 _0718_ (.A1(_0118_),
    .A2(_0264_),
    .B1(_0266_),
    .Y(_0086_));
 sky130_fd_sc_hd__clkbuf_4 _0719_ (.A(_0265_),
    .X(_0267_));
 sky130_fd_sc_hd__clkbuf_4 _0720_ (.A(_0116_),
    .X(_0268_));
 sky130_fd_sc_hd__o31ai_1 _0721_ (.A1(net21),
    .A2(net22),
    .A3(_0134_),
    .B1(net24),
    .Y(_0269_));
 sky130_fd_sc_hd__and3_1 _0722_ (.A(_0268_),
    .B(_0135_),
    .C(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__buf_2 _0723_ (.A(_0115_),
    .X(_0271_));
 sky130_fd_sc_hd__a31o_1 _0724_ (.A1(_0138_),
    .A2(_0253_),
    .A3(_0255_),
    .B1(_0256_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _0725_ (.A(_0258_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__clkbuf_4 _0726_ (.A(_0116_),
    .X(_0274_));
 sky130_fd_sc_hd__o21ai_4 _0727_ (.A1(_0115_),
    .A2(_0274_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .Y(_0275_));
 sky130_fd_sc_hd__clkbuf_4 _0728_ (.A(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__a31o_1 _0729_ (.A1(_0271_),
    .A2(_0259_),
    .A3(_0273_),
    .B1(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__o22a_1 _0730_ (.A1(net104),
    .A2(_0267_),
    .B1(_0270_),
    .B2(_0277_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_4 _0731_ (.A(_0115_),
    .X(_0278_));
 sky130_fd_sc_hd__o211ai_1 _0732_ (.A1(_0256_),
    .A2(_0254_),
    .B1(_0253_),
    .C1(_0138_),
    .Y(_0279_));
 sky130_fd_sc_hd__a211o_1 _0733_ (.A1(_0138_),
    .A2(_0253_),
    .B1(_0254_),
    .C1(_0256_),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _0734_ (.A(net21),
    .B(_0134_),
    .X(_0281_));
 sky130_fd_sc_hd__o31ai_2 _0735_ (.A1(net21),
    .A2(net22),
    .A3(_0134_),
    .B1(_0274_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _0736_ (.A1(net22),
    .A2(_0281_),
    .B1(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__a31o_1 _0737_ (.A1(_0278_),
    .A2(_0279_),
    .A3(_0280_),
    .B1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net61),
    .A1(_0284_),
    .S(_0265_),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0285_),
    .X(_0084_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(_0271_),
    .B(_0253_),
    .Y(_0286_));
 sky130_fd_sc_hd__a41oi_1 _0741_ (.A1(_0252_),
    .A2(_0245_),
    .A3(_0247_),
    .A4(_0250_),
    .B1(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__clkbuf_4 _0742_ (.A(_0268_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _0743_ (.A(net21),
    .B(_0134_),
    .Y(_0289_));
 sky130_fd_sc_hd__a31o_1 _0744_ (.A1(_0288_),
    .A2(_0281_),
    .A3(_0289_),
    .B1(_0276_),
    .X(_0290_));
 sky130_fd_sc_hd__o22a_1 _0745_ (.A1(net94),
    .A2(_0267_),
    .B1(_0287_),
    .B2(_0290_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _0746_ (.A(_0226_),
    .B(_0233_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(_0291_),
    .B(_0244_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _0748_ (.A(_0237_),
    .Y(_0293_));
 sky130_fd_sc_hd__a211oi_1 _0749_ (.A1(_0246_),
    .A2(_0292_),
    .B1(_0293_),
    .C1(_0240_),
    .Y(_0294_));
 sky130_fd_sc_hd__o21ai_1 _0750_ (.A1(_0235_),
    .A2(_0294_),
    .B1(_0234_),
    .Y(_0295_));
 sky130_fd_sc_hd__or3_1 _0751_ (.A(_0234_),
    .B(_0235_),
    .C(_0294_),
    .X(_0296_));
 sky130_fd_sc_hd__and3_1 _0752_ (.A(_0271_),
    .B(_0295_),
    .C(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__or2_1 _0753_ (.A(net19),
    .B(_0133_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(net20),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__a31o_1 _0755_ (.A1(_0288_),
    .A2(_0134_),
    .A3(_0299_),
    .B1(_0276_),
    .X(_0300_));
 sky130_fd_sc_hd__o22a_1 _0756_ (.A1(net102),
    .A2(_0267_),
    .B1(_0297_),
    .B2(_0300_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_1 _0757_ (.A(net19),
    .B(_0133_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21oi_1 _0758_ (.A1(_0246_),
    .A2(_0292_),
    .B1(_0240_),
    .Y(_0302_));
 sky130_fd_sc_hd__xnor2_1 _0759_ (.A(_0293_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__a32o_1 _0760_ (.A1(_0268_),
    .A2(_0298_),
    .A3(_0301_),
    .B1(_0303_),
    .B2(_0278_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _0761_ (.A0(net58),
    .A1(_0304_),
    .S(_0265_),
    .X(_0305_));
 sky130_fd_sc_hd__clkbuf_1 _0762_ (.A(_0305_),
    .X(_0081_));
 sky130_fd_sc_hd__a21oi_1 _0763_ (.A1(_0242_),
    .A2(_0292_),
    .B1(_0241_),
    .Y(_0306_));
 sky130_fd_sc_hd__clkbuf_4 _0764_ (.A(_0262_),
    .X(_0307_));
 sky130_fd_sc_hd__a31o_1 _0765_ (.A1(_0241_),
    .A2(_0242_),
    .A3(_0292_),
    .B1(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__nor2_1 _0766_ (.A(_0306_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__or2_1 _0767_ (.A(net17),
    .B(_0132_),
    .X(_0310_));
 sky130_fd_sc_hd__nand2_1 _0768_ (.A(net18),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__a31o_1 _0769_ (.A1(_0288_),
    .A2(_0133_),
    .A3(_0311_),
    .B1(_0276_),
    .X(_0312_));
 sky130_fd_sc_hd__o22a_1 _0770_ (.A1(net87),
    .A2(_0267_),
    .B1(_0309_),
    .B2(_0312_),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _0771_ (.A(_0291_),
    .B(_0244_),
    .Y(_0313_));
 sky130_fd_sc_hd__and3_1 _0772_ (.A(_0271_),
    .B(_0292_),
    .C(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _0773_ (.A(net17),
    .B(_0132_),
    .Y(_0315_));
 sky130_fd_sc_hd__a31o_1 _0774_ (.A1(_0288_),
    .A2(_0310_),
    .A3(_0315_),
    .B1(_0276_),
    .X(_0316_));
 sky130_fd_sc_hd__o22a_1 _0775_ (.A1(net89),
    .A2(_0267_),
    .B1(_0314_),
    .B2(_0316_),
    .X(_0079_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(net15),
    .B(_0131_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _0777_ (.A(net16),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__and3_1 _0778_ (.A(_0268_),
    .B(_0132_),
    .C(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _0779_ (.A1(_0184_),
    .A2(_0197_),
    .B1(_0215_),
    .X(_0320_));
 sky130_fd_sc_hd__a311o_1 _0780_ (.A1(_0213_),
    .A2(_0217_),
    .A3(_0320_),
    .B1(_0223_),
    .C1(_0216_),
    .X(_0321_));
 sky130_fd_sc_hd__a211o_1 _0781_ (.A1(_0228_),
    .A2(_0321_),
    .B1(_0207_),
    .C1(_0220_),
    .X(_0322_));
 sky130_fd_sc_hd__a211o_1 _0782_ (.A1(_0230_),
    .A2(_0322_),
    .B1(_0200_),
    .C1(_0210_),
    .X(_0323_));
 sky130_fd_sc_hd__a21oi_1 _0783_ (.A1(_0199_),
    .A2(_0323_),
    .B1(_0203_),
    .Y(_0324_));
 sky130_fd_sc_hd__a31o_1 _0784_ (.A1(_0199_),
    .A2(_0203_),
    .A3(_0323_),
    .B1(_0307_),
    .X(_0325_));
 sky130_fd_sc_hd__o21ai_1 _0785_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0118_),
    .Y(_0326_));
 sky130_fd_sc_hd__o22a_1 _0786_ (.A1(net91),
    .A2(_0267_),
    .B1(_0319_),
    .B2(_0326_),
    .X(_0078_));
 sky130_fd_sc_hd__a21o_1 _0787_ (.A1(_0230_),
    .A2(_0322_),
    .B1(_0210_),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_1 _0788_ (.A(_0200_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_1 _0789_ (.A(net15),
    .B(_0131_),
    .Y(_0329_));
 sky130_fd_sc_hd__and3_1 _0790_ (.A(_0116_),
    .B(_0317_),
    .C(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__a31o_1 _0791_ (.A1(_0278_),
    .A2(_0323_),
    .A3(_0328_),
    .B1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net54),
    .A1(_0331_),
    .S(_0265_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0793_ (.A(_0332_),
    .X(_0077_));
 sky130_fd_sc_hd__a21oi_1 _0794_ (.A1(_0205_),
    .A2(_0322_),
    .B1(_0211_),
    .Y(_0333_));
 sky130_fd_sc_hd__a31o_1 _0795_ (.A1(_0205_),
    .A2(_0211_),
    .A3(_0322_),
    .B1(_0307_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_1 _0796_ (.A(_0333_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__or3_1 _0797_ (.A(net10),
    .B(net11),
    .C(_0129_),
    .X(_0336_));
 sky130_fd_sc_hd__or2_1 _0798_ (.A(net13),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__nand2_1 _0799_ (.A(net14),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__a31o_1 _0800_ (.A1(_0288_),
    .A2(_0131_),
    .A3(_0338_),
    .B1(_0276_),
    .X(_0339_));
 sky130_fd_sc_hd__o22a_1 _0801_ (.A1(net92),
    .A2(_0267_),
    .B1(_0335_),
    .B2(_0339_),
    .X(_0076_));
 sky130_fd_sc_hd__nand2_1 _0802_ (.A(net13),
    .B(_0336_),
    .Y(_0340_));
 sky130_fd_sc_hd__and3_1 _0803_ (.A(_0268_),
    .B(_0337_),
    .C(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__o311ai_1 _0804_ (.A1(_0218_),
    .A2(_0224_),
    .A3(_0320_),
    .B1(_0229_),
    .C1(_0207_),
    .Y(_0342_));
 sky130_fd_sc_hd__a31o_1 _0805_ (.A1(_0271_),
    .A2(_0322_),
    .A3(_0342_),
    .B1(_0276_),
    .X(_0343_));
 sky130_fd_sc_hd__o22a_1 _0806_ (.A1(net90),
    .A2(_0267_),
    .B1(_0341_),
    .B2(_0343_),
    .X(_0075_));
 sky130_fd_sc_hd__or2_1 _0807_ (.A(net10),
    .B(_0129_),
    .X(_0344_));
 sky130_fd_sc_hd__nand2_1 _0808_ (.A(net11),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _0809_ (.A(_0219_),
    .B(_0220_),
    .Y(_0346_));
 sky130_fd_sc_hd__a311oi_2 _0810_ (.A1(_0213_),
    .A2(_0217_),
    .A3(_0320_),
    .B1(_0223_),
    .C1(_0216_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_1 _0811_ (.A(_0221_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_1 _0812_ (.A(_0346_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a32o_1 _0813_ (.A1(_0268_),
    .A2(_0336_),
    .A3(_0345_),
    .B1(_0349_),
    .B2(_0278_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(net50),
    .A1(_0350_),
    .S(_0265_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0815_ (.A(_0351_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2_1 _0816_ (.A(net10),
    .B(_0129_),
    .Y(_0352_));
 sky130_fd_sc_hd__o211a_1 _0817_ (.A1(_0218_),
    .A2(_0320_),
    .B1(_0227_),
    .C1(_0223_),
    .X(_0353_));
 sky130_fd_sc_hd__nor2_1 _0818_ (.A(_0347_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__a32o_1 _0819_ (.A1(_0274_),
    .A2(_0344_),
    .A3(_0352_),
    .B1(_0354_),
    .B2(_0278_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(net49),
    .A1(_0355_),
    .S(_0265_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0821_ (.A(_0356_),
    .X(_0073_));
 sky130_fd_sc_hd__or3_1 _0822_ (.A(net8),
    .B(_0127_),
    .C(_0128_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(net9),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _0824_ (.A(_0213_),
    .B(_0320_),
    .Y(_0359_));
 sky130_fd_sc_hd__xnor2_1 _0825_ (.A(_0218_),
    .B(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hd__a32o_1 _0826_ (.A1(_0274_),
    .A2(_0129_),
    .A3(_0358_),
    .B1(_0360_),
    .B2(_0278_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _0827_ (.A0(net48),
    .A1(_0361_),
    .S(_0117_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0362_),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _0829_ (.A(_0184_),
    .B(_0197_),
    .C(_0215_),
    .X(_0363_));
 sky130_fd_sc_hd__and3b_1 _0830_ (.A_N(_0363_),
    .B(_0271_),
    .C(_0320_),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_1 _0831_ (.A1(_0127_),
    .A2(_0128_),
    .B1(net8),
    .Y(_0365_));
 sky130_fd_sc_hd__a31o_1 _0832_ (.A1(_0288_),
    .A2(_0357_),
    .A3(_0365_),
    .B1(_0276_),
    .X(_0366_));
 sky130_fd_sc_hd__o22a_1 _0833_ (.A1(net99),
    .A2(_0267_),
    .B1(_0364_),
    .B2(_0366_),
    .X(_0071_));
 sky130_fd_sc_hd__a21o_1 _0834_ (.A1(_0155_),
    .A2(_0161_),
    .B1(_0163_),
    .X(_0367_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(_0367_),
    .B(_0173_),
    .X(_0368_));
 sky130_fd_sc_hd__a21o_1 _0836_ (.A1(_0189_),
    .A2(_0368_),
    .B1(_0178_),
    .X(_0369_));
 sky130_fd_sc_hd__a211o_1 _0837_ (.A1(_0191_),
    .A2(_0369_),
    .B1(_0174_),
    .C1(_0180_),
    .X(_0370_));
 sky130_fd_sc_hd__o21ai_1 _0838_ (.A1(net6),
    .A2(_0194_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__xnor2_1 _0839_ (.A(_0175_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__or2_1 _0840_ (.A(net6),
    .B(_0127_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(net7),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__o21a_1 _0842_ (.A1(_0127_),
    .A2(_0128_),
    .B1(_0274_),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _0843_ (.A1(_0115_),
    .A2(_0372_),
    .B1(_0374_),
    .B2(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(net46),
    .A1(_0376_),
    .S(_0117_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0377_),
    .X(_0070_));
 sky130_fd_sc_hd__a21o_1 _0846_ (.A1(_0191_),
    .A2(_0369_),
    .B1(_0180_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _0847_ (.A(_0174_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _0848_ (.A(net6),
    .B(_0127_),
    .Y(_0380_));
 sky130_fd_sc_hd__and3_1 _0849_ (.A(_0116_),
    .B(_0373_),
    .C(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__a31o_1 _0850_ (.A1(_0278_),
    .A2(_0370_),
    .A3(_0379_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _0851_ (.A0(net45),
    .A1(_0382_),
    .S(_0117_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0852_ (.A(_0383_),
    .X(_0069_));
 sky130_fd_sc_hd__or3_1 _0853_ (.A(net4),
    .B(_0125_),
    .C(_0126_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _0854_ (.A(net5),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__nand2_1 _0855_ (.A(_0176_),
    .B(_0369_),
    .Y(_0386_));
 sky130_fd_sc_hd__xnor2_1 _0856_ (.A(_0181_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__a32o_1 _0857_ (.A1(_0274_),
    .A2(_0127_),
    .A3(_0385_),
    .B1(_0387_),
    .B2(_0278_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(net44),
    .A1(_0388_),
    .S(_0117_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0859_ (.A(_0389_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _0860_ (.A(_0178_),
    .B(_0189_),
    .C(_0368_),
    .X(_0390_));
 sky130_fd_sc_hd__and3b_1 _0861_ (.A_N(_0390_),
    .B(_0271_),
    .C(_0369_),
    .X(_0391_));
 sky130_fd_sc_hd__o21ai_1 _0862_ (.A1(_0125_),
    .A2(_0126_),
    .B1(net4),
    .Y(_0392_));
 sky130_fd_sc_hd__a31o_1 _0863_ (.A1(_0288_),
    .A2(_0384_),
    .A3(_0392_),
    .B1(_0275_),
    .X(_0393_));
 sky130_fd_sc_hd__o22a_1 _0864_ (.A1(net97),
    .A2(_0118_),
    .B1(_0391_),
    .B2(_0393_),
    .X(_0067_));
 sky130_fd_sc_hd__or3_1 _0865_ (.A(_0367_),
    .B(_0169_),
    .C(_0172_),
    .X(_0394_));
 sky130_fd_sc_hd__a21oi_1 _0866_ (.A1(_0186_),
    .A2(_0394_),
    .B1(_0165_),
    .Y(_0395_));
 sky130_fd_sc_hd__o21ba_1 _0867_ (.A1(_0187_),
    .A2(net2),
    .B1_N(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__xnor2_1 _0868_ (.A(_0164_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(net2),
    .B(_0125_),
    .X(_0398_));
 sky130_fd_sc_hd__o21ai_1 _0870_ (.A1(net3),
    .A2(_0398_),
    .B1(_0274_),
    .Y(_0399_));
 sky130_fd_sc_hd__a21o_1 _0871_ (.A1(net3),
    .A2(_0398_),
    .B1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__o211a_1 _0872_ (.A1(_0307_),
    .A2(_0397_),
    .B1(_0400_),
    .C1(_0265_),
    .X(_0401_));
 sky130_fd_sc_hd__a21oi_1 _0873_ (.A1(_0185_),
    .A2(_0276_),
    .B1(_0401_),
    .Y(_0066_));
 sky130_fd_sc_hd__and3_1 _0874_ (.A(_0165_),
    .B(_0186_),
    .C(_0394_),
    .X(_0402_));
 sky130_fd_sc_hd__nor3_1 _0875_ (.A(_0307_),
    .B(_0395_),
    .C(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _0876_ (.A(net2),
    .B(_0125_),
    .Y(_0404_));
 sky130_fd_sc_hd__a31o_1 _0877_ (.A1(_0288_),
    .A2(_0398_),
    .A3(_0404_),
    .B1(_0275_),
    .X(_0405_));
 sky130_fd_sc_hd__o22a_1 _0878_ (.A1(net41),
    .A2(_0118_),
    .B1(_0403_),
    .B2(_0405_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_2 _0879_ (.A(_0121_),
    .B(_0122_),
    .X(_0406_));
 sky130_fd_sc_hd__or3_1 _0880_ (.A(net31),
    .B(_0406_),
    .C(_0123_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(net32),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__and3_1 _0882_ (.A(_0268_),
    .B(_0125_),
    .C(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_1 _0883_ (.A(_0367_),
    .B(_0172_),
    .X(_0410_));
 sky130_fd_sc_hd__a21oi_1 _0884_ (.A1(_0170_),
    .A2(_0410_),
    .B1(_0169_),
    .Y(_0411_));
 sky130_fd_sc_hd__a31o_1 _0885_ (.A1(_0169_),
    .A2(_0170_),
    .A3(_0410_),
    .B1(_0307_),
    .X(_0412_));
 sky130_fd_sc_hd__o21ai_1 _0886_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0265_),
    .Y(_0413_));
 sky130_fd_sc_hd__o22a_1 _0887_ (.A1(net88),
    .A2(_0118_),
    .B1(_0409_),
    .B2(_0413_),
    .X(_0064_));
 sky130_fd_sc_hd__o21ai_1 _0888_ (.A1(_0406_),
    .A2(_0123_),
    .B1(net31),
    .Y(_0414_));
 sky130_fd_sc_hd__and3_1 _0889_ (.A(_0268_),
    .B(_0407_),
    .C(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(_0367_),
    .B(_0172_),
    .Y(_0416_));
 sky130_fd_sc_hd__a31o_1 _0891_ (.A1(_0271_),
    .A2(_0410_),
    .A3(_0416_),
    .B1(_0275_),
    .X(_0417_));
 sky130_fd_sc_hd__o22a_1 _0892_ (.A1(net95),
    .A2(_0118_),
    .B1(_0415_),
    .B2(_0417_),
    .X(_0063_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(net29),
    .B(_0406_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _0894_ (.A(net30),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__o211a_1 _0895_ (.A1(_0406_),
    .A2(_0123_),
    .B1(_0419_),
    .C1(_0288_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _0896_ (.A(net68),
    .B(_0156_),
    .Y(_0421_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(_0421_),
    .B(_0162_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21o_1 _0898_ (.A1(_0155_),
    .A2(_0160_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__or2b_1 _0899_ (.A(_0158_),
    .B_N(_0157_),
    .X(_0424_));
 sky130_fd_sc_hd__a21oi_1 _0900_ (.A1(_0421_),
    .A2(_0423_),
    .B1(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a31o_1 _0901_ (.A1(_0421_),
    .A2(_0424_),
    .A3(_0423_),
    .B1(_0307_),
    .X(_0426_));
 sky130_fd_sc_hd__o21ai_1 _0902_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0265_),
    .Y(_0427_));
 sky130_fd_sc_hd__o22a_1 _0903_ (.A1(net93),
    .A2(_0118_),
    .B1(_0420_),
    .B2(_0427_),
    .X(_0062_));
 sky130_fd_sc_hd__nand3_1 _0904_ (.A(_0155_),
    .B(_0160_),
    .C(_0422_),
    .Y(_0428_));
 sky130_fd_sc_hd__and3_1 _0905_ (.A(_0271_),
    .B(_0423_),
    .C(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(net29),
    .B(_0406_),
    .Y(_0430_));
 sky130_fd_sc_hd__a31o_1 _0907_ (.A1(_0288_),
    .A2(_0418_),
    .A3(_0430_),
    .B1(_0275_),
    .X(_0431_));
 sky130_fd_sc_hd__o22a_1 _0908_ (.A1(net101),
    .A2(_0118_),
    .B1(_0429_),
    .B2(_0431_),
    .X(_0061_));
 sky130_fd_sc_hd__or2_1 _0909_ (.A(net27),
    .B(_0121_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _0910_ (.A(net28),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a31o_1 _0911_ (.A1(_0139_),
    .A2(_0140_),
    .A3(_0146_),
    .B1(_0154_),
    .X(_0434_));
 sky130_fd_sc_hd__o21ai_1 _0912_ (.A1(_0434_),
    .A2(_0152_),
    .B1(_0150_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_1 _0913_ (.A(_0149_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__a32o_1 _0914_ (.A1(_0274_),
    .A2(_0406_),
    .A3(_0433_),
    .B1(_0436_),
    .B2(_0278_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _0915_ (.A0(net67),
    .A1(_0437_),
    .S(_0117_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _0916_ (.A(_0438_),
    .X(_0060_));
 sky130_fd_sc_hd__nand2_1 _0917_ (.A(net27),
    .B(_0121_),
    .Y(_0439_));
 sky130_fd_sc_hd__xor2_1 _0918_ (.A(_0434_),
    .B(_0152_),
    .X(_0440_));
 sky130_fd_sc_hd__a32o_1 _0919_ (.A1(_0274_),
    .A2(_0432_),
    .A3(_0439_),
    .B1(_0440_),
    .B2(_0278_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(net66),
    .A1(_0441_),
    .S(_0117_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0442_),
    .X(_0059_));
 sky130_fd_sc_hd__and2b_1 _0922_ (.A_N(net75),
    .B(net65),
    .X(_0443_));
 sky130_fd_sc_hd__a211o_1 _0923_ (.A1(_0140_),
    .A2(_0146_),
    .B1(_0443_),
    .C1(_0154_),
    .X(_0444_));
 sky130_fd_sc_hd__o211ai_1 _0924_ (.A1(_0443_),
    .A2(_0154_),
    .B1(_0140_),
    .C1(_0146_),
    .Y(_0445_));
 sky130_fd_sc_hd__and3_1 _0925_ (.A(_0271_),
    .B(_0444_),
    .C(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__or2_1 _0926_ (.A(net12),
    .B(_0112_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _0927_ (.A(net23),
    .B(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_1 _0928_ (.A(net26),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a31o_1 _0929_ (.A1(_0268_),
    .A2(net74),
    .A3(_0449_),
    .B1(_0275_),
    .X(_0450_));
 sky130_fd_sc_hd__o22a_1 _0930_ (.A1(net96),
    .A2(_0118_),
    .B1(_0446_),
    .B2(_0450_),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_1 _0931_ (.A(net23),
    .B(_0447_),
    .Y(_0451_));
 sky130_fd_sc_hd__o21a_1 _0932_ (.A1(_0141_),
    .A2(_0145_),
    .B1(_0115_),
    .X(_0452_));
 sky130_fd_sc_hd__a32o_1 _0933_ (.A1(_0274_),
    .A2(_0448_),
    .A3(_0451_),
    .B1(_0452_),
    .B2(_0146_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net62),
    .A1(_0453_),
    .S(_0117_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0454_),
    .X(_0057_));
 sky130_fd_sc_hd__a21oi_1 _0936_ (.A1(_0142_),
    .A2(_0143_),
    .B1(_0307_),
    .Y(_0455_));
 sky130_fd_sc_hd__o21a_1 _0937_ (.A1(_0142_),
    .A2(_0143_),
    .B1(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(net12),
    .B(_0112_),
    .Y(_0457_));
 sky130_fd_sc_hd__a31o_1 _0939_ (.A1(_0268_),
    .A2(_0447_),
    .A3(_0457_),
    .B1(_0275_),
    .X(_0458_));
 sky130_fd_sc_hd__o22a_1 _0940_ (.A1(net108),
    .A2(_0118_),
    .B1(_0456_),
    .B2(_0458_),
    .X(_0056_));
 sky130_fd_sc_hd__o21ai_1 _0941_ (.A1(net40),
    .A2(_0307_),
    .B1(_0120_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(_0112_),
    .B(_0307_),
    .Y(_0460_));
 sky130_fd_sc_hd__o21a_1 _0943_ (.A1(_0276_),
    .A2(_0460_),
    .B1(net40),
    .X(_0461_));
 sky130_fd_sc_hd__a31o_1 _0944_ (.A1(_0112_),
    .A2(_0267_),
    .A3(_0459_),
    .B1(_0461_),
    .X(_0055_));
 sky130_fd_sc_hd__and3b_1 _0945_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .X(_0462_));
 sky130_fd_sc_hd__nor2_1 _0946_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .Y(_0463_));
 sky130_fd_sc_hd__and3_1 _0947_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0462_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__or2_1 _0948_ (.A(net26),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .X(_0465_));
 sky130_fd_sc_hd__or2_1 _0949_ (.A(net23),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .X(_0466_));
 sky130_fd_sc_hd__nand2_1 _0950_ (.A(net12),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .Y(_0467_));
 sky130_fd_sc_hd__or2_1 _0951_ (.A(net12),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .X(_0468_));
 sky130_fd_sc_hd__and4_1 _0952_ (.A(_0112_),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .C(_0467_),
    .D(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__a21o_1 _0953_ (.A1(net12),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _0954_ (.A(net23),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .Y(_0471_));
 sky130_fd_sc_hd__a21bo_1 _0955_ (.A1(_0466_),
    .A2(_0470_),
    .B1_N(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_1 _0956_ (.A(net26),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .Y(_0473_));
 sky130_fd_sc_hd__a21bo_1 _0957_ (.A1(_0465_),
    .A2(_0472_),
    .B1_N(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__xnor2_1 _0958_ (.A(net27),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .Y(_0475_));
 sky130_fd_sc_hd__xnor2_1 _0959_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__and3b_1 _0960_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0462_),
    .C(_0463_),
    .X(_0477_));
 sky130_fd_sc_hd__inv_2 _0961_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .Y(_0478_));
 sky130_fd_sc_hd__and3_1 _0962_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .X(_0479_));
 sky130_fd_sc_hd__and2_1 _0963_ (.A(net64),
    .B(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__and4b_1 _0964_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0462_),
    .C(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .D(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0481_));
 sky130_fd_sc_hd__a21boi_1 _0965_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0480_),
    .B1_N(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__or3_1 _0966_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .X(_0483_));
 sky130_fd_sc_hd__a21oi_1 _0967_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0479_),
    .B1(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__xor2_1 _0968_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(_0462_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nor3_2 _0970_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(_0487_));
 sky130_fd_sc_hd__a31o_1 _0971_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0481_),
    .A3(_0480_),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .X(_0488_));
 sky130_fd_sc_hd__a31o_1 _0972_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0487_),
    .A3(_0479_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__o41a_1 _0973_ (.A1(_0478_),
    .A2(_0482_),
    .A3(_0484_),
    .A4(_0486_),
    .B1(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__a221o_1 _0974_ (.A1(_0464_),
    .A2(_0476_),
    .B1(_0477_),
    .B2(net27),
    .C1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o21a_1 _0975_ (.A1(_0462_),
    .A2(_0487_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _0976_ (.A0(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A1(_0491_),
    .S(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_1 _0977_ (.A(_0493_),
    .X(_0054_));
 sky130_fd_sc_hd__or2b_1 _0978_ (.A(_0486_),
    .B_N(_0492_),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0473_),
    .B(_0465_),
    .Y(_0495_));
 sky130_fd_sc_hd__xnor2_1 _0980_ (.A(_0495_),
    .B(_0472_),
    .Y(_0496_));
 sky130_fd_sc_hd__o21a_1 _0981_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0479_),
    .B1(_0484_),
    .X(_0497_));
 sky130_fd_sc_hd__or2_1 _0982_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .B(_0480_),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _0983_ (.A1(net26),
    .A2(_0477_),
    .B1(_0498_),
    .B2(_0482_),
    .X(_0499_));
 sky130_fd_sc_hd__a211o_1 _0984_ (.A1(_0464_),
    .A2(_0496_),
    .B1(_0497_),
    .C1(_0499_),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _0985_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0494_),
    .B1(_0500_),
    .B2(_0492_),
    .X(_0053_));
 sky130_fd_sc_hd__buf_2 _0986_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand3_1 _0988_ (.A(_0466_),
    .B(_0471_),
    .C(_0470_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21o_1 _0989_ (.A1(_0466_),
    .A2(_0471_),
    .B1(_0470_),
    .X(_0504_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0480_),
    .Y(_0505_));
 sky130_fd_sc_hd__a31o_1 _0991_ (.A1(net64),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A3(_0501_),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .X(_0506_));
 sky130_fd_sc_hd__a32o_1 _0992_ (.A1(_0481_),
    .A2(_0505_),
    .A3(_0506_),
    .B1(_0477_),
    .B2(net23),
    .X(_0507_));
 sky130_fd_sc_hd__a31oi_1 _0993_ (.A1(_0464_),
    .A2(_0503_),
    .A3(_0504_),
    .B1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__o31ai_1 _0994_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0483_),
    .A3(_0502_),
    .B1(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__a21o_1 _0995_ (.A1(_0487_),
    .A2(_0502_),
    .B1(_0494_),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _0996_ (.A1(_0492_),
    .A2(_0509_),
    .B1(_0510_),
    .B2(net98),
    .X(_0052_));
 sky130_fd_sc_hd__or2_1 _0997_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(_0501_),
    .X(_0511_));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(net64),
    .B(_0501_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_1 _0999_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__a22o_1 _1000_ (.A1(_0112_),
    .A2(_0501_),
    .B1(_0467_),
    .B2(_0468_),
    .X(_0514_));
 sky130_fd_sc_hd__and3b_1 _1001_ (.A_N(_0469_),
    .B(_0464_),
    .C(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__a221o_1 _1002_ (.A1(net12),
    .A2(_0477_),
    .B1(_0513_),
    .B2(_0481_),
    .C1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a31o_1 _1003_ (.A1(_0487_),
    .A2(_0502_),
    .A3(_0511_),
    .B1(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__a22o_1 _1004_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A2(_0494_),
    .B1(_0517_),
    .B2(_0492_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _1005_ (.A(net64),
    .B(_0501_),
    .X(_0518_));
 sky130_fd_sc_hd__a21boi_1 _1006_ (.A1(_0112_),
    .A2(_0501_),
    .B1_N(_0464_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_1 _1007_ (.A1(_0477_),
    .A2(_0519_),
    .B1(_0112_),
    .Y(_0520_));
 sky130_fd_sc_hd__o21ai_1 _1008_ (.A1(_0501_),
    .A2(_0483_),
    .B1(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__a31o_1 _1009_ (.A1(_0481_),
    .A2(_0512_),
    .A3(_0518_),
    .B1(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(_0494_),
    .B(_0519_),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _1011_ (.A1(_0492_),
    .A2(_0522_),
    .B1(_0523_),
    .B2(_0501_),
    .X(_0050_));
 sky130_fd_sc_hd__or2_1 _1012_ (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .B(net81),
    .X(_0524_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(net79),
    .B(_0524_),
    .Y(\manchester_baby_instance.BASE_0.s_tickNext ));
 sky130_fd_sc_hd__and3b_1 _1014_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .X(_0525_));
 sky130_fd_sc_hd__and4b_1 _1015_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .C(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .D(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1016_ (.A(_0526_),
    .X(net72));
 sky130_fd_sc_hd__xor2_1 _1017_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .X(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ));
 sky130_fd_sc_hd__a21boi_1 _1018_ (.A1(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .B1_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .Y(_0527_));
 sky130_fd_sc_hd__or2_1 _1019_ (.A(_0525_),
    .B(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1020_ (.A(_0528_),
    .X(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ));
 sky130_fd_sc_hd__and2b_1 _1021_ (.A_N(net73),
    .B(net34),
    .X(_0529_));
 sky130_fd_sc_hd__buf_1 _1022_ (.A(_0529_),
    .X(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ));
 sky130_fd_sc_hd__nor3_2 _1023_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .Y(_0530_));
 sky130_fd_sc_hd__a22o_1 _1024_ (.A1(_0101_),
    .A2(_0463_),
    .B1(_0485_),
    .B2(_0525_),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _1025_ (.A1(_0501_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net35));
 sky130_fd_sc_hd__a22o_1 _1026_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net36));
 sky130_fd_sc_hd__a22o_1 _1027_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net37));
 sky130_fd_sc_hd__a22o_1 _1028_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net38));
 sky130_fd_sc_hd__a22o_1 _1029_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net39));
 sky130_fd_sc_hd__and2b_1 _1030_ (.A_N(net76),
    .B(net77),
    .X(_0532_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0532_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _1032_ (.A(net33),
    .X(_0533_));
 sky130_fd_sc_hd__buf_4 _1033_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(_0534_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(_0534_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(_0534_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(_0534_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(_0534_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(_0534_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(_0534_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1041_ (.A(_0534_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(_0534_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(_0534_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_4 _1044_ (.A(net33),
    .X(_0535_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(_0535_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(_0535_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(_0535_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(_0535_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(_0535_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(_0535_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(_0535_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(_0535_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(_0535_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(_0535_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_4 _1055_ (.A(net33),
    .X(_0536_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0536_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0536_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0536_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0536_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0536_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0536_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0536_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0536_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(_0536_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(_0536_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_4 _1066_ (.A(net33),
    .X(_0537_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0537_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0537_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0537_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0537_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0537_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0537_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0537_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0537_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(_0537_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0537_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(_0533_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(_0533_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(_0533_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(_0533_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(_0533_),
    .Y(_0045_));
 sky130_fd_sc_hd__or2b_1 _1082_ (.A(net83),
    .B_N(\manchester_baby_instance.BASE_0.s_tickReg ),
    .X(_0538_));
 sky130_fd_sc_hd__xnor2_1 _1083_ (.A(net77),
    .B(net84),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(_0533_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(_0533_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1086_ (.A(_0533_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(_0533_),
    .Y(_0049_));
 sky130_fd_sc_hd__and2b_1 _1088_ (.A_N(\manchester_baby_instance.BASE_0.s_tickReg ),
    .B(net83),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1089_ (.A(_0539_),
    .X(_0097_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(net78),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _1091_ (.A(net78),
    .B(net81),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1092_ (.A(_0524_),
    .B(_0540_),
    .Y(_0099_));
 sky130_fd_sc_hd__and2_1 _1093_ (.A(net79),
    .B(_0524_),
    .X(_0541_));
 sky130_fd_sc_hd__clkbuf_1 _1094_ (.A(_0541_),
    .X(_0100_));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_2_1__leaf_clock),
    .D(net76),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _1096_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0000_),
    .Q(\manchester_baby_instance.CIRCUIT_0.Acc.tick ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0050_),
    .RESET_B(_0001_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1098_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0051_),
    .RESET_B(_0002_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1099_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0052_),
    .RESET_B(_0003_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1100_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0053_),
    .RESET_B(_0004_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1101_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0054_),
    .RESET_B(_0005_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0055_),
    .RESET_B(_0006_),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0056_),
    .RESET_B(_0007_),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0057_),
    .RESET_B(_0008_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0058_),
    .RESET_B(_0009_),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0059_),
    .RESET_B(_0010_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0060_),
    .RESET_B(_0011_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0061_),
    .RESET_B(_0012_),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0062_),
    .RESET_B(_0013_),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0063_),
    .RESET_B(_0014_),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0064_),
    .RESET_B(_0015_),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0065_),
    .RESET_B(_0016_),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0066_),
    .RESET_B(_0017_),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0067_),
    .RESET_B(_0018_),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_2 _1115_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0068_),
    .RESET_B(_0019_),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_2 _1116_ (.CLK(clknet_2_2__leaf_clock),
    .D(_0069_),
    .RESET_B(_0020_),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_2 _1117_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0070_),
    .RESET_B(_0021_),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0071_),
    .RESET_B(_0022_),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0072_),
    .RESET_B(_0023_),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0073_),
    .RESET_B(_0024_),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0074_),
    .RESET_B(_0025_),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0075_),
    .RESET_B(_0026_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0076_),
    .RESET_B(_0027_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0077_),
    .RESET_B(_0028_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0078_),
    .RESET_B(_0029_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0079_),
    .RESET_B(_0030_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0080_),
    .RESET_B(_0031_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0081_),
    .RESET_B(_0032_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_2 _1129_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0082_),
    .RESET_B(_0033_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_2_0__leaf_clock),
    .D(_0083_),
    .RESET_B(_0034_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0084_),
    .RESET_B(_0035_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0085_),
    .RESET_B(_0036_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_4 _1133_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0086_),
    .RESET_B(_0037_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0087_),
    .RESET_B(_0038_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0088_),
    .RESET_B(_0039_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0089_),
    .RESET_B(_0040_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0090_),
    .RESET_B(_0041_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0091_),
    .RESET_B(_0042_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _1139_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0092_),
    .RESET_B(_0043_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ));
 sky130_fd_sc_hd__dfrtp_4 _1140_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0093_),
    .RESET_B(_0044_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ));
 sky130_fd_sc_hd__dfrtp_4 _1141_ (.CLK(clknet_2_3__leaf_clock),
    .D(_0094_),
    .RESET_B(_0045_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0095_),
    .Q(\manchester_baby_instance.BASE_1.s_derivedClock ));
 sky130_fd_sc_hd__dfrtp_4 _1143_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[0] ),
    .RESET_B(_0046_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1144_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[1] ),
    .RESET_B(_0047_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1145_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue[2] ),
    .RESET_B(_0048_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(clknet_2_1__leaf_clock),
    .D(net86),
    .RESET_B(_0049_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _1147_ (.CLK(clknet_2_1__leaf_clock),
    .D(net77),
    .Q(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1148_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0097_),
    .Q(\manchester_baby_instance.BASE_1.s_counterValue ));
 sky130_fd_sc_hd__dfxtp_1 _1149_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0098_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1150_ (.CLK(clknet_2_1__leaf_clock),
    .D(net82),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1151_ (.CLK(clknet_2_1__leaf_clock),
    .D(_0100_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1152_ (.CLK(clknet_2_1__leaf_clock),
    .D(net80),
    .Q(\manchester_baby_instance.BASE_0.s_tickReg ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clock (.A(clock),
    .X(clknet_0_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clock (.A(clknet_0_clock),
    .X(clknet_2_0__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clock (.A(clknet_0_clock),
    .X(clknet_2_1__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clock (.A(clknet_0_clock),
    .X(clknet_2_2__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clock (.A(clknet_0_clock),
    .X(clknet_2_3__leaf_clock));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\manchester_baby_instance.BASE_1.s_counterValue ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0538_),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net73),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0096_),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net57),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net71),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net56),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net52),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(net55),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net53),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net69),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net60),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net70),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net65),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net43),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net47),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net68),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net59),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net63),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net51),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\manchester_baby_instance.BASE_0.s_tickNext ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0099_),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input1 (.A(ram_data_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(ram_data_i[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(ram_data_i[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(ram_data_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(ram_data_i[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(ram_data_i[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(ram_data_i[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(ram_data_i[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(ram_data_i[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(ram_data_i[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(ram_data_i[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ram_data_i[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(ram_data_i[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(ram_data_i[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(ram_data_i[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(ram_data_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(ram_data_i[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(ram_data_i[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_8 input26 (.A(ram_data_i[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(ram_data_i[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(ram_data_i[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(ram_data_i[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(ram_data_i[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(ram_data_i[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(ram_data_i[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(ram_data_i[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(reset_i),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input4 (.A(ram_data_i[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(ram_data_i[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(ram_data_i[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ram_data_i[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(ram_data_i[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(ram_data_i[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output34 (.A(net34),
    .X(clock_o));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net35),
    .X(ram_addr_o[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(ram_addr_o[1]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(ram_addr_o[2]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(ram_addr_o[3]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(ram_addr_o[4]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(ram_data_o[0]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(ram_data_o[10]));
 sky130_fd_sc_hd__buf_2 output42 (.A(net42),
    .X(ram_data_o[11]));
 sky130_fd_sc_hd__buf_2 output43 (.A(net43),
    .X(ram_data_o[12]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(ram_data_o[13]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(ram_data_o[14]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(ram_data_o[15]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(ram_data_o[16]));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(ram_data_o[17]));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(ram_data_o[18]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(ram_data_o[19]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(ram_data_o[1]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(ram_data_o[20]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(ram_data_o[21]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(ram_data_o[22]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(ram_data_o[23]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(ram_data_o[24]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(ram_data_o[25]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(ram_data_o[26]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(ram_data_o[27]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(ram_data_o[28]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(ram_data_o[29]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(ram_data_o[2]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(ram_data_o[30]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(ram_data_o[31]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(ram_data_o[3]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(ram_data_o[4]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(ram_data_o[5]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(ram_data_o[6]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(ram_data_o[7]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(ram_data_o[8]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ram_data_o[9]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(ram_rw_en_o));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(stop_lamp_o));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(_0121_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net26),
    .X(net75));
endmodule

