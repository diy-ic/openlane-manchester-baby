magic
tech sky130A
magscale 1 2
timestamp 1700142112
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 934 2128 38902 37584
<< metal2 >>
rect 15474 39200 15530 40000
rect 17406 39200 17462 40000
rect 19338 39200 19394 40000
rect 21914 39200 21970 40000
rect 23202 39200 23258 40000
rect 10966 0 11022 800
rect 14186 0 14242 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 23202 0 23258 800
rect 25134 0 25190 800
rect 28998 0 29054 800
<< obsm2 >>
rect 938 39144 15418 39200
rect 15586 39144 17350 39200
rect 17518 39144 19282 39200
rect 19450 39144 21858 39200
rect 22026 39144 23146 39200
rect 23314 39144 38898 39200
rect 938 856 38898 39144
rect 938 800 10910 856
rect 11078 800 14130 856
rect 14298 800 17994 856
rect 18162 800 18638 856
rect 18806 800 19282 856
rect 19450 800 21214 856
rect 21382 800 23146 856
rect 23314 800 25078 856
rect 25246 800 28942 856
rect 29110 800 38898 856
<< metal3 >>
rect 0 29928 800 30048
rect 39200 25848 40000 25968
rect 0 25168 800 25288
rect 39200 25168 40000 25288
rect 0 24488 800 24608
rect 39200 24488 40000 24608
rect 39200 23128 40000 23248
rect 0 22448 800 22568
rect 0 21768 800 21888
rect 0 20408 800 20528
rect 0 19728 800 19848
rect 39200 19728 40000 19848
rect 39200 19048 40000 19168
rect 0 18368 800 18488
rect 39200 18368 40000 18488
rect 39200 17688 40000 17808
rect 39200 17008 40000 17128
rect 39200 16328 40000 16448
rect 0 15648 800 15768
rect 39200 15648 40000 15768
rect 39200 14968 40000 15088
rect 39200 14288 40000 14408
rect 0 13608 800 13728
rect 39200 12248 40000 12368
rect 0 11568 800 11688
rect 39200 10208 40000 10328
rect 39200 8168 40000 8288
<< obsm3 >>
rect 800 30128 39200 37569
rect 880 29848 39200 30128
rect 800 26048 39200 29848
rect 800 25768 39120 26048
rect 800 25368 39200 25768
rect 880 25088 39120 25368
rect 800 24688 39200 25088
rect 880 24408 39120 24688
rect 800 23328 39200 24408
rect 800 23048 39120 23328
rect 800 22648 39200 23048
rect 880 22368 39200 22648
rect 800 21968 39200 22368
rect 880 21688 39200 21968
rect 800 20608 39200 21688
rect 880 20328 39200 20608
rect 800 19928 39200 20328
rect 880 19648 39120 19928
rect 800 19248 39200 19648
rect 800 18968 39120 19248
rect 800 18568 39200 18968
rect 880 18288 39120 18568
rect 800 17888 39200 18288
rect 800 17608 39120 17888
rect 800 17208 39200 17608
rect 800 16928 39120 17208
rect 800 16528 39200 16928
rect 800 16248 39120 16528
rect 800 15848 39200 16248
rect 880 15568 39120 15848
rect 800 15168 39200 15568
rect 800 14888 39120 15168
rect 800 14488 39200 14888
rect 800 14208 39120 14488
rect 800 13808 39200 14208
rect 880 13528 39200 13808
rect 800 12448 39200 13528
rect 800 12168 39120 12448
rect 800 11768 39200 12168
rect 880 11488 39200 11768
rect 800 10408 39200 11488
rect 800 10128 39120 10408
rect 800 8368 39200 10128
rect 800 8088 39120 8368
rect 800 2143 39200 8088
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2128 5188 37584
rect 34928 2128 35248 37584
rect 35588 2128 35908 37584
<< obsm4 >>
rect 18643 16491 25149 23221
<< metal5 >>
rect 1056 36642 38872 36962
rect 1056 35982 38872 36302
rect 1056 6006 38872 6326
rect 1056 5346 38872 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38872 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38872 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38872 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38872 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 29928 800 30048 6 clock
port 3 nsew signal input
rlabel metal2 s 19338 39200 19394 40000 6 ram_addr_o[0]
port 4 nsew signal output
rlabel metal2 s 17406 39200 17462 40000 6 ram_addr_o[1]
port 5 nsew signal output
rlabel metal2 s 15474 39200 15530 40000 6 ram_addr_o[2]
port 6 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 ram_addr_o[3]
port 7 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 ram_addr_o[4]
port 8 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 ram_data_io[0]
port 9 nsew signal bidirectional
rlabel metal2 s 18050 0 18106 800 6 ram_data_io[10]
port 10 nsew signal bidirectional
rlabel metal2 s 21270 0 21326 800 6 ram_data_io[11]
port 11 nsew signal bidirectional
rlabel metal2 s 18694 0 18750 800 6 ram_data_io[12]
port 12 nsew signal bidirectional
rlabel metal2 s 19338 0 19394 800 6 ram_data_io[13]
port 13 nsew signal bidirectional
rlabel metal3 s 39200 16328 40000 16448 6 ram_data_io[14]
port 14 nsew signal bidirectional
rlabel metal3 s 39200 14288 40000 14408 6 ram_data_io[15]
port 15 nsew signal bidirectional
rlabel metal2 s 23202 0 23258 800 6 ram_data_io[16]
port 16 nsew signal bidirectional
rlabel metal2 s 25134 0 25190 800 6 ram_data_io[17]
port 17 nsew signal bidirectional
rlabel metal2 s 28998 0 29054 800 6 ram_data_io[18]
port 18 nsew signal bidirectional
rlabel metal3 s 39200 10208 40000 10328 6 ram_data_io[19]
port 19 nsew signal bidirectional
rlabel metal3 s 0 21768 800 21888 6 ram_data_io[1]
port 20 nsew signal bidirectional
rlabel metal3 s 39200 12248 40000 12368 6 ram_data_io[20]
port 21 nsew signal bidirectional
rlabel metal3 s 39200 14968 40000 15088 6 ram_data_io[21]
port 22 nsew signal bidirectional
rlabel metal3 s 39200 15648 40000 15768 6 ram_data_io[22]
port 23 nsew signal bidirectional
rlabel metal3 s 39200 18368 40000 18488 6 ram_data_io[23]
port 24 nsew signal bidirectional
rlabel metal3 s 39200 19728 40000 19848 6 ram_data_io[24]
port 25 nsew signal bidirectional
rlabel metal3 s 39200 24488 40000 24608 6 ram_data_io[25]
port 26 nsew signal bidirectional
rlabel metal3 s 39200 25848 40000 25968 6 ram_data_io[26]
port 27 nsew signal bidirectional
rlabel metal3 s 39200 25168 40000 25288 6 ram_data_io[27]
port 28 nsew signal bidirectional
rlabel metal3 s 39200 23128 40000 23248 6 ram_data_io[28]
port 29 nsew signal bidirectional
rlabel metal3 s 39200 17688 40000 17808 6 ram_data_io[29]
port 30 nsew signal bidirectional
rlabel metal3 s 0 22448 800 22568 6 ram_data_io[2]
port 31 nsew signal bidirectional
rlabel metal3 s 39200 19048 40000 19168 6 ram_data_io[30]
port 32 nsew signal bidirectional
rlabel metal2 s 23202 39200 23258 40000 6 ram_data_io[31]
port 33 nsew signal bidirectional
rlabel metal3 s 0 19728 800 19848 6 ram_data_io[3]
port 34 nsew signal bidirectional
rlabel metal3 s 0 18368 800 18488 6 ram_data_io[4]
port 35 nsew signal bidirectional
rlabel metal3 s 0 15648 800 15768 6 ram_data_io[5]
port 36 nsew signal bidirectional
rlabel metal3 s 0 13608 800 13728 6 ram_data_io[6]
port 37 nsew signal bidirectional
rlabel metal3 s 0 11568 800 11688 6 ram_data_io[7]
port 38 nsew signal bidirectional
rlabel metal2 s 10966 0 11022 800 6 ram_data_io[8]
port 39 nsew signal bidirectional
rlabel metal2 s 14186 0 14242 800 6 ram_data_io[9]
port 40 nsew signal bidirectional
rlabel metal3 s 39200 8168 40000 8288 6 ram_rw_en_o
port 41 nsew signal output
rlabel metal3 s 39200 17008 40000 17128 6 reset_i
port 42 nsew signal input
rlabel metal2 s 21914 39200 21970 40000 6 stop_lamp_o
port 43 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2673270
string GDS_FILE /openlane/designs/openlane-manchester-baby/runs/RUN_2023.11.16_13.39.35/results/signoff/openlane_manchester_baby.magic.gds
string GDS_START 584702
<< end >>

