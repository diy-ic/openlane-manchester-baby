// This is the unpowered netlist.
module openlane_manchester_baby (clock,
    ram_rw_en_o,
    reset_i,
    stop_lamp_o,
    ram_addr_o,
    ram_data_io);
 input clock;
 output ram_rw_en_o;
 input reset_i;
 output stop_lamp_o;
 output [4:0] ram_addr_o;
 inout [31:0] ram_data_io;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire clknet_0_clock;
 wire clknet_3_0__leaf_clock;
 wire clknet_3_1__leaf_clock;
 wire clknet_3_2__leaf_clock;
 wire clknet_3_3__leaf_clock;
 wire clknet_3_4__leaf_clock;
 wire clknet_3_5__leaf_clock;
 wire clknet_3_6__leaf_clock;
 wire clknet_3_7__leaf_clock;
 wire \manchester_baby_instance.BASE_0.s_countReg[0] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[10] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[11] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[12] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[13] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[14] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[15] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[16] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[17] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[18] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[19] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[1] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[20] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[21] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[22] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[23] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[24] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[25] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[2] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[3] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[4] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[5] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[6] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[7] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[8] ;
 wire \manchester_baby_instance.BASE_0.s_countReg[9] ;
 wire \manchester_baby_instance.BASE_0.s_tickNext ;
 wire \manchester_baby_instance.BASE_0.s_tickReg ;
 wire \manchester_baby_instance.BASE_1.s_bufferRegs[0] ;
 wire \manchester_baby_instance.BASE_1.s_counterValue ;
 wire \manchester_baby_instance.BASE_1.s_derivedClock ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.Acc.tick ;
 wire \manchester_baby_instance.CIRCUIT_0.GATES_13.input1 ;
 wire \manchester_baby_instance.CIRCUIT_0.GATES_13.result ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[13] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[14] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[15] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[2] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[3] ;
 wire \manchester_baby_instance.CIRCUIT_0.IR.q[4] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ;
 wire \manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ;
 wire \manchester_baby_instance.ram_data_i_0 ;
 wire \manchester_baby_instance.ram_data_i_1 ;
 wire \manchester_baby_instance.ram_data_i_10 ;
 wire \manchester_baby_instance.ram_data_i_11 ;
 wire \manchester_baby_instance.ram_data_i_12 ;
 wire \manchester_baby_instance.ram_data_i_13 ;
 wire \manchester_baby_instance.ram_data_i_14 ;
 wire \manchester_baby_instance.ram_data_i_15 ;
 wire \manchester_baby_instance.ram_data_i_16 ;
 wire \manchester_baby_instance.ram_data_i_17 ;
 wire \manchester_baby_instance.ram_data_i_18 ;
 wire \manchester_baby_instance.ram_data_i_19 ;
 wire \manchester_baby_instance.ram_data_i_2 ;
 wire \manchester_baby_instance.ram_data_i_20 ;
 wire \manchester_baby_instance.ram_data_i_21 ;
 wire \manchester_baby_instance.ram_data_i_22 ;
 wire \manchester_baby_instance.ram_data_i_23 ;
 wire \manchester_baby_instance.ram_data_i_24 ;
 wire \manchester_baby_instance.ram_data_i_25 ;
 wire \manchester_baby_instance.ram_data_i_26 ;
 wire \manchester_baby_instance.ram_data_i_27 ;
 wire \manchester_baby_instance.ram_data_i_28 ;
 wire \manchester_baby_instance.ram_data_i_29 ;
 wire \manchester_baby_instance.ram_data_i_3 ;
 wire \manchester_baby_instance.ram_data_i_30 ;
 wire \manchester_baby_instance.ram_data_i_31 ;
 wire \manchester_baby_instance.ram_data_i_4 ;
 wire \manchester_baby_instance.ram_data_i_5 ;
 wire \manchester_baby_instance.ram_data_i_6 ;
 wire \manchester_baby_instance.ram_data_i_7 ;
 wire \manchester_baby_instance.ram_data_i_8 ;
 wire \manchester_baby_instance.ram_data_i_9 ;
 wire \manchester_baby_instance.ram_data_o_0 ;
 wire \manchester_baby_instance.ram_data_o_1 ;
 wire \manchester_baby_instance.ram_data_o_10 ;
 wire \manchester_baby_instance.ram_data_o_11 ;
 wire \manchester_baby_instance.ram_data_o_12 ;
 wire \manchester_baby_instance.ram_data_o_13 ;
 wire \manchester_baby_instance.ram_data_o_14 ;
 wire \manchester_baby_instance.ram_data_o_15 ;
 wire \manchester_baby_instance.ram_data_o_16 ;
 wire \manchester_baby_instance.ram_data_o_17 ;
 wire \manchester_baby_instance.ram_data_o_18 ;
 wire \manchester_baby_instance.ram_data_o_19 ;
 wire \manchester_baby_instance.ram_data_o_2 ;
 wire \manchester_baby_instance.ram_data_o_20 ;
 wire \manchester_baby_instance.ram_data_o_21 ;
 wire \manchester_baby_instance.ram_data_o_22 ;
 wire \manchester_baby_instance.ram_data_o_23 ;
 wire \manchester_baby_instance.ram_data_o_24 ;
 wire \manchester_baby_instance.ram_data_o_25 ;
 wire \manchester_baby_instance.ram_data_o_26 ;
 wire \manchester_baby_instance.ram_data_o_27 ;
 wire \manchester_baby_instance.ram_data_o_28 ;
 wire \manchester_baby_instance.ram_data_o_29 ;
 wire \manchester_baby_instance.ram_data_o_3 ;
 wire \manchester_baby_instance.ram_data_o_30 ;
 wire \manchester_baby_instance.ram_data_o_31 ;
 wire \manchester_baby_instance.ram_data_o_4 ;
 wire \manchester_baby_instance.ram_data_o_5 ;
 wire \manchester_baby_instance.ram_data_o_6 ;
 wire \manchester_baby_instance.ram_data_o_7 ;
 wire \manchester_baby_instance.ram_data_o_8 ;
 wire \manchester_baby_instance.ram_data_o_9 ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net24;
 wire net25;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net52;
 wire net54;
 wire net55;
 wire net56;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net65;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_206 ();
 sky130_fd_sc_hd__and3b_1 _0676_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .C(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .X(_0124_));
 sky130_fd_sc_hd__nor2_1 _0677_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .Y(_0125_));
 sky130_fd_sc_hd__and2_1 _0678_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0125_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__or2_1 _0680_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .X(_0128_));
 sky130_fd_sc_hd__nor2_2 _0681_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__o21a_1 _0682_ (.A1(_0124_),
    .A2(_0129_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .X(_0130_));
 sky130_fd_sc_hd__a21bo_1 _0683_ (.A1(_0124_),
    .A2(_0127_),
    .B1_N(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_4 _0684_ (.A(\manchester_baby_instance.ram_data_i_2 ),
    .X(_0132_));
 sky130_fd_sc_hd__nor2_1 _0685_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0132_),
    .Y(_0133_));
 sky130_fd_sc_hd__buf_2 _0686_ (.A(\manchester_baby_instance.ram_data_i_1 ),
    .X(_0134_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _0688_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .Y(_0136_));
 sky130_fd_sc_hd__or2_1 _0689_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(_0134_),
    .X(_0137_));
 sky130_fd_sc_hd__and3b_1 _0690_ (.A_N(_0136_),
    .B(_0137_),
    .C(_0135_),
    .X(_0138_));
 sky130_fd_sc_hd__inv_2 _0691_ (.A(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__and2_1 _0692_ (.A(_0135_),
    .B(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0132_),
    .Y(_0141_));
 sky130_fd_sc_hd__o21ai_1 _0694_ (.A1(_0133_),
    .A2(_0140_),
    .B1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__o21a_1 _0695_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(\manchester_baby_instance.ram_data_i_3 ),
    .B1(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _0696_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(\manchester_baby_instance.ram_data_i_3 ),
    .B1(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__xnor2_1 _0697_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__and2_1 _0698_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__nor2_1 _0699_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0145_),
    .Y(_0147_));
 sky130_fd_sc_hd__and3_2 _0700_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0124_),
    .C(_0125_),
    .X(_0148_));
 sky130_fd_sc_hd__o21a_1 _0701_ (.A1(_0146_),
    .A2(_0147_),
    .B1(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__and3b_1 _0702_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0124_),
    .C(_0126_),
    .X(_0150_));
 sky130_fd_sc_hd__inv_2 _0703_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .Y(_0151_));
 sky130_fd_sc_hd__o21a_1 _0704_ (.A1(_0129_),
    .A2(_0150_),
    .B1(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__and3_1 _0705_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .C(\manchester_baby_instance.ram_data_o_31 ),
    .X(_0153_));
 sky130_fd_sc_hd__a21boi_1 _0706_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0153_),
    .B1_N(_0150_),
    .Y(_0154_));
 sky130_fd_sc_hd__and3_1 _0707_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .C(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .X(_0155_));
 sky130_fd_sc_hd__and2b_1 _0708_ (.A_N(_0155_),
    .B(_0129_),
    .X(_0156_));
 sky130_fd_sc_hd__o31a_1 _0709_ (.A1(_0152_),
    .A2(_0154_),
    .A3(_0156_),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .X(_0157_));
 sky130_fd_sc_hd__and3b_1 _0710_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .B(_0124_),
    .C(_0125_),
    .X(_0158_));
 sky130_fd_sc_hd__a21o_1 _0711_ (.A1(\manchester_baby_instance.ram_data_o_31 ),
    .A2(_0150_),
    .B1(_0129_),
    .X(_0159_));
 sky130_fd_sc_hd__and4b_1 _0712_ (.A_N(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .C(_0155_),
    .D(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__a21oi_1 _0713_ (.A1(\manchester_baby_instance.ram_data_i_4 ),
    .A2(_0158_),
    .B1(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__or3b_1 _0714_ (.A(_0149_),
    .B(_0157_),
    .C_N(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _0715_ (.A1(net68),
    .A2(_0131_),
    .B1(_0162_),
    .B2(_0130_),
    .X(_0123_));
 sky130_fd_sc_hd__xnor2_1 _0716_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .B(\manchester_baby_instance.ram_data_i_3 ),
    .Y(_0163_));
 sky130_fd_sc_hd__xnor2_1 _0717_ (.A(_0142_),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__a22o_1 _0718_ (.A1(\manchester_baby_instance.ram_data_i_3 ),
    .A2(_0158_),
    .B1(_0164_),
    .B2(_0148_),
    .X(_0165_));
 sky130_fd_sc_hd__a31o_1 _0719_ (.A1(_0151_),
    .A2(_0155_),
    .A3(_0159_),
    .B1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__or3_1 _0720_ (.A(_0131_),
    .B(_0154_),
    .C(_0156_),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _0721_ (.A1(_0130_),
    .A2(_0166_),
    .B1(_0167_),
    .B2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .X(_0122_));
 sky130_fd_sc_hd__a21o_1 _0722_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A2(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .X(_0168_));
 sky130_fd_sc_hd__or2_1 _0723_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0132_),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_1 _0724_ (.A(_0141_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__xor2_1 _0725_ (.A(_0140_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__or2_1 _0726_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .B(_0153_),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(_0148_),
    .A2(_0171_),
    .B1(_0172_),
    .B2(_0154_),
    .X(_0173_));
 sky130_fd_sc_hd__a221o_1 _0728_ (.A1(_0132_),
    .A2(_0158_),
    .B1(_0168_),
    .B2(_0156_),
    .C1(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _0729_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0131_),
    .B1(_0174_),
    .B2(_0130_),
    .X(_0121_));
 sky130_fd_sc_hd__xor2_1 _0730_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .X(_0175_));
 sky130_fd_sc_hd__a21bo_1 _0731_ (.A1(_0135_),
    .A2(_0137_),
    .B1_N(_0136_),
    .X(_0176_));
 sky130_fd_sc_hd__a21oi_1 _0732_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .A2(\manchester_baby_instance.ram_data_o_31 ),
    .B1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _0733_ (.A(_0153_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__a32o_1 _0734_ (.A1(_0148_),
    .A2(_0139_),
    .A3(_0176_),
    .B1(_0178_),
    .B2(_0150_),
    .X(_0179_));
 sky130_fd_sc_hd__a221o_1 _0735_ (.A1(_0134_),
    .A2(_0158_),
    .B1(_0175_),
    .B2(_0129_),
    .C1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _0736_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A2(_0131_),
    .B1(_0180_),
    .B2(_0130_),
    .X(_0120_));
 sky130_fd_sc_hd__inv_2 _0737_ (.A(\manchester_baby_instance.ram_data_o_31 ),
    .Y(_0181_));
 sky130_fd_sc_hd__a22o_1 _0738_ (.A1(_0148_),
    .A2(_0136_),
    .B1(_0150_),
    .B2(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__inv_2 _0739_ (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .Y(_0183_));
 sky130_fd_sc_hd__a21o_1 _0740_ (.A1(_0148_),
    .A2(_0136_),
    .B1(_0158_),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _0741_ (.A1(_0183_),
    .A2(_0159_),
    .B1(_0184_),
    .B2(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0185_));
 sky130_fd_sc_hd__a21o_1 _0742_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .A2(_0182_),
    .B1(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _0743_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .A2(_0131_),
    .B1(_0186_),
    .B2(_0130_),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0745_ (.A(_0187_),
    .B(_0128_),
    .Y(_0188_));
 sky130_fd_sc_hd__a41o_1 _0746_ (.A1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .A2(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A3(_0126_),
    .A4(_0188_),
    .B1(net60),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _0747_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .Y(_0089_));
 sky130_fd_sc_hd__and4_1 _0748_ (.A(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .B(_0089_),
    .C(_0187_),
    .D(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .X(_0189_));
 sky130_fd_sc_hd__buf_2 _0749_ (.A(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .A1(\manchester_baby_instance.ram_data_i_15 ),
    .S(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0191_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .A1(\manchester_baby_instance.ram_data_i_14 ),
    .S(_0190_),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0192_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .A1(\manchester_baby_instance.ram_data_i_13 ),
    .S(_0190_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_1 _0755_ (.A(_0193_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(net72),
    .A1(\manchester_baby_instance.ram_data_i_4 ),
    .S(_0190_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0194_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(net75),
    .A1(\manchester_baby_instance.ram_data_i_3 ),
    .S(_0190_),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _0759_ (.A(_0195_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(net73),
    .A1(_0132_),
    .S(_0190_),
    .X(_0196_));
 sky130_fd_sc_hd__clkbuf_1 _0761_ (.A(_0196_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0762_ (.A0(net71),
    .A1(_0134_),
    .S(_0190_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_1 _0763_ (.A(_0197_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(net70),
    .A1(\manchester_baby_instance.ram_data_i_0 ),
    .S(_0190_),
    .X(_0198_));
 sky130_fd_sc_hd__clkbuf_1 _0765_ (.A(_0198_),
    .X(_0079_));
 sky130_fd_sc_hd__and2b_1 _0766_ (.A_N(\manchester_baby_instance.ram_data_o_29 ),
    .B(\manchester_baby_instance.ram_data_i_29 ),
    .X(_0199_));
 sky130_fd_sc_hd__and2b_1 _0767_ (.A_N(\manchester_baby_instance.ram_data_o_30 ),
    .B(\manchester_baby_instance.ram_data_i_30 ),
    .X(_0200_));
 sky130_fd_sc_hd__and2b_1 _0768_ (.A_N(\manchester_baby_instance.ram_data_i_30 ),
    .B(\manchester_baby_instance.ram_data_o_30 ),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(_0200_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__or2_1 _0770_ (.A(_0199_),
    .B(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__inv_2 _0771_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .Y(_0204_));
 sky130_fd_sc_hd__and2b_1 _0772_ (.A_N(\manchester_baby_instance.ram_data_i_29 ),
    .B(\manchester_baby_instance.ram_data_o_29 ),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _0773_ (.A(_0199_),
    .B(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__o21a_1 _0774_ (.A1(\manchester_baby_instance.ram_data_o_28 ),
    .A2(_0204_),
    .B1(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__xor2_1 _0775_ (.A(\manchester_baby_instance.ram_data_o_28 ),
    .B(\manchester_baby_instance.ram_data_i_28 ),
    .X(_0208_));
 sky130_fd_sc_hd__or2b_1 _0776_ (.A(\manchester_baby_instance.ram_data_o_27 ),
    .B_N(\manchester_baby_instance.ram_data_i_27 ),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _0777_ (.A(_0208_),
    .B(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__and2b_1 _0778_ (.A_N(\manchester_baby_instance.ram_data_o_6 ),
    .B(\manchester_baby_instance.ram_data_i_6 ),
    .X(_0211_));
 sky130_fd_sc_hd__xnor2_1 _0779_ (.A(\manchester_baby_instance.ram_data_o_7 ),
    .B(\manchester_baby_instance.ram_data_i_7 ),
    .Y(_0212_));
 sky130_fd_sc_hd__xnor2_1 _0780_ (.A(_0211_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__and2b_1 _0781_ (.A_N(\manchester_baby_instance.ram_data_o_5 ),
    .B(\manchester_baby_instance.ram_data_i_5 ),
    .X(_0214_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(\manchester_baby_instance.ram_data_o_6 ),
    .B(\manchester_baby_instance.ram_data_i_6 ),
    .Y(_0215_));
 sky130_fd_sc_hd__xnor2_2 _0783_ (.A(_0214_),
    .B(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _0784_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .Y(_0217_));
 sky130_fd_sc_hd__xor2_1 _0785_ (.A(\manchester_baby_instance.ram_data_o_5 ),
    .B(\manchester_baby_instance.ram_data_i_5 ),
    .X(_0218_));
 sky130_fd_sc_hd__o21ai_1 _0786_ (.A1(_0217_),
    .A2(\manchester_baby_instance.ram_data_o_4 ),
    .B1(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__xor2_2 _0787_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(\manchester_baby_instance.ram_data_o_4 ),
    .X(_0220_));
 sky130_fd_sc_hd__nand2b_2 _0788_ (.A_N(\manchester_baby_instance.ram_data_o_3 ),
    .B(\manchester_baby_instance.ram_data_i_3 ),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _0789_ (.A(_0220_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__or3_1 _0790_ (.A(_0217_),
    .B(\manchester_baby_instance.ram_data_o_4 ),
    .C(_0218_),
    .X(_0223_));
 sky130_fd_sc_hd__a21bo_1 _0791_ (.A1(_0219_),
    .A2(_0222_),
    .B1_N(_0223_),
    .X(_0224_));
 sky130_fd_sc_hd__or2_1 _0792_ (.A(_0214_),
    .B(_0215_),
    .X(_0225_));
 sky130_fd_sc_hd__a21o_1 _0793_ (.A1(_0211_),
    .A2(_0212_),
    .B1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _0794_ (.A(_0211_),
    .B(_0212_),
    .X(_0227_));
 sky130_fd_sc_hd__o311a_1 _0795_ (.A1(_0213_),
    .A2(_0216_),
    .A3(_0224_),
    .B1(_0226_),
    .C1(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__or2_1 _0796_ (.A(_0213_),
    .B(_0216_),
    .X(_0229_));
 sky130_fd_sc_hd__or2b_1 _0797_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B_N(\manchester_baby_instance.ram_data_o_3 ),
    .X(_0230_));
 sky130_fd_sc_hd__and4b_1 _0798_ (.A_N(\manchester_baby_instance.ram_data_o_2 ),
    .B(_0221_),
    .C(_0230_),
    .D(_0132_),
    .X(_0231_));
 sky130_fd_sc_hd__inv_2 _0799_ (.A(\manchester_baby_instance.ram_data_i_0 ),
    .Y(_0232_));
 sky130_fd_sc_hd__and2b_1 _0800_ (.A_N(\manchester_baby_instance.ram_data_o_1 ),
    .B(_0134_),
    .X(_0233_));
 sky130_fd_sc_hd__and2b_1 _0801_ (.A_N(_0134_),
    .B(\manchester_baby_instance.ram_data_o_1 ),
    .X(_0234_));
 sky130_fd_sc_hd__o22a_2 _0802_ (.A1(_0232_),
    .A2(\manchester_baby_instance.ram_data_o_0 ),
    .B1(_0233_),
    .B2(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__xor2_2 _0803_ (.A(_0132_),
    .B(\manchester_baby_instance.ram_data_o_2 ),
    .X(_0236_));
 sky130_fd_sc_hd__xnor2_2 _0804_ (.A(_0236_),
    .B(_0233_),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _0805_ (.A(_0132_),
    .Y(_0238_));
 sky130_fd_sc_hd__o2bb2a_1 _0806_ (.A1_N(_0221_),
    .A2_N(_0230_),
    .B1(_0238_),
    .B2(\manchester_baby_instance.ram_data_o_2 ),
    .X(_0239_));
 sky130_fd_sc_hd__inv_2 _0807_ (.A(_0134_),
    .Y(_0240_));
 sky130_fd_sc_hd__o21a_1 _0808_ (.A1(_0240_),
    .A2(\manchester_baby_instance.ram_data_o_1 ),
    .B1(_0236_),
    .X(_0241_));
 sky130_fd_sc_hd__a211oi_2 _0809_ (.A1(_0235_),
    .A2(_0237_),
    .B1(_0239_),
    .C1(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__xor2_2 _0810_ (.A(_0220_),
    .B(_0221_),
    .X(_0243_));
 sky130_fd_sc_hd__nand3_1 _0811_ (.A(_0219_),
    .B(_0223_),
    .C(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__or4_1 _0812_ (.A(_0229_),
    .B(_0231_),
    .C(_0242_),
    .D(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xnor2_1 _0813_ (.A(\manchester_baby_instance.ram_data_o_11 ),
    .B(\manchester_baby_instance.ram_data_i_11 ),
    .Y(_0246_));
 sky130_fd_sc_hd__and2b_1 _0814_ (.A_N(\manchester_baby_instance.ram_data_o_10 ),
    .B(\manchester_baby_instance.ram_data_i_10 ),
    .X(_0247_));
 sky130_fd_sc_hd__xnor2_1 _0815_ (.A(_0246_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__and2b_1 _0816_ (.A_N(\manchester_baby_instance.ram_data_i_10 ),
    .B(\manchester_baby_instance.ram_data_o_10 ),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(_0247_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__and2b_1 _0818_ (.A_N(\manchester_baby_instance.ram_data_o_9 ),
    .B(\manchester_baby_instance.ram_data_i_9 ),
    .X(_0251_));
 sky130_fd_sc_hd__xnor2_1 _0819_ (.A(_0250_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_1 _0820_ (.A(\manchester_baby_instance.ram_data_o_9 ),
    .B(\manchester_baby_instance.ram_data_i_9 ),
    .Y(_0253_));
 sky130_fd_sc_hd__and2b_1 _0821_ (.A_N(\manchester_baby_instance.ram_data_o_8 ),
    .B(\manchester_baby_instance.ram_data_i_8 ),
    .X(_0254_));
 sky130_fd_sc_hd__or2_1 _0822_ (.A(_0253_),
    .B(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(_0253_),
    .B(_0254_),
    .Y(_0256_));
 sky130_fd_sc_hd__nand2_1 _0824_ (.A(_0255_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_1 _0825_ (.A(\manchester_baby_instance.ram_data_o_8 ),
    .B(\manchester_baby_instance.ram_data_i_8 ),
    .Y(_0258_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(\manchester_baby_instance.ram_data_i_7 ),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _0827_ (.A(\manchester_baby_instance.ram_data_o_7 ),
    .Y(_0260_));
 sky130_fd_sc_hd__a21o_1 _0828_ (.A1(_0260_),
    .A2(\manchester_baby_instance.ram_data_i_7 ),
    .B1(_0258_),
    .X(_0261_));
 sky130_fd_sc_hd__o21a_1 _0829_ (.A1(\manchester_baby_instance.ram_data_o_7 ),
    .A2(_0259_),
    .B1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__or4b_1 _0830_ (.A(_0248_),
    .B(_0252_),
    .C(_0257_),
    .D_N(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__xnor2_1 _0831_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(\manchester_baby_instance.ram_data_o_15 ),
    .Y(_0264_));
 sky130_fd_sc_hd__and2b_1 _0832_ (.A_N(\manchester_baby_instance.ram_data_o_14 ),
    .B(\manchester_baby_instance.ram_data_i_14 ),
    .X(_0265_));
 sky130_fd_sc_hd__xnor2_1 _0833_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__xnor2_1 _0834_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B(\manchester_baby_instance.ram_data_o_14 ),
    .Y(_0267_));
 sky130_fd_sc_hd__and2b_1 _0835_ (.A_N(\manchester_baby_instance.ram_data_o_13 ),
    .B(\manchester_baby_instance.ram_data_i_13 ),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(_0267_),
    .B(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_1 _0837_ (.A(_0267_),
    .B(_0268_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0269_),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__xnor2_1 _0839_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B(\manchester_baby_instance.ram_data_o_13 ),
    .Y(_0272_));
 sky130_fd_sc_hd__and2b_1 _0840_ (.A_N(\manchester_baby_instance.ram_data_o_12 ),
    .B(\manchester_baby_instance.ram_data_i_12 ),
    .X(_0273_));
 sky130_fd_sc_hd__xnor2_1 _0841_ (.A(_0272_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__xor2_1 _0842_ (.A(\manchester_baby_instance.ram_data_o_12 ),
    .B(\manchester_baby_instance.ram_data_i_12 ),
    .X(_0275_));
 sky130_fd_sc_hd__nand2b_1 _0843_ (.A_N(\manchester_baby_instance.ram_data_o_11 ),
    .B(\manchester_baby_instance.ram_data_i_11 ),
    .Y(_0276_));
 sky130_fd_sc_hd__xnor2_1 _0844_ (.A(_0275_),
    .B(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__nor2_1 _0845_ (.A(_0274_),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__or3b_1 _0846_ (.A(_0266_),
    .B(_0271_),
    .C_N(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__a211o_1 _0847_ (.A1(_0228_),
    .A2(_0245_),
    .B1(_0263_),
    .C1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__a21bo_1 _0848_ (.A1(_0255_),
    .A2(_0261_),
    .B1_N(_0256_),
    .X(_0281_));
 sky130_fd_sc_hd__a211o_1 _0849_ (.A1(_0246_),
    .A2(_0247_),
    .B1(_0250_),
    .C1(_0251_),
    .X(_0282_));
 sky130_fd_sc_hd__or2_1 _0850_ (.A(_0246_),
    .B(_0247_),
    .X(_0283_));
 sky130_fd_sc_hd__o311a_1 _0851_ (.A1(_0248_),
    .A2(_0252_),
    .A3(_0281_),
    .B1(_0282_),
    .C1(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a2bb2o_1 _0852_ (.A1_N(_0272_),
    .A2_N(_0273_),
    .B1(_0275_),
    .B2(_0276_),
    .X(_0285_));
 sky130_fd_sc_hd__a21bo_1 _0853_ (.A1(_0272_),
    .A2(_0273_),
    .B1_N(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__a21o_1 _0854_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0269_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _0855_ (.A(_0264_),
    .B(_0265_),
    .X(_0288_));
 sky130_fd_sc_hd__o311a_1 _0856_ (.A1(_0266_),
    .A2(_0271_),
    .A3(_0286_),
    .B1(_0287_),
    .C1(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__o21a_1 _0857_ (.A1(_0279_),
    .A2(_0284_),
    .B1(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__and2b_1 _0858_ (.A_N(\manchester_baby_instance.ram_data_o_22 ),
    .B(\manchester_baby_instance.ram_data_i_22 ),
    .X(_0291_));
 sky130_fd_sc_hd__or2b_1 _0859_ (.A(\manchester_baby_instance.ram_data_o_23 ),
    .B_N(\manchester_baby_instance.ram_data_i_23 ),
    .X(_0292_));
 sky130_fd_sc_hd__or2b_1 _0860_ (.A(\manchester_baby_instance.ram_data_i_23 ),
    .B_N(\manchester_baby_instance.ram_data_o_23 ),
    .X(_0293_));
 sky130_fd_sc_hd__and3_1 _0861_ (.A(_0291_),
    .B(_0292_),
    .C(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _0862_ (.A1(_0292_),
    .A2(_0293_),
    .B1(_0291_),
    .X(_0295_));
 sky130_fd_sc_hd__or2b_1 _0863_ (.A(_0294_),
    .B_N(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__xnor2_1 _0864_ (.A(\manchester_baby_instance.ram_data_o_22 ),
    .B(\manchester_baby_instance.ram_data_i_22 ),
    .Y(_0297_));
 sky130_fd_sc_hd__and2b_1 _0865_ (.A_N(\manchester_baby_instance.ram_data_o_21 ),
    .B(\manchester_baby_instance.ram_data_i_21 ),
    .X(_0298_));
 sky130_fd_sc_hd__or2_1 _0866_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _0867_ (.A(_0297_),
    .B(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _0868_ (.A(_0299_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _0869_ (.A(_0296_),
    .B(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__and2b_1 _0870_ (.A_N(\manchester_baby_instance.ram_data_i_21 ),
    .B(\manchester_baby_instance.ram_data_o_21 ),
    .X(_0303_));
 sky130_fd_sc_hd__nor2_1 _0871_ (.A(_0298_),
    .B(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__and2b_1 _0872_ (.A_N(\manchester_baby_instance.ram_data_o_20 ),
    .B(\manchester_baby_instance.ram_data_i_20 ),
    .X(_0305_));
 sky130_fd_sc_hd__xor2_1 _0873_ (.A(_0304_),
    .B(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__and2b_1 _0874_ (.A_N(\manchester_baby_instance.ram_data_i_20 ),
    .B(\manchester_baby_instance.ram_data_o_20 ),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _0875_ (.A(_0305_),
    .B(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__inv_2 _0876_ (.A(\manchester_baby_instance.ram_data_i_19 ),
    .Y(_0309_));
 sky130_fd_sc_hd__or2_1 _0877_ (.A(\manchester_baby_instance.ram_data_o_19 ),
    .B(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__xor2_1 _0878_ (.A(_0308_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(_0306_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__or2b_1 _0880_ (.A(_0302_),
    .B_N(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _0881_ (.A(\manchester_baby_instance.ram_data_o_19 ),
    .B(_0309_),
    .Y(_0314_));
 sky130_fd_sc_hd__and2b_1 _0882_ (.A_N(\manchester_baby_instance.ram_data_o_18 ),
    .B(\manchester_baby_instance.ram_data_i_18 ),
    .X(_0315_));
 sky130_fd_sc_hd__and3_1 _0883_ (.A(_0310_),
    .B(_0314_),
    .C(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__a21oi_2 _0884_ (.A1(_0310_),
    .A2(_0314_),
    .B1(_0315_),
    .Y(_0317_));
 sky130_fd_sc_hd__xnor2_1 _0885_ (.A(\manchester_baby_instance.ram_data_o_18 ),
    .B(\manchester_baby_instance.ram_data_i_18 ),
    .Y(_0318_));
 sky130_fd_sc_hd__and2b_1 _0886_ (.A_N(\manchester_baby_instance.ram_data_o_17 ),
    .B(\manchester_baby_instance.ram_data_i_17 ),
    .X(_0319_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(_0318_),
    .B(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_1 _0888_ (.A(_0318_),
    .B(_0319_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _0889_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__or3_1 _0890_ (.A(_0316_),
    .B(_0317_),
    .C(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__and2b_1 _0891_ (.A_N(\manchester_baby_instance.ram_data_o_16 ),
    .B(\manchester_baby_instance.ram_data_i_16 ),
    .X(_0324_));
 sky130_fd_sc_hd__xnor2_1 _0892_ (.A(\manchester_baby_instance.ram_data_o_17 ),
    .B(\manchester_baby_instance.ram_data_i_17 ),
    .Y(_0325_));
 sky130_fd_sc_hd__or2_1 _0893_ (.A(_0324_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0894_ (.A(_0324_),
    .B(_0325_),
    .Y(_0327_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(_0326_),
    .B(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__inv_2 _0896_ (.A(\manchester_baby_instance.ram_data_o_15 ),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _0897_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__and2b_1 _0898_ (.A_N(\manchester_baby_instance.ram_data_i_16 ),
    .B(\manchester_baby_instance.ram_data_o_16 ),
    .X(_0331_));
 sky130_fd_sc_hd__nor2_1 _0899_ (.A(_0324_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__xnor2_1 _0900_ (.A(_0330_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _0901_ (.A(_0328_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__or2_1 _0902_ (.A(_0323_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__a211o_1 _0903_ (.A1(_0280_),
    .A2(_0290_),
    .B1(_0313_),
    .C1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _0904_ (.A(_0308_),
    .B(_0310_),
    .Y(_0337_));
 sky130_fd_sc_hd__o21a_1 _0905_ (.A1(_0304_),
    .A2(_0305_),
    .B1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _0906_ (.A1(_0304_),
    .A2(_0305_),
    .B1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__o221a_1 _0907_ (.A1(_0294_),
    .A2(_0299_),
    .B1(_0302_),
    .B2(_0339_),
    .C1(_0295_),
    .X(_0340_));
 sky130_fd_sc_hd__a21o_1 _0908_ (.A1(\manchester_baby_instance.ram_data_i_15 ),
    .A2(_0329_),
    .B1(_0332_),
    .X(_0341_));
 sky130_fd_sc_hd__a21bo_1 _0909_ (.A1(_0326_),
    .A2(_0341_),
    .B1_N(_0327_),
    .X(_0342_));
 sky130_fd_sc_hd__inv_2 _0910_ (.A(_0317_),
    .Y(_0343_));
 sky130_fd_sc_hd__o221a_1 _0911_ (.A1(_0316_),
    .A2(_0320_),
    .B1(_0323_),
    .B2(_0342_),
    .C1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__or2_1 _0912_ (.A(_0313_),
    .B(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__inv_2 _0913_ (.A(\manchester_baby_instance.ram_data_o_24 ),
    .Y(_0346_));
 sky130_fd_sc_hd__and2b_1 _0914_ (.A_N(\manchester_baby_instance.ram_data_o_25 ),
    .B(\manchester_baby_instance.ram_data_i_25 ),
    .X(_0347_));
 sky130_fd_sc_hd__and2b_1 _0915_ (.A_N(\manchester_baby_instance.ram_data_i_25 ),
    .B(\manchester_baby_instance.ram_data_o_25 ),
    .X(_0348_));
 sky130_fd_sc_hd__nor2_1 _0916_ (.A(_0347_),
    .B(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a21o_1 _0917_ (.A1(_0346_),
    .A2(\manchester_baby_instance.ram_data_i_24 ),
    .B1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__and3_1 _0918_ (.A(_0346_),
    .B(\manchester_baby_instance.ram_data_i_24 ),
    .C(_0349_),
    .X(_0351_));
 sky130_fd_sc_hd__inv_2 _0919_ (.A(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0920_ (.A(_0350_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__xnor2_1 _0921_ (.A(\manchester_baby_instance.ram_data_o_24 ),
    .B(\manchester_baby_instance.ram_data_i_24 ),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_2 _0922_ (.A(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _0923_ (.A(_0292_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__or2_1 _0924_ (.A(_0292_),
    .B(_0355_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_1 _0925_ (.A(_0356_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__or2_1 _0926_ (.A(_0353_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__or2b_1 _0927_ (.A(\manchester_baby_instance.ram_data_i_27 ),
    .B_N(\manchester_baby_instance.ram_data_o_27 ),
    .X(_0360_));
 sky130_fd_sc_hd__inv_2 _0928_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .Y(_0361_));
 sky130_fd_sc_hd__o2bb2a_1 _0929_ (.A1_N(_0209_),
    .A2_N(_0360_),
    .B1(\manchester_baby_instance.ram_data_o_26 ),
    .B2(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__and4b_1 _0930_ (.A_N(\manchester_baby_instance.ram_data_o_26 ),
    .B(\manchester_baby_instance.ram_data_i_26 ),
    .C(_0209_),
    .D(_0360_),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _0931_ (.A(_0362_),
    .B(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__xnor2_1 _0932_ (.A(\manchester_baby_instance.ram_data_o_26 ),
    .B(\manchester_baby_instance.ram_data_i_26 ),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _0933_ (.A(_0365_),
    .B(_0347_),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_2 _0934_ (.A(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _0935_ (.A(_0365_),
    .B(_0347_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _0936_ (.A(_0367_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__or2_1 _0937_ (.A(_0364_),
    .B(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__a311o_1 _0938_ (.A1(_0336_),
    .A2(_0340_),
    .A3(_0345_),
    .B1(_0359_),
    .C1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a21o_1 _0939_ (.A1(_0350_),
    .A2(_0356_),
    .B1(_0351_),
    .X(_0372_));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(_0362_),
    .Y(_0373_));
 sky130_fd_sc_hd__o221a_1 _0941_ (.A1(_0363_),
    .A2(_0367_),
    .B1(_0370_),
    .B2(_0372_),
    .C1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nor2_1 _0942_ (.A(_0208_),
    .B(_0209_),
    .Y(_0375_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(_0210_),
    .B(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_2 _0944_ (.A1(_0371_),
    .A2(_0374_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or3_2 _0945_ (.A(\manchester_baby_instance.ram_data_o_28 ),
    .B(_0204_),
    .C(_0206_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _0946_ (.A(_0199_),
    .B(_0202_),
    .Y(_0379_));
 sky130_fd_sc_hd__and2_1 _0947_ (.A(_0203_),
    .B(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__o311ai_4 _0948_ (.A1(_0207_),
    .A2(_0210_),
    .A3(_0377_),
    .B1(_0378_),
    .C1(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_1 _0949_ (.A(\manchester_baby_instance.ram_data_o_31 ),
    .B(\manchester_baby_instance.ram_data_i_31 ),
    .Y(_0382_));
 sky130_fd_sc_hd__xnor2_1 _0950_ (.A(_0200_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0951_ (.A1(_0203_),
    .A2(_0381_),
    .B1(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__or4b_1 _0952_ (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .B(_0187_),
    .C(_0128_),
    .D_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_4 _0953_ (.A(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a31o_1 _0954_ (.A1(_0203_),
    .A2(_0381_),
    .A3(_0383_),
    .B1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__and4bb_2 _0955_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B_N(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .C(_0188_),
    .D(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .X(_0388_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(\manchester_baby_instance.ram_data_i_31 ),
    .Y(_0390_));
 sky130_fd_sc_hd__and4_1 _0958_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B(\manchester_baby_instance.ram_data_i_2 ),
    .C(\manchester_baby_instance.ram_data_i_1 ),
    .D(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_2 _0959_ (.A(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _0960_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(\manchester_baby_instance.ram_data_i_5 ),
    .X(_0393_));
 sky130_fd_sc_hd__and4_1 _0961_ (.A(\manchester_baby_instance.ram_data_i_6 ),
    .B(\manchester_baby_instance.ram_data_i_7 ),
    .C(_0392_),
    .D(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_2 _0962_ (.A(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__and4_1 _0963_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B(\manchester_baby_instance.ram_data_i_9 ),
    .C(\manchester_baby_instance.ram_data_i_10 ),
    .D(\manchester_baby_instance.ram_data_i_11 ),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _0964_ (.A(\manchester_baby_instance.ram_data_i_13 ),
    .B(\manchester_baby_instance.ram_data_i_12 ),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _0965_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(\manchester_baby_instance.ram_data_i_14 ),
    .X(_0398_));
 sky130_fd_sc_hd__and4_1 _0966_ (.A(_0395_),
    .B(_0396_),
    .C(_0397_),
    .D(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__and4_1 _0967_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(\manchester_baby_instance.ram_data_i_17 ),
    .C(\manchester_baby_instance.ram_data_i_18 ),
    .D(\manchester_baby_instance.ram_data_i_19 ),
    .X(_0400_));
 sky130_fd_sc_hd__and4_1 _0968_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B(\manchester_baby_instance.ram_data_i_21 ),
    .C(_0399_),
    .D(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__and3_1 _0969_ (.A(\manchester_baby_instance.ram_data_i_22 ),
    .B(\manchester_baby_instance.ram_data_i_23 ),
    .C(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__and3_1 _0970_ (.A(\manchester_baby_instance.ram_data_i_24 ),
    .B(\manchester_baby_instance.ram_data_i_25 ),
    .C(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _0971_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B(\manchester_baby_instance.ram_data_i_27 ),
    .C(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .B(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0973_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__and4_1 _0974_ (.A(\manchester_baby_instance.ram_data_i_29 ),
    .B(\manchester_baby_instance.ram_data_i_30 ),
    .C(_0390_),
    .D(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a31o_1 _0975_ (.A1(\manchester_baby_instance.ram_data_i_29 ),
    .A2(\manchester_baby_instance.ram_data_i_30 ),
    .A3(_0406_),
    .B1(_0390_),
    .X(_0408_));
 sky130_fd_sc_hd__or3b_1 _0976_ (.A(_0389_),
    .B(_0407_),
    .C_N(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__o21ai_1 _0977_ (.A1(_0384_),
    .A2(_0387_),
    .B1(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__and3b_1 _0978_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .B(_0188_),
    .C(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_4 _0979_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__o21ai_4 _0980_ (.A1(_0412_),
    .A2(_0388_),
    .B1(\manchester_baby_instance.CIRCUIT_0.Acc.tick ),
    .Y(_0413_));
 sky130_fd_sc_hd__clkbuf_4 _0981_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _0982_ (.A0(_0410_),
    .A1(\manchester_baby_instance.ram_data_o_31 ),
    .S(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0983_ (.A(_0415_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_4 _0984_ (.A(_0412_),
    .X(_0416_));
 sky130_fd_sc_hd__o31a_1 _0985_ (.A1(_0207_),
    .A2(_0210_),
    .A3(_0377_),
    .B1(_0378_),
    .X(_0417_));
 sky130_fd_sc_hd__or2_1 _0986_ (.A(_0380_),
    .B(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(\manchester_baby_instance.ram_data_i_29 ),
    .B(_0406_),
    .Y(_0419_));
 sky130_fd_sc_hd__xor2_1 _0988_ (.A(\manchester_baby_instance.ram_data_i_30 ),
    .B(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_4 _0989_ (.A(_0388_),
    .X(_0421_));
 sky130_fd_sc_hd__a32o_1 _0990_ (.A1(_0416_),
    .A2(_0381_),
    .A3(_0418_),
    .B1(_0420_),
    .B2(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(_0422_),
    .A1(\manchester_baby_instance.ram_data_o_30 ),
    .S(_0414_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0992_ (.A(_0423_),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_4 _0993_ (.A(_0412_),
    .X(_0424_));
 sky130_fd_sc_hd__and2b_1 _0994_ (.A_N(_0207_),
    .B(_0378_),
    .X(_0425_));
 sky130_fd_sc_hd__nor2_1 _0995_ (.A(_0210_),
    .B(_0377_),
    .Y(_0426_));
 sky130_fd_sc_hd__xnor2_1 _0996_ (.A(_0425_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__xnor2_1 _0997_ (.A(\manchester_baby_instance.ram_data_i_29 ),
    .B(_0406_),
    .Y(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _0998_ (.A(_0388_),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _0999_ (.A1(_0424_),
    .A2(_0427_),
    .B1(_0428_),
    .B2(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _1000_ (.A0(_0430_),
    .A1(\manchester_baby_instance.ram_data_o_29 ),
    .S(_0414_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _1001_ (.A(_0431_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(\manchester_baby_instance.ram_data_i_28 ),
    .B(_0404_),
    .Y(_0432_));
 sky130_fd_sc_hd__o21ai_1 _1003_ (.A1(_0406_),
    .A2(_0432_),
    .B1(_0421_),
    .Y(_0433_));
 sky130_fd_sc_hd__a311o_1 _1004_ (.A1(_0376_),
    .A2(_0371_),
    .A3(_0374_),
    .B1(_0377_),
    .C1(_0386_),
    .X(_0434_));
 sky130_fd_sc_hd__nand2_1 _1005_ (.A(_0433_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__mux2_1 _1006_ (.A0(_0435_),
    .A1(\manchester_baby_instance.ram_data_o_28 ),
    .S(_0414_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _1007_ (.A(_0436_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _1008_ (.A(_0336_),
    .B(_0340_),
    .C(_0345_),
    .X(_0437_));
 sky130_fd_sc_hd__or2_1 _1009_ (.A(_0437_),
    .B(_0359_),
    .X(_0438_));
 sky130_fd_sc_hd__a21o_1 _1010_ (.A1(_0438_),
    .A2(_0372_),
    .B1(_0369_),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _1011_ (.A1(_0367_),
    .A2(_0439_),
    .B1(_0364_),
    .Y(_0440_));
 sky130_fd_sc_hd__a31o_1 _1012_ (.A1(_0364_),
    .A2(_0367_),
    .A3(_0439_),
    .B1(_0386_),
    .X(_0441_));
 sky130_fd_sc_hd__a21oi_1 _1013_ (.A1(\manchester_baby_instance.ram_data_i_26 ),
    .A2(_0403_),
    .B1(\manchester_baby_instance.ram_data_i_27 ),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_1 _1014_ (.A1(_0404_),
    .A2(_0442_),
    .B1(_0421_),
    .Y(_0443_));
 sky130_fd_sc_hd__o21ai_1 _1015_ (.A1(_0440_),
    .A2(_0441_),
    .B1(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(_0444_),
    .A1(\manchester_baby_instance.ram_data_o_27 ),
    .S(_0414_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0445_),
    .X(_0074_));
 sky130_fd_sc_hd__nand3_1 _1018_ (.A(_0369_),
    .B(_0438_),
    .C(_0372_),
    .Y(_0446_));
 sky130_fd_sc_hd__xnor2_1 _1019_ (.A(\manchester_baby_instance.ram_data_i_26 ),
    .B(_0403_),
    .Y(_0447_));
 sky130_fd_sc_hd__a32o_1 _1020_ (.A1(_0416_),
    .A2(_0439_),
    .A3(_0446_),
    .B1(_0447_),
    .B2(_0421_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(_0448_),
    .A1(\manchester_baby_instance.ram_data_o_26 ),
    .S(_0414_),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(_0449_),
    .X(_0073_));
 sky130_fd_sc_hd__or2_1 _1023_ (.A(_0437_),
    .B(_0358_),
    .X(_0450_));
 sky130_fd_sc_hd__a21oi_1 _1024_ (.A1(_0356_),
    .A2(_0450_),
    .B1(_0353_),
    .Y(_0451_));
 sky130_fd_sc_hd__a31o_1 _1025_ (.A1(_0353_),
    .A2(_0356_),
    .A3(_0450_),
    .B1(_0386_),
    .X(_0452_));
 sky130_fd_sc_hd__a21oi_1 _1026_ (.A1(\manchester_baby_instance.ram_data_i_24 ),
    .A2(_0402_),
    .B1(\manchester_baby_instance.ram_data_i_25 ),
    .Y(_0453_));
 sky130_fd_sc_hd__o21ai_1 _1027_ (.A1(_0403_),
    .A2(_0453_),
    .B1(_0421_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21ai_1 _1028_ (.A1(_0451_),
    .A2(_0452_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(_0455_),
    .A1(\manchester_baby_instance.ram_data_o_25 ),
    .S(_0414_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _1030_ (.A(_0456_),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _1031_ (.A(_0437_),
    .B(_0358_),
    .Y(_0457_));
 sky130_fd_sc_hd__xnor2_1 _1032_ (.A(\manchester_baby_instance.ram_data_i_24 ),
    .B(_0402_),
    .Y(_0458_));
 sky130_fd_sc_hd__a32o_1 _1033_ (.A1(_0416_),
    .A2(_0450_),
    .A3(_0457_),
    .B1(_0458_),
    .B2(_0421_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(_0459_),
    .A1(\manchester_baby_instance.ram_data_o_24 ),
    .S(_0414_),
    .X(_0460_));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(_0460_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _1036_ (.A(_0280_),
    .B(_0290_),
    .X(_0461_));
 sky130_fd_sc_hd__o21ai_1 _1037_ (.A1(_0461_),
    .A2(_0335_),
    .B1(_0344_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _1038_ (.A(_0312_),
    .B(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__a21o_1 _1039_ (.A1(_0339_),
    .A2(_0463_),
    .B1(_0301_),
    .X(_0464_));
 sky130_fd_sc_hd__a21oi_1 _1040_ (.A1(_0299_),
    .A2(_0464_),
    .B1(_0296_),
    .Y(_0465_));
 sky130_fd_sc_hd__a31o_1 _1041_ (.A1(_0296_),
    .A2(_0299_),
    .A3(_0464_),
    .B1(_0386_),
    .X(_0466_));
 sky130_fd_sc_hd__a21oi_1 _1042_ (.A1(\manchester_baby_instance.ram_data_i_22 ),
    .A2(_0401_),
    .B1(\manchester_baby_instance.ram_data_i_23 ),
    .Y(_0467_));
 sky130_fd_sc_hd__o21ai_1 _1043_ (.A1(_0402_),
    .A2(_0467_),
    .B1(_0421_),
    .Y(_0468_));
 sky130_fd_sc_hd__o21ai_1 _1044_ (.A1(_0465_),
    .A2(_0466_),
    .B1(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _1045_ (.A(_0413_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(_0469_),
    .A1(\manchester_baby_instance.ram_data_o_23 ),
    .S(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _1047_ (.A(_0471_),
    .X(_0070_));
 sky130_fd_sc_hd__nand3_1 _1048_ (.A(_0301_),
    .B(_0339_),
    .C(_0463_),
    .Y(_0472_));
 sky130_fd_sc_hd__xnor2_1 _1049_ (.A(\manchester_baby_instance.ram_data_i_22 ),
    .B(_0401_),
    .Y(_0473_));
 sky130_fd_sc_hd__a32o_1 _1050_ (.A1(_0416_),
    .A2(_0464_),
    .A3(_0472_),
    .B1(_0473_),
    .B2(_0421_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1051_ (.A0(_0474_),
    .A1(\manchester_baby_instance.ram_data_o_22 ),
    .S(_0470_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _1052_ (.A(_0475_),
    .X(_0069_));
 sky130_fd_sc_hd__nand2_1 _1053_ (.A(_0311_),
    .B(_0462_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _1054_ (.A(_0337_),
    .B(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__xor2_1 _1055_ (.A(_0306_),
    .B(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__and2_1 _1056_ (.A(_0395_),
    .B(_0396_),
    .X(_0479_));
 sky130_fd_sc_hd__and4_1 _1057_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B(\manchester_baby_instance.ram_data_i_13 ),
    .C(\manchester_baby_instance.ram_data_i_12 ),
    .D(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__and4_1 _1058_ (.A(\manchester_baby_instance.ram_data_i_15 ),
    .B(\manchester_baby_instance.ram_data_i_16 ),
    .C(\manchester_baby_instance.ram_data_i_17 ),
    .D(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _1059_ (.A(\manchester_baby_instance.ram_data_i_18 ),
    .B(\manchester_baby_instance.ram_data_i_19 ),
    .C(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__a21oi_1 _1060_ (.A1(\manchester_baby_instance.ram_data_i_20 ),
    .A2(_0482_),
    .B1(\manchester_baby_instance.ram_data_i_21 ),
    .Y(_0483_));
 sky130_fd_sc_hd__clkbuf_4 _1061_ (.A(_0388_),
    .X(_0484_));
 sky130_fd_sc_hd__o21a_1 _1062_ (.A1(_0401_),
    .A2(_0483_),
    .B1(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__a21o_1 _1063_ (.A1(_0424_),
    .A2(_0478_),
    .B1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(_0486_),
    .A1(\manchester_baby_instance.ram_data_o_21 ),
    .S(_0470_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _1065_ (.A(_0487_),
    .X(_0068_));
 sky130_fd_sc_hd__or2_1 _1066_ (.A(_0311_),
    .B(_0462_),
    .X(_0488_));
 sky130_fd_sc_hd__xnor2_1 _1067_ (.A(\manchester_baby_instance.ram_data_i_20 ),
    .B(_0482_),
    .Y(_0489_));
 sky130_fd_sc_hd__a32o_1 _1068_ (.A1(_0416_),
    .A2(_0476_),
    .A3(_0488_),
    .B1(_0489_),
    .B2(_0429_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1069_ (.A0(_0490_),
    .A1(\manchester_baby_instance.ram_data_o_20 ),
    .S(_0470_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_1 _1070_ (.A(_0491_),
    .X(_0067_));
 sky130_fd_sc_hd__or2_1 _1071_ (.A(_0461_),
    .B(_0334_),
    .X(_0492_));
 sky130_fd_sc_hd__a21o_1 _1072_ (.A1(_0342_),
    .A2(_0492_),
    .B1(_0322_),
    .X(_0493_));
 sky130_fd_sc_hd__a211o_1 _1073_ (.A1(_0320_),
    .A2(_0493_),
    .B1(_0316_),
    .C1(_0317_),
    .X(_0494_));
 sky130_fd_sc_hd__o211ai_1 _1074_ (.A1(_0316_),
    .A2(_0317_),
    .B1(_0320_),
    .C1(_0493_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(\manchester_baby_instance.ram_data_i_18 ),
    .B(_0481_),
    .Y(_0496_));
 sky130_fd_sc_hd__a21o_1 _1076_ (.A1(_0309_),
    .A2(_0496_),
    .B1(_0482_),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _1077_ (.A1(_0412_),
    .A2(_0494_),
    .A3(_0495_),
    .B1(_0497_),
    .B2(_0429_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1078_ (.A0(_0498_),
    .A1(\manchester_baby_instance.ram_data_o_19 ),
    .S(_0470_),
    .X(_0499_));
 sky130_fd_sc_hd__clkbuf_1 _1079_ (.A(_0499_),
    .X(_0066_));
 sky130_fd_sc_hd__nand3_1 _1080_ (.A(_0322_),
    .B(_0342_),
    .C(_0492_),
    .Y(_0500_));
 sky130_fd_sc_hd__and2_1 _1081_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(_0399_),
    .X(_0501_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(\manchester_baby_instance.ram_data_i_17 ),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__xor2_1 _1083_ (.A(\manchester_baby_instance.ram_data_i_18 ),
    .B(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a32o_1 _1084_ (.A1(_0412_),
    .A2(_0493_),
    .A3(_0500_),
    .B1(_0503_),
    .B2(_0429_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1085_ (.A0(_0504_),
    .A1(\manchester_baby_instance.ram_data_o_18 ),
    .S(_0470_),
    .X(_0505_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0505_),
    .X(_0065_));
 sky130_fd_sc_hd__nand2_1 _1087_ (.A(_0280_),
    .B(_0290_),
    .Y(_0506_));
 sky130_fd_sc_hd__a21bo_1 _1088_ (.A1(_0506_),
    .A2(_0333_),
    .B1_N(_0341_),
    .X(_0507_));
 sky130_fd_sc_hd__xor2_1 _1089_ (.A(_0328_),
    .B(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__or2_1 _1090_ (.A(\manchester_baby_instance.ram_data_i_17 ),
    .B(_0501_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _1091_ (.A(_0502_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__a22o_1 _1092_ (.A1(_0416_),
    .A2(_0508_),
    .B1(_0510_),
    .B2(_0429_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _1093_ (.A0(_0511_),
    .A1(\manchester_baby_instance.ram_data_o_17 ),
    .S(_0470_),
    .X(_0512_));
 sky130_fd_sc_hd__clkbuf_1 _1094_ (.A(_0512_),
    .X(_0064_));
 sky130_fd_sc_hd__xnor2_1 _1095_ (.A(\manchester_baby_instance.ram_data_i_16 ),
    .B(_0399_),
    .Y(_0513_));
 sky130_fd_sc_hd__xnor2_1 _1096_ (.A(_0461_),
    .B(_0333_),
    .Y(_0514_));
 sky130_fd_sc_hd__a22o_1 _1097_ (.A1(_0484_),
    .A2(_0513_),
    .B1(_0514_),
    .B2(_0424_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1098_ (.A0(_0515_),
    .A1(\manchester_baby_instance.ram_data_o_16 ),
    .S(_0470_),
    .X(_0516_));
 sky130_fd_sc_hd__clkbuf_1 _1099_ (.A(_0516_),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_1 _1100_ (.A1(_0228_),
    .A2(_0245_),
    .B1(_0263_),
    .X(_0517_));
 sky130_fd_sc_hd__nand2_1 _1101_ (.A(_0517_),
    .B(_0284_),
    .Y(_0518_));
 sky130_fd_sc_hd__a21boi_1 _1102_ (.A1(_0278_),
    .A2(_0518_),
    .B1_N(_0286_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_1 _1103_ (.A1(_0271_),
    .A2(_0519_),
    .B1(_0269_),
    .Y(_0520_));
 sky130_fd_sc_hd__xnor2_1 _1104_ (.A(_0266_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__and3_1 _1105_ (.A(_0395_),
    .B(_0396_),
    .C(_0397_),
    .X(_0522_));
 sky130_fd_sc_hd__a21oi_1 _1106_ (.A1(\manchester_baby_instance.ram_data_i_14 ),
    .A2(_0522_),
    .B1(\manchester_baby_instance.ram_data_i_15 ),
    .Y(_0523_));
 sky130_fd_sc_hd__o21a_1 _1107_ (.A1(_0399_),
    .A2(_0523_),
    .B1(_0484_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _1108_ (.A1(_0424_),
    .A2(_0521_),
    .B1(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _1109_ (.A0(_0525_),
    .A1(\manchester_baby_instance.ram_data_o_15 ),
    .S(_0470_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1110_ (.A(_0526_),
    .X(_0062_));
 sky130_fd_sc_hd__xnor2_1 _1111_ (.A(\manchester_baby_instance.ram_data_i_14 ),
    .B(_0522_),
    .Y(_0527_));
 sky130_fd_sc_hd__xor2_1 _1112_ (.A(_0271_),
    .B(_0519_),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _1113_ (.A1(_0484_),
    .A2(_0527_),
    .B1(_0528_),
    .B2(_0424_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _1114_ (.A0(_0529_),
    .A1(\manchester_baby_instance.ram_data_o_14 ),
    .S(_0470_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1115_ (.A(_0530_),
    .X(_0061_));
 sky130_fd_sc_hd__nand2_1 _1116_ (.A(_0275_),
    .B(_0276_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21o_1 _1117_ (.A1(_0517_),
    .A2(_0284_),
    .B1(_0277_),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1118_ (.A1(_0531_),
    .A2(_0532_),
    .B1(_0274_),
    .Y(_0533_));
 sky130_fd_sc_hd__a31o_1 _1119_ (.A1(_0274_),
    .A2(_0531_),
    .A3(_0532_),
    .B1(_0386_),
    .X(_0534_));
 sky130_fd_sc_hd__a21oi_1 _1120_ (.A1(\manchester_baby_instance.ram_data_i_12 ),
    .A2(_0479_),
    .B1(\manchester_baby_instance.ram_data_i_13 ),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_1 _1121_ (.A1(_0522_),
    .A2(_0535_),
    .B1(_0421_),
    .Y(_0536_));
 sky130_fd_sc_hd__o21ai_1 _1122_ (.A1(_0533_),
    .A2(_0534_),
    .B1(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__clkbuf_4 _1123_ (.A(_0413_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _1124_ (.A0(_0537_),
    .A1(\manchester_baby_instance.ram_data_o_13 ),
    .S(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1125_ (.A(_0539_),
    .X(_0060_));
 sky130_fd_sc_hd__xnor2_1 _1126_ (.A(\manchester_baby_instance.ram_data_i_12 ),
    .B(_0479_),
    .Y(_0540_));
 sky130_fd_sc_hd__xnor2_1 _1127_ (.A(_0277_),
    .B(_0518_),
    .Y(_0541_));
 sky130_fd_sc_hd__a22o_1 _1128_ (.A1(_0484_),
    .A2(_0540_),
    .B1(_0541_),
    .B2(_0424_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _1129_ (.A0(_0542_),
    .A1(\manchester_baby_instance.ram_data_o_12 ),
    .S(_0538_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1130_ (.A(_0543_),
    .X(_0059_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(_0228_),
    .B(_0245_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand3b_1 _1132_ (.A_N(_0257_),
    .B(_0262_),
    .C(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a21oi_1 _1133_ (.A1(_0281_),
    .A2(_0545_),
    .B1(_0252_),
    .Y(_0546_));
 sky130_fd_sc_hd__o21ba_1 _1134_ (.A1(_0250_),
    .A2(_0251_),
    .B1_N(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__xor2_1 _1135_ (.A(_0248_),
    .B(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__and3_1 _1136_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B(\manchester_baby_instance.ram_data_i_9 ),
    .C(_0395_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(\manchester_baby_instance.ram_data_i_10 ),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__xor2_1 _1138_ (.A(\manchester_baby_instance.ram_data_i_11 ),
    .B(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _1139_ (.A1(_0416_),
    .A2(_0548_),
    .B1(_0551_),
    .B2(_0429_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _1140_ (.A0(_0552_),
    .A1(\manchester_baby_instance.ram_data_o_11 ),
    .S(_0538_),
    .X(_0553_));
 sky130_fd_sc_hd__clkbuf_1 _1141_ (.A(_0553_),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _1142_ (.A(\manchester_baby_instance.ram_data_i_10 ),
    .B(_0549_),
    .X(_0554_));
 sky130_fd_sc_hd__nand2_1 _1143_ (.A(_0550_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__and3_1 _1144_ (.A(_0252_),
    .B(_0281_),
    .C(_0545_),
    .X(_0556_));
 sky130_fd_sc_hd__nor2_1 _1145_ (.A(_0546_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a22o_1 _1146_ (.A1(_0484_),
    .A2(_0555_),
    .B1(_0557_),
    .B2(_0424_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _1147_ (.A0(_0558_),
    .A1(\manchester_baby_instance.ram_data_o_10 ),
    .S(_0538_),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_1 _1148_ (.A(_0559_),
    .X(_0057_));
 sky130_fd_sc_hd__a21bo_1 _1149_ (.A1(_0544_),
    .A2(_0262_),
    .B1_N(_0261_),
    .X(_0560_));
 sky130_fd_sc_hd__xnor2_1 _1150_ (.A(_0257_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _1151_ (.A1(\manchester_baby_instance.ram_data_i_8 ),
    .A2(_0395_),
    .B1(\manchester_baby_instance.ram_data_i_9 ),
    .Y(_0562_));
 sky130_fd_sc_hd__or2_1 _1152_ (.A(_0549_),
    .B(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _1153_ (.A1(_0416_),
    .A2(_0561_),
    .B1(_0563_),
    .B2(_0429_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(_0564_),
    .A1(\manchester_baby_instance.ram_data_o_9 ),
    .S(_0538_),
    .X(_0565_));
 sky130_fd_sc_hd__clkbuf_1 _1155_ (.A(_0565_),
    .X(_0056_));
 sky130_fd_sc_hd__xnor2_1 _1156_ (.A(\manchester_baby_instance.ram_data_i_8 ),
    .B(_0395_),
    .Y(_0566_));
 sky130_fd_sc_hd__xor2_1 _1157_ (.A(_0544_),
    .B(_0262_),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _1158_ (.A1(_0484_),
    .A2(_0566_),
    .B1(_0567_),
    .B2(_0424_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_1 _1159_ (.A0(_0568_),
    .A1(\manchester_baby_instance.ram_data_o_8 ),
    .S(_0538_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_1 _1160_ (.A(_0569_),
    .X(_0055_));
 sky130_fd_sc_hd__o31ai_1 _1161_ (.A1(_0231_),
    .A2(_0242_),
    .A3(_0244_),
    .B1(_0224_),
    .Y(_0570_));
 sky130_fd_sc_hd__or2b_1 _1162_ (.A(_0216_),
    .B_N(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__a21oi_1 _1163_ (.A1(_0225_),
    .A2(_0571_),
    .B1(_0213_),
    .Y(_0572_));
 sky130_fd_sc_hd__a31o_1 _1164_ (.A1(_0213_),
    .A2(_0225_),
    .A3(_0571_),
    .B1(_0386_),
    .X(_0573_));
 sky130_fd_sc_hd__a31o_1 _1165_ (.A1(\manchester_baby_instance.ram_data_i_6 ),
    .A2(_0392_),
    .A3(_0393_),
    .B1(\manchester_baby_instance.ram_data_i_7 ),
    .X(_0574_));
 sky130_fd_sc_hd__or2b_1 _1166_ (.A(_0395_),
    .B_N(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__a2bb2o_1 _1167_ (.A1_N(_0572_),
    .A2_N(_0573_),
    .B1(_0575_),
    .B2(_0484_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(_0576_),
    .A1(\manchester_baby_instance.ram_data_o_7 ),
    .S(_0538_),
    .X(_0577_));
 sky130_fd_sc_hd__clkbuf_1 _1169_ (.A(_0577_),
    .X(_0054_));
 sky130_fd_sc_hd__and2_1 _1170_ (.A(_0392_),
    .B(_0393_),
    .X(_0578_));
 sky130_fd_sc_hd__xnor2_1 _1171_ (.A(\manchester_baby_instance.ram_data_i_6 ),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__xnor2_1 _1172_ (.A(_0216_),
    .B(_0570_),
    .Y(_0580_));
 sky130_fd_sc_hd__a22o_1 _1173_ (.A1(_0484_),
    .A2(_0579_),
    .B1(_0580_),
    .B2(_0424_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(_0581_),
    .A1(\manchester_baby_instance.ram_data_o_6 ),
    .S(_0538_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_1 _1175_ (.A(_0582_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _1176_ (.A(_0219_),
    .B(_0223_),
    .Y(_0583_));
 sky130_fd_sc_hd__nor2_1 _1177_ (.A(_0231_),
    .B(_0242_),
    .Y(_0584_));
 sky130_fd_sc_hd__a21bo_1 _1178_ (.A1(_0584_),
    .A2(_0243_),
    .B1_N(_0222_),
    .X(_0585_));
 sky130_fd_sc_hd__xnor2_1 _1179_ (.A(_0583_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__a21oi_1 _1180_ (.A1(\manchester_baby_instance.ram_data_i_4 ),
    .A2(_0392_),
    .B1(\manchester_baby_instance.ram_data_i_5 ),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _1181_ (.A(_0578_),
    .B(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _1182_ (.A1(_0416_),
    .A2(_0586_),
    .B1(_0588_),
    .B2(_0429_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _1183_ (.A0(_0589_),
    .A1(\manchester_baby_instance.ram_data_o_5 ),
    .S(_0538_),
    .X(_0590_));
 sky130_fd_sc_hd__clkbuf_1 _1184_ (.A(_0590_),
    .X(_0052_));
 sky130_fd_sc_hd__xor2_1 _1185_ (.A(_0584_),
    .B(_0243_),
    .X(_0591_));
 sky130_fd_sc_hd__xnor2_1 _1186_ (.A(\manchester_baby_instance.ram_data_i_4 ),
    .B(_0392_),
    .Y(_0592_));
 sky130_fd_sc_hd__a22o_1 _1187_ (.A1(_0416_),
    .A2(_0591_),
    .B1(_0592_),
    .B2(_0484_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(_0593_),
    .A1(\manchester_baby_instance.ram_data_o_4 ),
    .S(_0538_),
    .X(_0594_));
 sky130_fd_sc_hd__clkbuf_1 _1189_ (.A(_0594_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _1190_ (.A1(_0235_),
    .A2(_0237_),
    .B1(_0241_),
    .X(_0595_));
 sky130_fd_sc_hd__nor2_1 _1191_ (.A(_0231_),
    .B(_0239_),
    .Y(_0596_));
 sky130_fd_sc_hd__xnor2_1 _1192_ (.A(_0595_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__and3_1 _1193_ (.A(_0132_),
    .B(_0134_),
    .C(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _1194_ (.A(\manchester_baby_instance.ram_data_i_3 ),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_1 _1195_ (.A1(_0392_),
    .A2(_0599_),
    .B1(_0421_),
    .Y(_0600_));
 sky130_fd_sc_hd__o21ai_1 _1196_ (.A1(_0386_),
    .A2(_0597_),
    .B1(_0600_),
    .Y(_0601_));
 sky130_fd_sc_hd__mux2_1 _1197_ (.A0(_0601_),
    .A1(\manchester_baby_instance.ram_data_o_3 ),
    .S(_0413_),
    .X(_0602_));
 sky130_fd_sc_hd__clkbuf_1 _1198_ (.A(_0602_),
    .X(_0050_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(_0235_),
    .B(_0237_),
    .Y(_0603_));
 sky130_fd_sc_hd__or2_1 _1200_ (.A(_0235_),
    .B(_0237_),
    .X(_0604_));
 sky130_fd_sc_hd__a21oi_1 _1201_ (.A1(_0134_),
    .A2(\manchester_baby_instance.ram_data_i_0 ),
    .B1(_0132_),
    .Y(_0605_));
 sky130_fd_sc_hd__or2_1 _1202_ (.A(_0598_),
    .B(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__a32o_1 _1203_ (.A1(_0412_),
    .A2(_0603_),
    .A3(_0604_),
    .B1(_0606_),
    .B2(_0429_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _1204_ (.A0(_0607_),
    .A1(\manchester_baby_instance.ram_data_o_2 ),
    .S(_0413_),
    .X(_0608_));
 sky130_fd_sc_hd__clkbuf_1 _1205_ (.A(_0608_),
    .X(_0049_));
 sky130_fd_sc_hd__inv_2 _1206_ (.A(_0235_),
    .Y(_0609_));
 sky130_fd_sc_hd__or4_1 _1207_ (.A(_0232_),
    .B(\manchester_baby_instance.ram_data_o_0 ),
    .C(_0233_),
    .D(_0234_),
    .X(_0610_));
 sky130_fd_sc_hd__xnor2_1 _1208_ (.A(_0134_),
    .B(\manchester_baby_instance.ram_data_i_0 ),
    .Y(_0611_));
 sky130_fd_sc_hd__a32o_1 _1209_ (.A1(_0412_),
    .A2(_0609_),
    .A3(_0610_),
    .B1(_0611_),
    .B2(_0429_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(_0612_),
    .A1(\manchester_baby_instance.ram_data_o_1 ),
    .S(_0413_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_1 _1211_ (.A(_0613_),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _1212_ (.A1(_0232_),
    .A2(_0424_),
    .B1(_0414_),
    .X(_0614_));
 sky130_fd_sc_hd__a21oi_1 _1213_ (.A1(\manchester_baby_instance.ram_data_o_0 ),
    .A2(_0389_),
    .B1(_0414_),
    .Y(_0615_));
 sky130_fd_sc_hd__a22o_1 _1214_ (.A1(net69),
    .A2(_0614_),
    .B1(_0615_),
    .B2(\manchester_baby_instance.ram_data_i_0 ),
    .X(_0047_));
 sky130_fd_sc_hd__inv_2 _1215_ (.A(net59),
    .Y(_0616_));
 sky130_fd_sc_hd__or4_4 _1216_ (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .C(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .D(\manchester_baby_instance.BASE_0.s_countReg[3] ),
    .X(_0617_));
 sky130_fd_sc_hd__or4_4 _1217_ (.A(\manchester_baby_instance.BASE_0.s_countReg[4] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[5] ),
    .C(\manchester_baby_instance.BASE_0.s_countReg[6] ),
    .D(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__or4_4 _1218_ (.A(\manchester_baby_instance.BASE_0.s_countReg[7] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[8] ),
    .C(net49),
    .D(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__or4_4 _1219_ (.A(\manchester_baby_instance.BASE_0.s_countReg[10] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[11] ),
    .C(net29),
    .D(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__or4_4 _1220_ (.A(\manchester_baby_instance.BASE_0.s_countReg[13] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[14] ),
    .C(\manchester_baby_instance.BASE_0.s_countReg[15] ),
    .D(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__buf_6 _1221_ (.A(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__or2_1 _1222_ (.A(\manchester_baby_instance.BASE_0.s_countReg[16] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[17] ),
    .X(_0623_));
 sky130_fd_sc_hd__or4_4 _1223_ (.A(\manchester_baby_instance.BASE_0.s_countReg[18] ),
    .B(net38),
    .C(_0622_),
    .D(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or3_4 _1224_ (.A(\manchester_baby_instance.BASE_0.s_countReg[20] ),
    .B(net21),
    .C(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__or2_4 _1225_ (.A(_0625_),
    .B(\manchester_baby_instance.BASE_0.s_countReg[22] ),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_4 _1226_ (.A(net76),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_2 _1227_ (.A(_0616_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__or2_1 _1228_ (.A(\manchester_baby_instance.BASE_0.s_countReg[25] ),
    .B(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__buf_6 _1229_ (.A(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__inv_4 _1230_ (.A(_0630_),
    .Y(\manchester_baby_instance.BASE_0.s_tickNext ));
 sky130_fd_sc_hd__nand2_1 _1231_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .Y(_0631_));
 sky130_fd_sc_hd__nor2_1 _1232_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__and4b_1 _1233_ (.A_N(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ),
    .B(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ),
    .C(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_1 _1234_ (.A(_0633_),
    .X(net7));
 sky130_fd_sc_hd__and2b_1 _1235_ (.A_N(net18),
    .B(net19),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_1 _1236_ (.A(_0634_),
    .X(_0000_));
 sky130_fd_sc_hd__and2b_1 _1237_ (.A_N(net8),
    .B(\manchester_baby_instance.CIRCUIT_0.GATES_13.input1 ),
    .X(_0635_));
 sky130_fd_sc_hd__clkbuf_1 _1238_ (.A(_0635_),
    .X(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ));
 sky130_fd_sc_hd__and3b_1 _1239_ (.A_N(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ),
    .B(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ),
    .C(_0187_),
    .X(_0636_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1240_ (.A(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__a22o_1 _1241_ (.A1(_0125_),
    .A2(_0188_),
    .B1(_0632_),
    .B2(_0127_),
    .X(_0638_));
 sky130_fd_sc_hd__a22o_1 _1242_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net2));
 sky130_fd_sc_hd__a22o_1 _1243_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net3));
 sky130_fd_sc_hd__a22o_1 _1244_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net4));
 sky130_fd_sc_hd__a22o_1 _1245_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net5));
 sky130_fd_sc_hd__a22o_1 _1246_ (.A1(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .A2(_0637_),
    .B1(_0638_),
    .B2(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net6));
 sky130_fd_sc_hd__buf_4 _1247_ (.A(net1),
    .X(_0639_));
 sky130_fd_sc_hd__buf_4 _1248_ (.A(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__inv_2 _1249_ (.A(_0640_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1250_ (.A(_0640_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(_0640_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1252_ (.A(_0640_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1253_ (.A(_0640_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1254_ (.A(_0640_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1255_ (.A(_0640_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1256_ (.A(_0640_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1257_ (.A(_0640_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1258_ (.A(_0640_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_4 _1259_ (.A(_0639_),
    .X(_0641_));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(_0641_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1261_ (.A(_0641_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1262_ (.A(_0641_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1263_ (.A(_0641_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1264_ (.A(_0641_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1265_ (.A(_0641_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1266_ (.A(_0641_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1267_ (.A(_0641_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1268_ (.A(_0641_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1269_ (.A(_0641_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_4 _1270_ (.A(_0639_),
    .X(_0642_));
 sky130_fd_sc_hd__inv_2 _1271_ (.A(_0642_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1272_ (.A(_0642_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1273_ (.A(_0642_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1274_ (.A(_0642_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1275_ (.A(_0642_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1276_ (.A(_0642_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1277_ (.A(_0642_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1278_ (.A(_0642_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(_0642_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1280_ (.A(_0642_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_4 _1281_ (.A(_0639_),
    .X(_0643_));
 sky130_fd_sc_hd__inv_2 _1282_ (.A(_0643_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1283_ (.A(_0643_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1284_ (.A(_0643_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1285_ (.A(_0643_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(_0643_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1287_ (.A(_0643_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(_0643_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1289_ (.A(_0643_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1290_ (.A(_0643_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1291_ (.A(_0643_),
    .Y(_0040_));
 sky130_fd_sc_hd__or2b_1 _1292_ (.A(net55),
    .B_N(\manchester_baby_instance.BASE_0.s_tickReg ),
    .X(_0644_));
 sky130_fd_sc_hd__xnor2_1 _1293_ (.A(net19),
    .B(net56),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1294_ (.A(_0639_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(_0128_),
    .B(_0631_),
    .Y(_0090_));
 sky130_fd_sc_hd__and2_1 _1296_ (.A(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ),
    .B(_0128_),
    .X(_0645_));
 sky130_fd_sc_hd__or2_1 _1297_ (.A(_0129_),
    .B(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_1 _1298_ (.A(_0646_),
    .X(_0091_));
 sky130_fd_sc_hd__and2b_1 _1299_ (.A_N(net63),
    .B(net55),
    .X(_0647_));
 sky130_fd_sc_hd__clkbuf_1 _1300_ (.A(_0647_),
    .X(_0092_));
 sky130_fd_sc_hd__inv_2 _1301_ (.A(net20),
    .Y(_0093_));
 sky130_fd_sc_hd__xnor2_1 _1302_ (.A(net17),
    .B(net61),
    .Y(_0094_));
 sky130_fd_sc_hd__or3_1 _1303_ (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .B(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .C(net44),
    .X(_0648_));
 sky130_fd_sc_hd__o21ai_1 _1304_ (.A1(net20),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .B1(net44),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _1305_ (.A(_0648_),
    .B(net45),
    .Y(_0095_));
 sky130_fd_sc_hd__nand2_1 _1306_ (.A(\manchester_baby_instance.BASE_0.s_countReg[3] ),
    .B(_0648_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _1307_ (.A(_0617_),
    .B(net24),
    .Y(_0096_));
 sky130_fd_sc_hd__or2_1 _1308_ (.A(\manchester_baby_instance.BASE_0.s_countReg[4] ),
    .B(_0617_),
    .X(_0651_));
 sky130_fd_sc_hd__nand2_1 _1309_ (.A(net42),
    .B(_0617_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _1310_ (.A(_0651_),
    .B(net43),
    .Y(_0097_));
 sky130_fd_sc_hd__xnor2_1 _1311_ (.A(\manchester_baby_instance.BASE_0.s_countReg[5] ),
    .B(_0651_),
    .Y(_0098_));
 sky130_fd_sc_hd__o21ai_1 _1312_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[5] ),
    .A2(_0651_),
    .B1(\manchester_baby_instance.BASE_0.s_countReg[6] ),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _1313_ (.A(_0618_),
    .B(net27),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(\manchester_baby_instance.BASE_0.s_countReg[7] ),
    .B(_0618_),
    .Y(_0654_));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(\manchester_baby_instance.BASE_0.s_countReg[7] ),
    .B(_0618_),
    .X(_0655_));
 sky130_fd_sc_hd__o21a_1 _1316_ (.A1(_0654_),
    .A2(_0655_),
    .B1(_0630_),
    .X(_0100_));
 sky130_fd_sc_hd__xnor2_1 _1317_ (.A(\manchester_baby_instance.BASE_0.s_countReg[8] ),
    .B(_0654_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _1318_ (.A(\manchester_baby_instance.BASE_0.s_tickNext ),
    .B(net67),
    .Y(_0101_));
 sky130_fd_sc_hd__o31ai_1 _1319_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[7] ),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[8] ),
    .A3(_0618_),
    .B1(net49),
    .Y(_0657_));
 sky130_fd_sc_hd__a21oi_1 _1320_ (.A1(_0619_),
    .A2(net50),
    .B1(\manchester_baby_instance.BASE_0.s_tickNext ),
    .Y(_0102_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(\manchester_baby_instance.BASE_0.s_countReg[10] ),
    .B(_0619_),
    .Y(_0658_));
 sky130_fd_sc_hd__and2_1 _1322_ (.A(\manchester_baby_instance.BASE_0.s_countReg[10] ),
    .B(_0619_),
    .X(_0659_));
 sky130_fd_sc_hd__o21a_1 _1323_ (.A1(_0658_),
    .A2(_0659_),
    .B1(_0630_),
    .X(_0103_));
 sky130_fd_sc_hd__xnor2_1 _1324_ (.A(\manchester_baby_instance.BASE_0.s_countReg[11] ),
    .B(_0658_),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_1 _1325_ (.A(\manchester_baby_instance.BASE_0.s_tickNext ),
    .B(net65),
    .Y(_0104_));
 sky130_fd_sc_hd__o31ai_1 _1326_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[10] ),
    .A2(\manchester_baby_instance.BASE_0.s_countReg[11] ),
    .A3(_0619_),
    .B1(net29),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(_0620_),
    .B(net30),
    .Y(_0105_));
 sky130_fd_sc_hd__or2_1 _1328_ (.A(\manchester_baby_instance.BASE_0.s_countReg[13] ),
    .B(_0620_),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _1329_ (.A(\manchester_baby_instance.BASE_0.s_countReg[13] ),
    .B(_0620_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _1330_ (.A(_0662_),
    .B(net48),
    .Y(_0106_));
 sky130_fd_sc_hd__xnor2_1 _1331_ (.A(\manchester_baby_instance.BASE_0.s_countReg[14] ),
    .B(_0662_),
    .Y(_0107_));
 sky130_fd_sc_hd__o21ai_1 _1332_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[14] ),
    .A2(_0662_),
    .B1(net34),
    .Y(_0664_));
 sky130_fd_sc_hd__nand2_1 _1333_ (.A(_0622_),
    .B(net35),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_1 _1334_ (.A(\manchester_baby_instance.BASE_0.s_countReg[16] ),
    .B(_0622_),
    .Y(_0665_));
 sky130_fd_sc_hd__and2_1 _1335_ (.A(net74),
    .B(_0622_),
    .X(_0666_));
 sky130_fd_sc_hd__o21a_1 _1336_ (.A1(_0665_),
    .A2(_0666_),
    .B1(_0630_),
    .X(_0109_));
 sky130_fd_sc_hd__xor2_1 _1337_ (.A(net36),
    .B(_0665_),
    .X(_0110_));
 sky130_fd_sc_hd__or3_1 _1338_ (.A(net62),
    .B(_0622_),
    .C(_0623_),
    .X(_0667_));
 sky130_fd_sc_hd__o21ai_1 _1339_ (.A1(_0622_),
    .A2(_0623_),
    .B1(net62),
    .Y(_0668_));
 sky130_fd_sc_hd__a21oi_1 _1340_ (.A1(_0667_),
    .A2(_0668_),
    .B1(\manchester_baby_instance.BASE_0.s_tickNext ),
    .Y(_0111_));
 sky130_fd_sc_hd__o31ai_1 _1341_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[18] ),
    .A2(_0622_),
    .A3(_0623_),
    .B1(net38),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _1342_ (.A(_0624_),
    .B(net39),
    .Y(_0112_));
 sky130_fd_sc_hd__xnor2_1 _1343_ (.A(\manchester_baby_instance.BASE_0.s_countReg[20] ),
    .B(_0624_),
    .Y(_0113_));
 sky130_fd_sc_hd__o21ai_1 _1344_ (.A1(\manchester_baby_instance.BASE_0.s_countReg[20] ),
    .A2(_0624_),
    .B1(net21),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0625_),
    .B(net22),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2_1 _1346_ (.A(\manchester_baby_instance.BASE_0.s_countReg[22] ),
    .B(_0625_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _1347_ (.A(_0626_),
    .B(_0671_),
    .Y(_0115_));
 sky130_fd_sc_hd__and2_1 _1348_ (.A(\manchester_baby_instance.BASE_0.s_countReg[23] ),
    .B(_0626_),
    .X(_0672_));
 sky130_fd_sc_hd__or2_1 _1349_ (.A(_0627_),
    .B(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_1 _1350_ (.A(_0673_),
    .X(_0116_));
 sky130_fd_sc_hd__or4b_4 _1351_ (.A(net77),
    .B(_0626_),
    .C(net59),
    .D_N(\manchester_baby_instance.BASE_0.s_countReg[25] ),
    .X(_0674_));
 sky130_fd_sc_hd__o21ai_1 _1352_ (.A1(_0616_),
    .A2(_0627_),
    .B1(_0674_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _1353_ (.A(net40),
    .B(_0628_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_1 _1354_ (.A(_0630_),
    .B(_0675_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1355_ (.A(_0639_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(_0639_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1357_ (.A(_0639_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(_0639_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1359_ (.A(_0639_),
    .Y(_0046_));
 sky130_fd_sc_hd__dfrtp_1 _1360_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0047_),
    .RESET_B(_0001_),
    .Q(\manchester_baby_instance.ram_data_o_0 ));
 sky130_fd_sc_hd__dfrtp_1 _1361_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0048_),
    .RESET_B(_0002_),
    .Q(\manchester_baby_instance.ram_data_o_1 ));
 sky130_fd_sc_hd__dfrtp_2 _1362_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0049_),
    .RESET_B(_0003_),
    .Q(\manchester_baby_instance.ram_data_o_2 ));
 sky130_fd_sc_hd__dfrtp_1 _1363_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0050_),
    .RESET_B(_0004_),
    .Q(\manchester_baby_instance.ram_data_o_3 ));
 sky130_fd_sc_hd__dfrtp_2 _1364_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0051_),
    .RESET_B(_0005_),
    .Q(\manchester_baby_instance.ram_data_o_4 ));
 sky130_fd_sc_hd__dfrtp_1 _1365_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0052_),
    .RESET_B(_0006_),
    .Q(\manchester_baby_instance.ram_data_o_5 ));
 sky130_fd_sc_hd__dfrtp_1 _1366_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0053_),
    .RESET_B(_0007_),
    .Q(\manchester_baby_instance.ram_data_o_6 ));
 sky130_fd_sc_hd__dfrtp_2 _1367_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0054_),
    .RESET_B(_0008_),
    .Q(\manchester_baby_instance.ram_data_o_7 ));
 sky130_fd_sc_hd__dfrtp_1 _1368_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0055_),
    .RESET_B(_0009_),
    .Q(\manchester_baby_instance.ram_data_o_8 ));
 sky130_fd_sc_hd__dfrtp_1 _1369_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0056_),
    .RESET_B(_0010_),
    .Q(\manchester_baby_instance.ram_data_o_9 ));
 sky130_fd_sc_hd__dfrtp_1 _1370_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0057_),
    .RESET_B(_0011_),
    .Q(\manchester_baby_instance.ram_data_o_10 ));
 sky130_fd_sc_hd__dfrtp_1 _1371_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0058_),
    .RESET_B(_0012_),
    .Q(\manchester_baby_instance.ram_data_o_11 ));
 sky130_fd_sc_hd__dfrtp_1 _1372_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0059_),
    .RESET_B(_0013_),
    .Q(\manchester_baby_instance.ram_data_o_12 ));
 sky130_fd_sc_hd__dfrtp_1 _1373_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0060_),
    .RESET_B(_0014_),
    .Q(\manchester_baby_instance.ram_data_o_13 ));
 sky130_fd_sc_hd__dfrtp_1 _1374_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0061_),
    .RESET_B(_0015_),
    .Q(\manchester_baby_instance.ram_data_o_14 ));
 sky130_fd_sc_hd__dfrtp_1 _1375_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0062_),
    .RESET_B(_0016_),
    .Q(\manchester_baby_instance.ram_data_o_15 ));
 sky130_fd_sc_hd__dfrtp_1 _1376_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0063_),
    .RESET_B(_0017_),
    .Q(\manchester_baby_instance.ram_data_o_16 ));
 sky130_fd_sc_hd__dfrtp_1 _1377_ (.CLK(clknet_3_4__leaf_clock),
    .D(_0064_),
    .RESET_B(_0018_),
    .Q(\manchester_baby_instance.ram_data_o_17 ));
 sky130_fd_sc_hd__dfrtp_1 _1378_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0065_),
    .RESET_B(_0019_),
    .Q(\manchester_baby_instance.ram_data_o_18 ));
 sky130_fd_sc_hd__dfrtp_1 _1379_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0066_),
    .RESET_B(_0020_),
    .Q(\manchester_baby_instance.ram_data_o_19 ));
 sky130_fd_sc_hd__dfrtp_1 _1380_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0067_),
    .RESET_B(_0021_),
    .Q(\manchester_baby_instance.ram_data_o_20 ));
 sky130_fd_sc_hd__dfrtp_1 _1381_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0068_),
    .RESET_B(_0022_),
    .Q(\manchester_baby_instance.ram_data_o_21 ));
 sky130_fd_sc_hd__dfrtp_1 _1382_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0069_),
    .RESET_B(_0023_),
    .Q(\manchester_baby_instance.ram_data_o_22 ));
 sky130_fd_sc_hd__dfrtp_1 _1383_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0070_),
    .RESET_B(_0024_),
    .Q(\manchester_baby_instance.ram_data_o_23 ));
 sky130_fd_sc_hd__dfrtp_1 _1384_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0071_),
    .RESET_B(_0025_),
    .Q(\manchester_baby_instance.ram_data_o_24 ));
 sky130_fd_sc_hd__dfrtp_1 _1385_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0072_),
    .RESET_B(_0026_),
    .Q(\manchester_baby_instance.ram_data_o_25 ));
 sky130_fd_sc_hd__dfrtp_1 _1386_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0073_),
    .RESET_B(_0027_),
    .Q(\manchester_baby_instance.ram_data_o_26 ));
 sky130_fd_sc_hd__dfrtp_1 _1387_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0074_),
    .RESET_B(_0028_),
    .Q(\manchester_baby_instance.ram_data_o_27 ));
 sky130_fd_sc_hd__dfrtp_1 _1388_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0075_),
    .RESET_B(_0029_),
    .Q(\manchester_baby_instance.ram_data_o_28 ));
 sky130_fd_sc_hd__dfrtp_1 _1389_ (.CLK(clknet_3_5__leaf_clock),
    .D(_0076_),
    .RESET_B(_0030_),
    .Q(\manchester_baby_instance.ram_data_o_29 ));
 sky130_fd_sc_hd__dfrtp_1 _1390_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0077_),
    .RESET_B(_0031_),
    .Q(\manchester_baby_instance.ram_data_o_30 ));
 sky130_fd_sc_hd__dfrtp_4 _1391_ (.CLK(clknet_3_7__leaf_clock),
    .D(_0078_),
    .RESET_B(_0032_),
    .Q(\manchester_baby_instance.ram_data_o_31 ));
 sky130_fd_sc_hd__dfrtp_1 _1392_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0079_),
    .RESET_B(_0033_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1393_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0080_),
    .RESET_B(_0034_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1394_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0081_),
    .RESET_B(_0035_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1395_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0082_),
    .RESET_B(_0036_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1396_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0083_),
    .RESET_B(_0037_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1397_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0084_),
    .RESET_B(_0038_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1398_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0085_),
    .RESET_B(_0039_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1399_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0086_),
    .RESET_B(_0040_),
    .Q(\manchester_baby_instance.CIRCUIT_0.IR.q[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1400_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0087_),
    .Q(\manchester_baby_instance.BASE_1.s_derivedClock ));
 sky130_fd_sc_hd__dfrtp_1 _1401_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0088_),
    .RESET_B(_0041_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _1402_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(_0089_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1403_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(_0090_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1404_ (.CLK(\manchester_baby_instance.CIRCUIT_0.GATES_13.result ),
    .D(_0091_),
    .Q(\manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1405_ (.CLK(clknet_3_6__leaf_clock),
    .D(net19),
    .Q(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1406_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0092_),
    .Q(\manchester_baby_instance.BASE_1.s_counterValue ));
 sky130_fd_sc_hd__dfxtp_2 _1407_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0093_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1408_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0094_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1409_ (.CLK(clknet_3_2__leaf_clock),
    .D(net46),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1410_ (.CLK(clknet_3_0__leaf_clock),
    .D(net25),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1411_ (.CLK(clknet_3_0__leaf_clock),
    .D(_0097_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _1412_ (.CLK(clknet_3_1__leaf_clock),
    .D(net54),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _1413_ (.CLK(clknet_3_1__leaf_clock),
    .D(net28),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _1414_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0100_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _1415_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0101_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _1416_ (.CLK(clknet_3_1__leaf_clock),
    .D(_0102_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _1417_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0103_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _1418_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0104_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _1419_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0105_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[12] ));
 sky130_fd_sc_hd__dfxtp_1 _1420_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0106_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[13] ));
 sky130_fd_sc_hd__dfxtp_1 _1421_ (.CLK(clknet_3_2__leaf_clock),
    .D(net58),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[14] ));
 sky130_fd_sc_hd__dfxtp_1 _1422_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0108_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[15] ));
 sky130_fd_sc_hd__dfxtp_1 _1423_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0109_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[16] ));
 sky130_fd_sc_hd__dfxtp_1 _1424_ (.CLK(clknet_3_2__leaf_clock),
    .D(net37),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[17] ));
 sky130_fd_sc_hd__dfxtp_1 _1425_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0111_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[18] ));
 sky130_fd_sc_hd__dfxtp_1 _1426_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0112_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[19] ));
 sky130_fd_sc_hd__dfxtp_1 _1427_ (.CLK(clknet_3_2__leaf_clock),
    .D(net52),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[20] ));
 sky130_fd_sc_hd__dfxtp_1 _1428_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0114_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[21] ));
 sky130_fd_sc_hd__dfxtp_1 _1429_ (.CLK(clknet_3_2__leaf_clock),
    .D(net33),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[22] ));
 sky130_fd_sc_hd__dfxtp_1 _1430_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0116_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[23] ));
 sky130_fd_sc_hd__dfxtp_1 _1431_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0117_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[24] ));
 sky130_fd_sc_hd__dfxtp_1 _1432_ (.CLK(clknet_3_2__leaf_clock),
    .D(_0118_),
    .Q(\manchester_baby_instance.BASE_0.s_countReg[25] ));
 sky130_fd_sc_hd__dfxtp_1 _1433_ (.CLK(clknet_3_3__leaf_clock),
    .D(\manchester_baby_instance.BASE_0.s_tickNext ),
    .Q(\manchester_baby_instance.BASE_0.s_tickReg ));
 sky130_fd_sc_hd__dlxtn_2 _1434_ (.D(ram_data_io[0]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_0 ));
 sky130_fd_sc_hd__dlxtn_1 _1435_ (.D(ram_data_io[1]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_1 ));
 sky130_fd_sc_hd__dlxtn_1 _1436_ (.D(ram_data_io[2]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_2 ));
 sky130_fd_sc_hd__dlxtn_2 _1437_ (.D(ram_data_io[3]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_3 ));
 sky130_fd_sc_hd__dlxtn_2 _1438_ (.D(ram_data_io[4]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_4 ));
 sky130_fd_sc_hd__dlxtn_1 _1439_ (.D(ram_data_io[5]),
    .GATE_N(net9),
    .Q(\manchester_baby_instance.ram_data_i_5 ));
 sky130_fd_sc_hd__dlxtn_1 _1440_ (.D(ram_data_io[6]),
    .GATE_N(net9),
    .Q(\manchester_baby_instance.ram_data_i_6 ));
 sky130_fd_sc_hd__dlxtn_1 _1441_ (.D(ram_data_io[7]),
    .GATE_N(net9),
    .Q(\manchester_baby_instance.ram_data_i_7 ));
 sky130_fd_sc_hd__dlxtn_1 _1442_ (.D(ram_data_io[8]),
    .GATE_N(net9),
    .Q(\manchester_baby_instance.ram_data_i_8 ));
 sky130_fd_sc_hd__dlxtn_1 _1443_ (.D(ram_data_io[9]),
    .GATE_N(net9),
    .Q(\manchester_baby_instance.ram_data_i_9 ));
 sky130_fd_sc_hd__dlxtn_1 _1444_ (.D(ram_data_io[10]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_10 ));
 sky130_fd_sc_hd__dlxtn_1 _1445_ (.D(ram_data_io[11]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_11 ));
 sky130_fd_sc_hd__dlxtn_1 _1446_ (.D(ram_data_io[12]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_12 ));
 sky130_fd_sc_hd__dlxtn_1 _1447_ (.D(ram_data_io[13]),
    .GATE_N(net11),
    .Q(\manchester_baby_instance.ram_data_i_13 ));
 sky130_fd_sc_hd__dlxtn_2 _1448_ (.D(ram_data_io[14]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_14 ));
 sky130_fd_sc_hd__dlxtn_2 _1449_ (.D(ram_data_io[15]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_15 ));
 sky130_fd_sc_hd__dlxtn_1 _1450_ (.D(ram_data_io[16]),
    .GATE_N(net10),
    .Q(\manchester_baby_instance.ram_data_i_16 ));
 sky130_fd_sc_hd__dlxtn_1 _1451_ (.D(ram_data_io[17]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_17 ));
 sky130_fd_sc_hd__dlxtn_1 _1452_ (.D(ram_data_io[18]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_18 ));
 sky130_fd_sc_hd__dlxtn_1 _1453_ (.D(ram_data_io[19]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_19 ));
 sky130_fd_sc_hd__dlxtn_1 _1454_ (.D(ram_data_io[20]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_20 ));
 sky130_fd_sc_hd__dlxtn_1 _1455_ (.D(ram_data_io[21]),
    .GATE_N(net13),
    .Q(\manchester_baby_instance.ram_data_i_21 ));
 sky130_fd_sc_hd__dlxtn_1 _1456_ (.D(ram_data_io[22]),
    .GATE_N(net15),
    .Q(\manchester_baby_instance.ram_data_i_22 ));
 sky130_fd_sc_hd__dlxtn_1 _1457_ (.D(ram_data_io[23]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_23 ));
 sky130_fd_sc_hd__dlxtn_1 _1458_ (.D(ram_data_io[24]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_24 ));
 sky130_fd_sc_hd__dlxtn_1 _1459_ (.D(ram_data_io[25]),
    .GATE_N(net15),
    .Q(\manchester_baby_instance.ram_data_i_25 ));
 sky130_fd_sc_hd__dlxtn_2 _1460_ (.D(ram_data_io[26]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_26 ));
 sky130_fd_sc_hd__dlxtn_1 _1461_ (.D(ram_data_io[27]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_27 ));
 sky130_fd_sc_hd__dlxtn_1 _1462_ (.D(ram_data_io[28]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_28 ));
 sky130_fd_sc_hd__dlxtn_1 _1463_ (.D(ram_data_io[29]),
    .GATE_N(net14),
    .Q(\manchester_baby_instance.ram_data_i_29 ));
 sky130_fd_sc_hd__dlxtn_1 _1464_ (.D(ram_data_io[30]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_30 ));
 sky130_fd_sc_hd__dlxtn_1 _1465_ (.D(ram_data_io[31]),
    .GATE_N(net12),
    .Q(\manchester_baby_instance.ram_data_i_31 ));
 sky130_fd_sc_hd__dlxtp_1 _1466_ (.D(\manchester_baby_instance.ram_data_o_0 ),
    .GATE(net12),
    .Q(ram_data_io[0]));
 sky130_fd_sc_hd__dlxtp_1 _1467_ (.D(\manchester_baby_instance.ram_data_o_1 ),
    .GATE(net11),
    .Q(ram_data_io[1]));
 sky130_fd_sc_hd__dlxtp_1 _1468_ (.D(\manchester_baby_instance.ram_data_o_2 ),
    .GATE(net11),
    .Q(ram_data_io[2]));
 sky130_fd_sc_hd__dlxtp_1 _1469_ (.D(\manchester_baby_instance.ram_data_o_3 ),
    .GATE(net11),
    .Q(ram_data_io[3]));
 sky130_fd_sc_hd__dlxtp_1 _1470_ (.D(\manchester_baby_instance.ram_data_o_4 ),
    .GATE(net11),
    .Q(ram_data_io[4]));
 sky130_fd_sc_hd__dlxtp_1 _1471_ (.D(\manchester_baby_instance.ram_data_o_5 ),
    .GATE(net9),
    .Q(ram_data_io[5]));
 sky130_fd_sc_hd__dlxtp_1 _1472_ (.D(\manchester_baby_instance.ram_data_o_6 ),
    .GATE(net9),
    .Q(ram_data_io[6]));
 sky130_fd_sc_hd__dlxtp_1 _1473_ (.D(\manchester_baby_instance.ram_data_o_7 ),
    .GATE(net9),
    .Q(ram_data_io[7]));
 sky130_fd_sc_hd__dlxtp_1 _1474_ (.D(\manchester_baby_instance.ram_data_o_8 ),
    .GATE(net9),
    .Q(ram_data_io[8]));
 sky130_fd_sc_hd__dlxtp_1 _1475_ (.D(\manchester_baby_instance.ram_data_o_9 ),
    .GATE(net9),
    .Q(ram_data_io[9]));
 sky130_fd_sc_hd__dlxtp_1 _1476_ (.D(\manchester_baby_instance.ram_data_o_10 ),
    .GATE(net10),
    .Q(ram_data_io[10]));
 sky130_fd_sc_hd__dlxtp_1 _1477_ (.D(\manchester_baby_instance.ram_data_o_11 ),
    .GATE(net10),
    .Q(ram_data_io[11]));
 sky130_fd_sc_hd__dlxtp_1 _1478_ (.D(\manchester_baby_instance.ram_data_o_12 ),
    .GATE(net10),
    .Q(ram_data_io[12]));
 sky130_fd_sc_hd__dlxtp_1 _1479_ (.D(\manchester_baby_instance.ram_data_o_13 ),
    .GATE(net12),
    .Q(ram_data_io[13]));
 sky130_fd_sc_hd__dlxtp_1 _1480_ (.D(\manchester_baby_instance.ram_data_o_14 ),
    .GATE(net12),
    .Q(ram_data_io[14]));
 sky130_fd_sc_hd__dlxtp_1 _1481_ (.D(\manchester_baby_instance.ram_data_o_15 ),
    .GATE(net10),
    .Q(ram_data_io[15]));
 sky130_fd_sc_hd__dlxtp_1 _1482_ (.D(\manchester_baby_instance.ram_data_o_16 ),
    .GATE(net10),
    .Q(ram_data_io[16]));
 sky130_fd_sc_hd__dlxtp_1 _1483_ (.D(\manchester_baby_instance.ram_data_o_17 ),
    .GATE(net13),
    .Q(ram_data_io[17]));
 sky130_fd_sc_hd__dlxtp_1 _1484_ (.D(\manchester_baby_instance.ram_data_o_18 ),
    .GATE(net13),
    .Q(ram_data_io[18]));
 sky130_fd_sc_hd__dlxtp_1 _1485_ (.D(\manchester_baby_instance.ram_data_o_19 ),
    .GATE(net13),
    .Q(ram_data_io[19]));
 sky130_fd_sc_hd__dlxtp_1 _1486_ (.D(\manchester_baby_instance.ram_data_o_20 ),
    .GATE(net15),
    .Q(ram_data_io[20]));
 sky130_fd_sc_hd__dlxtp_1 _1487_ (.D(\manchester_baby_instance.ram_data_o_21 ),
    .GATE(net13),
    .Q(ram_data_io[21]));
 sky130_fd_sc_hd__dlxtp_1 _1488_ (.D(\manchester_baby_instance.ram_data_o_22 ),
    .GATE(net15),
    .Q(ram_data_io[22]));
 sky130_fd_sc_hd__dlxtp_1 _1489_ (.D(\manchester_baby_instance.ram_data_o_23 ),
    .GATE(net15),
    .Q(ram_data_io[23]));
 sky130_fd_sc_hd__dlxtp_1 _1490_ (.D(\manchester_baby_instance.ram_data_o_24 ),
    .GATE(net15),
    .Q(ram_data_io[24]));
 sky130_fd_sc_hd__dlxtp_1 _1491_ (.D(\manchester_baby_instance.ram_data_o_25 ),
    .GATE(net15),
    .Q(ram_data_io[25]));
 sky130_fd_sc_hd__dlxtp_1 _1492_ (.D(\manchester_baby_instance.ram_data_o_26 ),
    .GATE(net14),
    .Q(ram_data_io[26]));
 sky130_fd_sc_hd__dlxtp_1 _1493_ (.D(\manchester_baby_instance.ram_data_o_27 ),
    .GATE(net14),
    .Q(ram_data_io[27]));
 sky130_fd_sc_hd__dlxtp_1 _1494_ (.D(\manchester_baby_instance.ram_data_o_28 ),
    .GATE(net14),
    .Q(ram_data_io[28]));
 sky130_fd_sc_hd__dlxtp_1 _1495_ (.D(\manchester_baby_instance.ram_data_o_29 ),
    .GATE(net14),
    .Q(ram_data_io[29]));
 sky130_fd_sc_hd__dlxtp_1 _1496_ (.D(\manchester_baby_instance.ram_data_o_30 ),
    .GATE(net12),
    .Q(ram_data_io[30]));
 sky130_fd_sc_hd__dlxtp_1 _1497_ (.D(\manchester_baby_instance.ram_data_o_31 ),
    .GATE(net12),
    .Q(ram_data_io[31]));
 sky130_fd_sc_hd__dfxtp_1 _1498_ (.CLK(clknet_3_6__leaf_clock),
    .D(net18),
    .Q(\manchester_baby_instance.CIRCUIT_0.GATES_13.input1 ));
 sky130_fd_sc_hd__dfxtp_1 _1499_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0000_),
    .Q(\manchester_baby_instance.CIRCUIT_0.Acc.tick ));
 sky130_fd_sc_hd__dfrtp_4 _1500_ (.CLK(clknet_3_6__leaf_clock),
    .D(_0119_),
    .RESET_B(_0042_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1501_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0120_),
    .RESET_B(_0043_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1502_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0121_),
    .RESET_B(_0044_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1503_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0122_),
    .RESET_B(_0045_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[3] ));
 sky130_fd_sc_hd__dfrtp_2 _1504_ (.CLK(clknet_3_3__leaf_clock),
    .D(_0123_),
    .RESET_B(_0046_),
    .Q(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clock (.A(clock),
    .X(clknet_0_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clock (.A(clknet_0_clock),
    .X(clknet_3_0__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clock (.A(clknet_0_clock),
    .X(clknet_3_1__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clock (.A(clknet_0_clock),
    .X(clknet_3_2__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clock (.A(clknet_0_clock),
    .X(clknet_3_3__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clock (.A(clknet_0_clock),
    .X(clknet_3_4__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clock (.A(clknet_0_clock),
    .X(clknet_3_5__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clock (.A(clknet_0_clock),
    .X(clknet_3_6__leaf_clock));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clock (.A(clknet_0_clock),
    .X(clknet_3_7__leaf_clock));
 sky130_fd_sc_hd__clkbuf_2 fanout10 (.A(net16),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 fanout11 (.A(net16),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 fanout12 (.A(net16),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net15),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 fanout16 (.A(net7),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout9 (.A(net16),
    .X(net9));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0653_),
    .X(net27));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0099_),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\manchester_baby_instance.BASE_0.s_countReg[12] ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0661_),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0115_),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\manchester_baby_instance.BASE_0.s_countReg[15] ),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0664_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\manchester_baby_instance.BASE_1.s_bufferRegs[0] ),
    .X(net18));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\manchester_baby_instance.BASE_0.s_countReg[17] ),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0110_),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\manchester_baby_instance.BASE_0.s_countReg[19] ),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0669_),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\manchester_baby_instance.BASE_0.s_countReg[25] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\manchester_baby_instance.BASE_0.s_countReg[4] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_0652_),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\manchester_baby_instance.BASE_0.s_countReg[2] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_0649_),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\manchester_baby_instance.BASE_1.s_derivedClock ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0095_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0663_),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\manchester_baby_instance.BASE_0.s_countReg[9] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0657_),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0113_),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0098_),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\manchester_baby_instance.BASE_1.s_counterValue ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .X(net20));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0644_),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0107_),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\manchester_baby_instance.BASE_0.s_countReg[24] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net8),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\manchester_baby_instance.BASE_0.s_countReg[1] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\manchester_baby_instance.BASE_0.s_countReg[18] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\manchester_baby_instance.BASE_0.s_tickReg ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0660_),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\manchester_baby_instance.BASE_0.s_countReg[21] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0656_),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB[4] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\manchester_baby_instance.ram_data_o_0 ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[0] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[1] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[4] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[2] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\manchester_baby_instance.BASE_0.s_countReg[16] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\manchester_baby_instance.CIRCUIT_0.IR.q[3] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0670_),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\manchester_baby_instance.BASE_0.s_countReg[23] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\manchester_baby_instance.BASE_0.s_countReg[23] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0650_),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0096_),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input1 (.A(reset_i),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 output2 (.A(net2),
    .X(ram_addr_o[0]));
 sky130_fd_sc_hd__clkbuf_4 output3 (.A(net3),
    .X(ram_addr_o[1]));
 sky130_fd_sc_hd__clkbuf_4 output4 (.A(net4),
    .X(ram_addr_o[2]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(ram_addr_o[3]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(ram_addr_o[4]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net15),
    .X(ram_rw_en_o));
 sky130_fd_sc_hd__clkbuf_4 output8 (.A(net8),
    .X(stop_lamp_o));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\manchester_baby_instance.BASE_0.s_countReg[0] ),
    .X(net17));
endmodule

