VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO openlane_manchester_baby
  CLASS BLOCK ;
  FOREIGN openlane_manchester_baby ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 187.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 194.360 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 194.360 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 194.360 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 194.360 181.510 ;
    END
  END VPWR
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END clock
  PIN ram_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 200.000 ;
    END
  END ram_addr_o[0]
  PIN ram_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 200.000 ;
    END
  END ram_addr_o[1]
  PIN ram_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 77.370 196.000 77.650 200.000 ;
    END
  END ram_addr_o[2]
  PIN ram_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END ram_addr_o[3]
  PIN ram_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END ram_addr_o[4]
  PIN ram_data_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END ram_data_io[0]
  PIN ram_data_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END ram_data_io[10]
  PIN ram_data_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END ram_data_io[11]
  PIN ram_data_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END ram_data_io[12]
  PIN ram_data_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END ram_data_io[13]
  PIN ram_data_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 81.640 200.000 82.240 ;
    END
  END ram_data_io[14]
  PIN ram_data_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 71.440 200.000 72.040 ;
    END
  END ram_data_io[15]
  PIN ram_data_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END ram_data_io[16]
  PIN ram_data_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END ram_data_io[17]
  PIN ram_data_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END ram_data_io[18]
  PIN ram_data_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 51.040 200.000 51.640 ;
    END
  END ram_data_io[19]
  PIN ram_data_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END ram_data_io[1]
  PIN ram_data_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END ram_data_io[20]
  PIN ram_data_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 74.840 200.000 75.440 ;
    END
  END ram_data_io[21]
  PIN ram_data_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 200.000 78.840 ;
    END
  END ram_data_io[22]
  PIN ram_data_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 91.840 200.000 92.440 ;
    END
  END ram_data_io[23]
  PIN ram_data_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 98.640 200.000 99.240 ;
    END
  END ram_data_io[24]
  PIN ram_data_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 122.440 200.000 123.040 ;
    END
  END ram_data_io[25]
  PIN ram_data_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 129.240 200.000 129.840 ;
    END
  END ram_data_io[26]
  PIN ram_data_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 125.840 200.000 126.440 ;
    END
  END ram_data_io[27]
  PIN ram_data_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 115.640 200.000 116.240 ;
    END
  END ram_data_io[28]
  PIN ram_data_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 88.440 200.000 89.040 ;
    END
  END ram_data_io[29]
  PIN ram_data_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END ram_data_io[2]
  PIN ram_data_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 196.000 95.240 200.000 95.840 ;
    END
  END ram_data_io[30]
  PIN ram_data_io[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 116.010 196.000 116.290 200.000 ;
    END
  END ram_data_io[31]
  PIN ram_data_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END ram_data_io[3]
  PIN ram_data_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END ram_data_io[4]
  PIN ram_data_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END ram_data_io[5]
  PIN ram_data_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END ram_data_io[6]
  PIN ram_data_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ram_data_io[7]
  PIN ram_data_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END ram_data_io[8]
  PIN ram_data_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END ram_data_io[9]
  PIN ram_rw_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 40.840 200.000 41.440 ;
    END
  END ram_rw_en_o
  PIN reset_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 85.040 200.000 85.640 ;
    END
  END reset_i
  PIN stop_lamp_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 196.000 109.850 200.000 ;
    END
  END stop_lamp_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 187.765 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.510 187.920 ;
      LAYER met2 ;
        RECT 4.690 195.720 77.090 196.000 ;
        RECT 77.930 195.720 86.750 196.000 ;
        RECT 87.590 195.720 96.410 196.000 ;
        RECT 97.250 195.720 109.290 196.000 ;
        RECT 110.130 195.720 115.730 196.000 ;
        RECT 116.570 195.720 194.490 196.000 ;
        RECT 4.690 4.280 194.490 195.720 ;
        RECT 4.690 4.000 54.550 4.280 ;
        RECT 55.390 4.000 70.650 4.280 ;
        RECT 71.490 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 106.070 4.280 ;
        RECT 106.910 4.000 115.730 4.280 ;
        RECT 116.570 4.000 125.390 4.280 ;
        RECT 126.230 4.000 144.710 4.280 ;
        RECT 145.550 4.000 194.490 4.280 ;
      LAYER met3 ;
        RECT 4.000 150.640 196.000 187.845 ;
        RECT 4.400 149.240 196.000 150.640 ;
        RECT 4.000 130.240 196.000 149.240 ;
        RECT 4.000 128.840 195.600 130.240 ;
        RECT 4.000 126.840 196.000 128.840 ;
        RECT 4.400 125.440 195.600 126.840 ;
        RECT 4.000 123.440 196.000 125.440 ;
        RECT 4.400 122.040 195.600 123.440 ;
        RECT 4.000 116.640 196.000 122.040 ;
        RECT 4.000 115.240 195.600 116.640 ;
        RECT 4.000 113.240 196.000 115.240 ;
        RECT 4.400 111.840 196.000 113.240 ;
        RECT 4.000 109.840 196.000 111.840 ;
        RECT 4.400 108.440 196.000 109.840 ;
        RECT 4.000 103.040 196.000 108.440 ;
        RECT 4.400 101.640 196.000 103.040 ;
        RECT 4.000 99.640 196.000 101.640 ;
        RECT 4.400 98.240 195.600 99.640 ;
        RECT 4.000 96.240 196.000 98.240 ;
        RECT 4.000 94.840 195.600 96.240 ;
        RECT 4.000 92.840 196.000 94.840 ;
        RECT 4.400 91.440 195.600 92.840 ;
        RECT 4.000 89.440 196.000 91.440 ;
        RECT 4.000 88.040 195.600 89.440 ;
        RECT 4.000 86.040 196.000 88.040 ;
        RECT 4.000 84.640 195.600 86.040 ;
        RECT 4.000 82.640 196.000 84.640 ;
        RECT 4.000 81.240 195.600 82.640 ;
        RECT 4.000 79.240 196.000 81.240 ;
        RECT 4.400 77.840 195.600 79.240 ;
        RECT 4.000 75.840 196.000 77.840 ;
        RECT 4.000 74.440 195.600 75.840 ;
        RECT 4.000 72.440 196.000 74.440 ;
        RECT 4.000 71.040 195.600 72.440 ;
        RECT 4.000 69.040 196.000 71.040 ;
        RECT 4.400 67.640 196.000 69.040 ;
        RECT 4.000 62.240 196.000 67.640 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 58.840 196.000 60.840 ;
        RECT 4.400 57.440 196.000 58.840 ;
        RECT 4.000 52.040 196.000 57.440 ;
        RECT 4.000 50.640 195.600 52.040 ;
        RECT 4.000 41.840 196.000 50.640 ;
        RECT 4.000 40.440 195.600 41.840 ;
        RECT 4.000 10.715 196.000 40.440 ;
      LAYER met4 ;
        RECT 93.215 82.455 125.745 116.105 ;
  END
END openlane_manchester_baby
END LIBRARY

