* NGSPICE file created from manchester_baby.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

.subckt manchester_baby VGND VPWR clock clock_o ram_addr_o[0] ram_addr_o[1] ram_addr_o[2]
+ ram_addr_o[3] ram_addr_o[4] ram_data_i[0] ram_data_i[10] ram_data_i[11] ram_data_i[12]
+ ram_data_i[13] ram_data_i[14] ram_data_i[15] ram_data_i[16] ram_data_i[17] ram_data_i[18]
+ ram_data_i[19] ram_data_i[1] ram_data_i[20] ram_data_i[21] ram_data_i[22] ram_data_i[23]
+ ram_data_i[24] ram_data_i[25] ram_data_i[26] ram_data_i[27] ram_data_i[28] ram_data_i[29]
+ ram_data_i[2] ram_data_i[30] ram_data_i[31] ram_data_i[3] ram_data_i[4] ram_data_i[5]
+ ram_data_i[6] ram_data_i[7] ram_data_i[8] ram_data_i[9] ram_data_o[0] ram_data_o[10]
+ ram_data_o[11] ram_data_o[12] ram_data_o[13] ram_data_o[14] ram_data_o[15] ram_data_o[16]
+ ram_data_o[17] ram_data_o[18] ram_data_o[19] ram_data_o[1] ram_data_o[20] ram_data_o[21]
+ ram_data_o[22] ram_data_o[23] ram_data_o[24] ram_data_o[25] ram_data_o[26] ram_data_o[27]
+ ram_data_o[28] ram_data_o[29] ram_data_o[2] ram_data_o[30] ram_data_o[31] ram_data_o[3]
+ ram_data_o[4] ram_data_o[5] ram_data_o[6] ram_data_o[7] ram_data_o[8] ram_data_o[9]
+ ram_rw_en_o reset_i stop_lamp_o
XFILLER_0_43_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0985_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0494_ _0500_ _0492_
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_269 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0770_ net87 _0267_ _0309_ _0312_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__o22a_1
X_0968_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0899_ _0158_ _0157_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_2_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0822_ net8 _0127_ _0128_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or3_1
X_0753_ net19 _0133_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0684_ _0201_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__and2b_1
X_1098_ clknet_2_3__leaf_clock _0051_ _0002_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1021_ net73 net34 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_36_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0805_ _0271_ _0322_ _0342_ _0276_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0667_ net48 net9 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and2b_1
X_0598_ net67 net28 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and2b_1
X_0736_ net22 _0281_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 manchester_baby_instance.CIRCUIT_0.IR.q\[2\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_275 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0494_ _0517_ _0492_
+ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0719_ _0265_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput64 net64 VGND VGND VPWR VPWR ram_data_o[31] sky130_fd_sc_hd__clkbuf_4
Xoutput42 net42 VGND VGND VPWR VPWR ram_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput53 net53 VGND VGND VPWR VPWR ram_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0984_ _0464_ _0496_ _0497_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a211o_1
XFILLER_0_13_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0967_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0479_ _0483_ VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ _0155_ _0160_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0752_ _0271_ _0295_ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__and3_1
X_0821_ _0356_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ _0199_ _0202_ _0212_ _0229_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_24_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1097_ clknet_2_3__leaf_clock _0050_ _0001_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1020_ _0528_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0804_ _0218_ _0224_ _0320_ _0229_ _0207_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o311ai_1
X_0735_ net21 net22 _0134_ _0274_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o31ai_2
X_0597_ _0141_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__nand2_1
X_0666_ _0213_ _0214_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nand2_1
X_1149_ clknet_2_1__leaf_clock _0098_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold31 net63 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 net69 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1003_ _0487_ _0502_ _0511_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ _0118_ _0264_ _0266_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0649_ net54 net15 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_11_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput43 net43 VGND VGND VPWR VPWR ram_data_o[12] sky130_fd_sc_hd__buf_2
Xoutput54 net54 VGND VGND VPWR VPWR ram_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput65 net65 VGND VGND VPWR VPWR ram_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ net26 _0477_ _0498_ _0482_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0966_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR VPWR
+ _0483_ sky130_fd_sc_hd__or3_1
X_0897_ _0421_ _0162_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0751_ _0234_ _0235_ _0294_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0820_ net49 _0355_ _0265_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
X_0682_ _0204_ _0210_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or3_1
X_1096_ clknet_2_1__leaf_clock _0000_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.Acc.tick
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_29_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0949_ net23 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] VGND VGND VPWR
+ VPWR _0466_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_30_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0803_ _0268_ _0337_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and3_1
X_0665_ net47 net8 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__or2b_1
X_0734_ net21 _0134_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or2_1
X_0596_ _0142_ _0143_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1148_ clknet_2_1__leaf_clock _0097_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_counterValue
+ sky130_fd_sc_hd__dfxtp_1
X_1079_ _0533_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold10 manchester_baby_instance.BASE_1.s_counterValue VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 manchester_baby_instance.CIRCUIT_0.IR.q\[4\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net60 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ net12 _0477_ _0513_ _0481_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ net64 _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0648_ _0182_ _0189_ _0192_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__o211a_1
X_0579_ net7 net6 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput55 net55 VGND VGND VPWR VPWR ram_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR ram_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput66 net66 VGND VGND VPWR VPWR ram_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0982_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0480_ VGND VGND VPWR
+ VPWR _0498_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0965_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0480_ _0481_ VGND
+ VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a21boi_1
X_0896_ net68 _0156_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ _0235_ _0294_ _0234_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0681_ _0208_ net14 _0205_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o21a_1
X_1095_ clknet_2_1__leaf_clock net76 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfxtp_1
X_0948_ net26 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] VGND VGND VPWR
+ VPWR _0465_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_22_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0879_ _0121_ _0122_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0802_ net13 _0336_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0733_ _0138_ _0253_ _0254_ _0256_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0664_ net8 net47 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0595_ net12 net51 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1147_ clknet_2_1__leaf_clock net77 VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_bufferRegs\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1078_ _0533_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 _0538_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 net70 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 manchester_baby_instance.CIRCUIT_0.IR.q\[1\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ _0469_ _0464_ _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0578_ net5 net4 _0125_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__or4_4
X_0647_ net7 _0193_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a21o_1
X_0716_ _0117_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__buf_4
Xoutput34 net34 VGND VGND VPWR VPWR clock_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput56 net56 VGND VGND VPWR VPWR ram_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput67 net67 VGND VGND VPWR VPWR ram_data_o[5] sky130_fd_sc_hd__buf_2
Xoutput45 net45 VGND VGND VPWR VPWR ram_data_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_34_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0981_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0479_ _0484_ VGND
+ VGND VPWR VPWR _0497_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_14_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clock clock VGND VGND VPWR VPWR clknet_0_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0964_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0462_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__and4b_1
XFILLER_0_40_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0895_ _0406_ _0123_ _0419_ _0288_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0680_ _0224_ _0227_ _0228_ _0220_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__o22a_1
X_1094_ _0541_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0947_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0462_ _0463_ VGND VGND VPWR
+ VPWR _0464_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_30_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0878_ net41 _0118_ _0403_ _0405_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_132 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0801_ net92 _0267_ _0335_ _0339_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0732_ _0256_ _0254_ _0253_ _0138_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__o211ai_1
X_0594_ net40 _0112_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__or2b_1
X_0663_ _0204_ _0207_ _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ clknet_2_1__leaf_clock net86 _0049_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1077_ _0533_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold12 net73 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 manchester_baby_instance.CIRCUIT_0.IR.q\[3\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 net65 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _0112_ _0501_ _0467_ _0468_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0715_ _0120_ _0136_ _0261_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0577_ net2 net3 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__or2_1
X_0646_ net7 _0193_ _0194_ net6 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__o22a_1
X_1129_ clknet_2_1__leaf_clock _0082_ _0033_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dfrtp_2
Xoutput35 net35 VGND VGND VPWR VPWR ram_addr_o[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput46 net46 VGND VGND VPWR VPWR ram_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput57 net57 VGND VGND VPWR VPWR ram_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VGND VGND VPWR VPWR ram_data_o[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0629_ _0176_ _0177_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0495_ _0472_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0963_ net64 _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__and2_1
X_0894_ net30 _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ net79 _0524_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0946_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0877_ _0288_ _0398_ _0404_ _0275_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0800_ _0288_ _0131_ _0338_ _0276_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0731_ _0115_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_4
X_0593_ net12 net51 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__xnor2_1
X_0662_ _0209_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[2\]
+ _0048_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_35_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1076_ _0537_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0929_ _0268_ net74 _0449_ _0275_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_45_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold13 _0096_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 net43 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 net51 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0714_ _0137_ _0259_ _0260_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0645_ net45 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__inv_2
X_0576_ _0121_ _0122_ _0123_ _0124_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__or4_4
X_1128_ clknet_2_1__leaf_clock _0081_ _0032_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dfrtp_1
X_1059_ _0536_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput36 net36 VGND VGND VPWR VPWR ram_addr_o[1] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR ram_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_9_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput69 net69 VGND VGND VPWR VPWR ram_data_o[7] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR ram_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ net43 net4 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__or2b_1
X_0559_ _0110_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0962_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\]
+ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] VGND VGND VPWR VPWR _0479_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0893_ net29 _0406_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1092_ _0524_ _0540_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0945_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0462_ sky130_fd_sc_hd__and3b_1
XFILLER_0_2_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0876_ net2 _0125_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0730_ net104 _0267_ _0270_ _0277_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0661_ _0208_ net14 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0592_ net23 net62 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1144_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
+ _0047_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_35_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1075_ _0537_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ _0389_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_0928_ net26 _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__nand2_1
Xhold25 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] VGND VGND VPWR VPWR
+ net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 net57 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0713_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] _0119_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0644_ net46 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__inv_2
X_0575_ net31 net32 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__or2_1
X_1058_ _0536_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
X_1127_ clknet_2_0__leaf_clock _0080_ _0031_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput59 net59 VGND VGND VPWR VPWR ram_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR ram_addr_o[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput48 net48 VGND VGND VPWR VPWR ram_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_19_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0558_ net103 net23 _0104_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0627_ net4 net43 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0961_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] VGND VGND VPWR VPWR
+ _0478_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0892_ net95 _0118_ _0415_ _0417_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1091_ net78 net81 VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
X_0944_ _0112_ _0267_ _0459_ _0461_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0875_ _0307_ _0395_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0660_ _0208_ net14 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0591_ net23 net62 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1143_ manchester_baby_instance.CIRCUIT_0.GATES_13.result manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
+ _0046_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1074_ _0537_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0927_ net23 _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0789_ net15 _0131_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nand2_1
X_0858_ net44 _0388_ _0117_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
Xhold15 net71 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net47 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0712_ _0137_ _0259_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0574_ net29 net30 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__or2_1
X_0643_ _0174_ _0175_ _0180_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__or4_1
XFILLER_0_32_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1126_ clknet_2_0__leaf_clock _0079_ _0030_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dfrtp_1
X_1057_ _0536_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
Xoutput38 net38 VGND VGND VPWR VPWR ram_addr_o[3] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR ram_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_11_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0557_ _0109_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0626_ net7 net46 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__xor2_1
X_1109_ clknet_2_2__leaf_clock _0062_ _0013_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0609_ net30 net69 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0960_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0462_ _0463_ VGND VGND VPWR
+ VPWR _0477_ sky130_fd_sc_hd__and3b_1
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0891_ _0271_ _0410_ _0416_ _0275_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ net78 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
X_0874_ _0165_ _0186_ _0394_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and3_1
X_0943_ _0276_ _0460_ net40 VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0590_ net75 net65 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__or2b_1
X_1142_ clknet_2_1__leaf_clock _0095_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_1.s_derivedClock
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1073_ _0537_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0857_ _0274_ _0127_ _0385_ _0387_ _0278_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a32o_1
X_0926_ net12 _0112_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or2_1
Xhold27 manchester_baby_instance.CIRCUIT_0.IR.q\[0\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0788_ _0200_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__nand2_1
Xhold16 net56 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_2__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_2__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0711_ net64 net25 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0573_ net27 net28 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__or2_1
X_0642_ net5 _0190_ _0176_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__o21a_1
X_1125_ clknet_2_0__leaf_clock _0078_ _0029_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1056_ _0536_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
Xoutput39 net39 VGND VGND VPWR VPWR ram_addr_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0909_ net27 _0121_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0625_ net6 net45 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0556_ net107 net26 _0104_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1039_ _0534_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
X_1108_ clknet_2_2__leaf_clock _0061_ _0012_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0608_ net69 net30 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0890_ _0367_ _0172_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0942_ _0112_ _0307_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nor2_1
X_0873_ _0185_ _0276_ _0401_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1141_ clknet_2_3__leaf_clock _0094_ _0045_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_1072_ _0537_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0787_ _0230_ _0322_ _0210_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0856_ _0181_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__xnor2_1
X_0925_ _0271_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 net52 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 net68 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0710_ _0138_ _0253_ _0255_ _0256_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0641_ net44 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0572_ net26 net23 net12 net1 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__or4_4
X_1124_ clknet_2_0__leaf_clock _0077_ _0028_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dfrtp_1
X_1055_ net33 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0908_ net101 _0118_ _0429_ _0431_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__o22a_1
X_0839_ _0175_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0624_ _0166_ _0169_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0555_ _0108_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1038_ _0534_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1107_ clknet_2_2__leaf_clock _0060_ _0011_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0607_ net29 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0941_ net40 _0307_ _0120_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__o21ai_1
X_0872_ _0307_ _0397_ _0400_ _0265_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ _0537_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
X_1140_ clknet_2_3__leaf_clock _0093_ _0044_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0924_ _0443_ _0154_ _0140_ _0146_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0786_ net91 _0267_ _0319_ _0326_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__o22a_1
X_0855_ _0176_ _0369_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
Xhold29 net59 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 net55 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0571_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ _0119_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] VGND VGND VPWR VPWR _0120_
+ sky130_fd_sc_hd__or4b_1
X_0640_ _0185_ net3 _0166_ _0186_ _0188_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1123_ clknet_2_0__leaf_clock _0076_ _0027_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dfrtp_1
X_1054_ _0535_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0907_ _0288_ _0418_ _0430_ _0275_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0838_ net6 _0194_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o21ai_1
X_0769_ _0288_ _0133_ _0311_ _0276_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0554_ net105 net27 _0104_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0623_ _0170_ _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nand2_1
X_1106_ clknet_2_2__leaf_clock _0059_ _0010_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfrtp_1
X_1037_ _0534_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0606_ _0139_ _0140_ _0146_ _0153_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__a311o_1
XFILLER_0_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0940_ net108 _0118_ _0456_ _0458_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0871_ net3 _0398_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_38_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1070_ _0537_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0854_ net5 _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
X_0923_ _0140_ _0146_ _0443_ _0154_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0785_ _0324_ _0325_ _0118_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o21ai_1
Xhold19 net53 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0570_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0119_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ clknet_2_0__leaf_clock _0075_ _0026_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1053_ _0535_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0906_ net29 _0406_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0837_ _0191_ _0369_ _0174_ _0180_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a211o_1
X_0699_ net20 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__inv_2
X_0768_ net18 _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0553_ _0107_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_0622_ net70 net31 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__or2b_1
X_1105_ clknet_2_3__leaf_clock _0058_ _0009_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfrtp_1
X_1036_ _0534_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0605_ net65 net75 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__and2b_1
X_1019_ _0525_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_220 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ net3 _0398_ _0274_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0999_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0512_ VGND VGND VPWR
+ VPWR _0513_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ net4 _0125_ _0126_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or3_1
X_0922_ net75 net65 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0784_ _0199_ _0203_ _0323_ _0307_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 ram_data_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ clknet_2_0__leaf_clock _0074_ _0025_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dfrtp_1
X_1052_ _0535_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0836_ _0189_ _0368_ _0178_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a21o_1
X_0905_ _0271_ _0423_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__and3_1
X_0767_ net17 _0132_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0698_ _0238_ _0240_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0621_ net31 net70 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0552_ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] net5 _0104_ VGND VGND VPWR VPWR
+ _0107_ sky130_fd_sc_hd__mux2_1
X_1035_ _0534_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
X_1104_ clknet_2_3__leaf_clock _0057_ _0008_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0819_ _0274_ _0344_ _0352_ _0354_ _0278_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0604_ _0149_ _0152_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1018_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0527_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_14_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_135 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ net64 _0501_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0442_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0783_ _0199_ _0323_ _0203_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__a21oi_1
X_0852_ _0383_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 ram_data_i[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1120_ clknet_2_0__leaf_clock _0073_ _0024_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dfrtp_1
X_1051_ _0535_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0904_ _0155_ _0160_ _0422_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__nand3_1
X_0835_ _0367_ _0173_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__or2_1
X_0766_ _0306_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nor2_1
X_0697_ _0239_ _0242_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_44_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0551_ _0106_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_0620_ _0167_ _0168_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1034_ _0534_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1103_ clknet_2_2__leaf_clock _0056_ _0007_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _0347_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nor2_1
X_0749_ _0246_ _0292_ _0293_ _0240_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_38_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0603_ _0150_ _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1017_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\]
+ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0997_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0501_ VGND VGND VPWR
+ VPWR _0511_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ net66 _0441_ _0117_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
X_0782_ _0230_ _0322_ _0200_ _0210_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a211o_1
X_0851_ net45 _0382_ _0117_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 ram_data_i[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ _0535_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0903_ net93 _0118_ _0420_ _0427_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__o22a_1
X_0834_ _0155_ _0161_ _0163_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0696_ _0226_ _0233_ _0238_ _0241_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a2111o_1
X_0765_ _0241_ _0242_ _0292_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a31o_1
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0550_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] net6 _0104_ VGND VGND VPWR VPWR
+ _0106_ sky130_fd_sc_hd__mux2_1
X_1102_ clknet_2_3__leaf_clock _0055_ _0006_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1033_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__buf_4
X_0817_ _0218_ _0320_ _0227_ _0223_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0748_ _0237_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__inv_2
X_0679_ _0219_ _0221_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0602_ net66 net27 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1016_ _0526_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0996_ _0492_ _0509_ _0510_ net98 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ _0278_ _0370_ _0379_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0781_ _0228_ _0321_ _0207_ _0220_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a211o_1
Xinput4 ram_data_i[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_0979_ _0473_ _0465_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0902_ _0425_ _0426_ _0265_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__o21ai_1
X_0833_ net99 _0267_ _0364_ _0366_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__o22a_1
X_0764_ _0262_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0695_ _0242_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1101_ clknet_2_3__leaf_clock _0054_ _0005_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1032_ net33 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_16_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ net10 _0129_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0747_ _0291_ _0244_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0678_ _0213_ _0217_ _0216_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0601_ net27 net66 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1015_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[14\]
+ manchester_baby_instance.CIRCUIT_0.IR.q\[13\] _0525_ VGND VGND VPWR VPWR _0526_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_28_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0487_ _0502_ _0494_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0780_ _0213_ _0217_ _0320_ _0223_ _0216_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__a311o_1
XFILLER_0_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput5 ram_data_i[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_0978_ _0486_ _0492_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_40_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0901_ _0421_ _0424_ _0423_ _0307_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a31o_1
X_0832_ _0288_ _0357_ _0365_ _0276_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a31o_1
X_0763_ _0242_ _0292_ _0241_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0694_ net56 net17 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1100_ clknet_2_3__leaf_clock _0053_ _0004_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_1031_ _0532_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0815_ _0351_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
Xinput30 ram_data_i[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
X_0746_ _0226_ _0233_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0677_ _0184_ _0197_ _0212_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0600_ _0147_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR VPWR
+ _0525_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0729_ _0271_ _0259_ _0273_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0994_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0483_ _0502_ _0508_
+ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 ram_data_i[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ _0493_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0421_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21oi_1
X_0762_ _0305_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_0831_ _0127_ _0128_ net8 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o21ai_1
X_0693_ net17 net56 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1030_ net76 net77 VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2b_1
Xinput20 ram_data_i[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0814_ net50 _0350_ _0265_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
Xinput31 ram_data_i[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0676_ _0215_ _0218_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or3_1
X_0745_ net94 _0267_ _0287_ _0290_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ net79 _0524_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_tickNext
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0659_ net53 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0728_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _0464_ _0503_ _0504_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput7 ram_data_i[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
X_0976_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0491_ _0492_ VGND
+ VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0830_ _0363_ _0271_ _0320_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__and3b_1
X_0761_ net58 _0304_ _0265_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0692_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or2_1
X_0959_ _0474_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput21 ram_data_i[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput10 ram_data_i[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput32 ram_data_i[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_0813_ _0268_ _0336_ _0345_ _0349_ _0278_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a32o_1
X_0675_ _0219_ _0220_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0744_ _0288_ _0281_ _0289_ _0276_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a31o_1
X_1089_ _0539_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1012_ manchester_baby_instance.BASE_0.s_countReg\[0\] net81 VGND VGND VPWR VPWR
+ _0524_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0727_ _0115_ _0274_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0275_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0658_ _0205_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0589_ net21 net60 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0992_ _0481_ _0505_ _0506_ _0477_ net23 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a32o_1
Xclkbuf_2_1__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_1__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 ram_data_i[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_0975_ _0462_ _0487_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0760_ _0268_ _0298_ _0301_ _0303_ _0278_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0691_ net57 net18 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0958_ net27 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] VGND VGND VPWR
+ VPWR _0475_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0889_ _0268_ _0407_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput22 ram_data_i[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 ram_data_i[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
X_0812_ _0346_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_286 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 reset_i VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
X_0743_ net21 _0134_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nand2_1
X_0674_ _0221_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__or2_1
X_1088_ manchester_baby_instance.BASE_0.s_tickReg net83 VGND VGND VPWR VPWR _0539_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ _0492_ _0522_ _0523_ _0501_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0726_ _0116_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0588_ net24 net63 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_4_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0657_ net52 net13 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0709_ _0137_ _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ net64 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0501_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
+ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 ram_data_i[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_0_39_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0974_ _0464_ _0476_ _0477_ net27 _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0690_ net18 net57 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0957_ _0465_ _0472_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0888_ _0406_ _0123_ net31 VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 ram_data_i[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_4
Xinput23 ram_data_i[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_6
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ net49 net10 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__and2b_1
X_0811_ _0221_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__nor2_1
X_0742_ _0268_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1087_ _0533_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1010_ _0494_ _0519_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0725_ _0258_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nand2_1
X_0656_ net13 net52 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0587_ net25 _0135_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_4_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1139_ clknet_2_3__leaf_clock _0092_ _0043_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0708_ net63 net24 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or2b_1
X_0639_ _0185_ net3 net2 _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_13_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ _0480_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0478_ _0482_ _0484_ _0486_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o41a_1
XFILLER_0_13_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ net26 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] VGND VGND VPWR
+ VPWR _0473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_288 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ net88 _0118_ _0409_ _0413_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 ram_data_i[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_0810_ _0213_ _0217_ _0320_ _0223_ _0216_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a311oi_2
Xinput24 ram_data_i[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0672_ net10 net49 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__and2b_1
X_0741_ _0252_ _0245_ _0247_ _0250_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a41oi_1
X_1086_ _0533_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0939_ _0268_ _0447_ _0457_ _0275_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ _0138_ _0253_ _0255_ _0256_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a31o_1
X_0655_ _0200_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0586_ net21 net22 net24 _0134_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_4_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1138_ clknet_2_3__leaf_clock _0091_ _0042_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1069_ _0537_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0707_ net61 net22 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0638_ net41 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__inv_2
X_0569_ _0117_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0972_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0487_ _0479_ _0488_
+ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0955_ _0466_ _0470_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__a21bo_1
X_0886_ _0411_ _0412_ _0265_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput25 ram_data_i[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
Xinput14 ram_data_i[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_0740_ _0271_ _0253_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
X_0671_ net50 net11 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__and2b_1
X_1085_ _0533_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__inv_2
X_0869_ net2 _0125_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0938_ net12 _0112_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0723_ _0115_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0654_ _0201_ _0202_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0585_ net19 net20 _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__or3_4
X_1137_ clknet_2_3__leaf_clock _0090_ _0041_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1068_ _0537_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 manchester_baby_instance.BASE_1.s_bufferRegs\[0\] VGND VGND VPWR VPWR net76
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0706_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0637_ _0168_ _0170_ _0167_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a21o_1
X_0568_ _0115_ _0116_ manchester_baby_instance.CIRCUIT_0.Acc.tick VGND VGND VPWR VPWR
+ _0117_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0481_ _0480_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\]
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0954_ net23 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] VGND VGND VPWR
+ VPWR _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0885_ _0169_ _0170_ _0410_ _0307_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput26 ram_data_i[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_8
X_0670_ net11 net50 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__and2b_1
Xinput15 ram_data_i[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
X_1084_ _0533_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0937_ _0142_ _0143_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o21a_1
X_0868_ _0164_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__xnor2_1
X_0799_ net14 _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0653_ net55 net16 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2b_1
X_0722_ _0268_ _0135_ _0269_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and3_1
X_0584_ net17 net18 _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__or3_4
XFILLER_0_47_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1136_ clknet_2_3__leaf_clock _0089_ _0040_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1067_ _0537_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold4 manchester_baby_instance.BASE_1.s_derivedClock VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0705_ net22 net61 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__and2b_1
X_0636_ net42 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0567_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ _0101_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] VGND VGND VPWR VPWR _0116_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1119_ clknet_2_0__leaf_clock _0072_ _0023_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_160 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0619_ net32 net71 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0970_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR VPWR
+ _0487_ sky130_fd_sc_hd__nor3_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_130 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ net12 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0469_ VGND VGND
+ VPWR VPWR _0470_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0884_ _0170_ _0410_ _0169_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_222 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 ram_data_i[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
Xinput16 ram_data_i[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_1083_ net77 net84 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__xnor2_1
X_1152_ clknet_2_1__leaf_clock net80 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_tickReg
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0936_ _0142_ _0143_ _0307_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0798_ net13 _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or2_1
X_0867_ _0187_ net2 _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0652_ net16 net55 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__and2b_1
X_0583_ net15 net16 _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or3_4
X_0721_ net21 net22 _0134_ net24 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_26_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1135_ clknet_2_3__leaf_clock _0088_ _0039_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1066_ net33 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0919_ _0274_ _0432_ _0439_ _0440_ _0278_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 manchester_baby_instance.BASE_0.s_countReg\[0\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0566_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__buf_2
X_0635_ _0155_ _0161_ _0163_ _0183_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a211o_1
X_0704_ _0245_ _0247_ _0250_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_48_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1049_ _0535_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
X_1118_ clknet_2_0__leaf_clock _0071_ _0022_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0549_ _0105_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_0618_ net71 net32 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ _0112_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] _0467_ _0468_
+ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0883_ _0367_ _0172_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput17 ram_data_i[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
Xinput28 ram_data_i[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
X_1151_ clknet_2_1__leaf_clock _0100_ VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1082_ net83 manchester_baby_instance.BASE_0.s_tickReg VGND VGND VPWR VPWR _0538_
+ sky130_fd_sc_hd__or2b_1
X_0935_ _0454_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_0866_ _0186_ _0394_ _0165_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_21_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0797_ net10 net11 _0129_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ _0116_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_4
X_0582_ net10 net11 _0129_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__or4_4
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0651_ _0198_ _0199_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ clknet_2_3__leaf_clock _0087_ _0038_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.IR.q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1065_ _0536_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
X_0849_ _0116_ _0373_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and3_1
X_0918_ _0434_ _0152_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_3_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 manchester_baby_instance.BASE_0.s_countReg\[2\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0703_ _0138_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nand2_1
X_0565_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] _0101_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__and3b_1
X_0634_ _0173_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ clknet_2_0__leaf_clock _0070_ _0021_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1048_ _0535_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0548_ manchester_baby_instance.CIRCUIT_0.IR.q\[15\] net7 _0104_ VGND VGND VPWR VPWR
+ _0105_ sky130_fd_sc_hd__mux2_1
X_0617_ _0164_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0951_ net12 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] VGND VGND VPWR
+ VPWR _0468_ sky130_fd_sc_hd__or2_1
X_0882_ _0268_ _0125_ _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput18 ram_data_i[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
Xinput29 ram_data_i[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
X_1150_ clknet_2_1__leaf_clock net82 VGND VGND VPWR VPWR manchester_baby_instance.BASE_0.s_countReg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1081_ _0533_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0865_ _0367_ _0169_ _0172_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or3_1
X_0934_ net62 _0453_ _0117_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0796_ _0333_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0581_ net13 net14 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__or2_1
X_0650_ net15 net54 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__or2b_1
X_1133_ clknet_2_1__leaf_clock _0086_ _0037_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfrtp_4
X_1064_ _0536_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0779_ _0184_ _0197_ _0215_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a21o_1
X_0848_ net6 _0127_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nand2_1
X_0917_ net27 _0121_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 manchester_baby_instance.BASE_0.s_tickNext VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0633_ _0174_ _0175_ _0178_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__or4_1
X_0702_ net60 net21 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or2b_1
X_0564_ _0113_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ _0535_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1116_ clknet_2_2__leaf_clock _0069_ _0020_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0616_ net41 net2 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0547_ _0103_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ net12 manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] VGND VGND VPWR
+ VPWR _0467_ sky130_fd_sc_hd__nand2_1
X_0881_ net32 _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__nand2_1
Xinput19 ram_data_i[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
X_1080_ _0533_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0795_ _0205_ _0211_ _0322_ _0307_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__a31o_1
X_0864_ net97 _0118_ _0391_ _0393_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__o22a_1
X_0933_ _0274_ _0448_ _0451_ _0452_ _0146_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0580_ net8 net9 _0127_ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__or4_4
X_1132_ clknet_2_1__leaf_clock _0085_ _0036_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfrtp_1
X_1063_ _0536_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0916_ _0438_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0778_ _0268_ _0132_ _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__and3_1
X_0847_ _0174_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 manchester_baby_instance.BASE_0.s_countReg\[1\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0563_ net100 _0112_ _0104_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
X_0701_ net59 _0248_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0632_ _0179_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ _0535_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_6 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1115_ clknet_2_2__leaf_clock _0068_ _0019_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0546_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\] manchester_baby_instance.CIRCUIT_0.Acc.tick
+ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__and4b_1
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0615_ net42 net3 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1029_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[4\] _0530_ _0531_ manchester_baby_instance.CIRCUIT_0.IR.q\[4\]
+ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__a22o_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_226 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_56 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0880_ net31 _0406_ _0123_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0932_ _0141_ _0145_ _0115_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0794_ _0205_ _0322_ _0211_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a21oi_1
X_0863_ _0288_ _0384_ _0392_ _0275_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1131_ clknet_2_1__leaf_clock _0084_ _0035_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfrtp_1
X_1062_ _0536_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ net67 _0437_ _0117_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_254 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0777_ net16 _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nand2_1
X_0846_ _0191_ _0369_ _0180_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 _0099_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0700_ net59 _0248_ _0235_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0631_ net44 net5 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__and2b_1
X_0562_ net1 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1114_ clknet_2_2__leaf_clock _0067_ _0018_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ _0535_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0829_ _0184_ _0197_ _0215_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0545_ manchester_baby_instance.CIRCUIT_0.IR.q\[14\] manchester_baby_instance.CIRCUIT_0.IR.q\[13\]
+ _0102_ net85 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0614_ _0157_ _0162_ _0158_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__a21oi_1
X_1028_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[3\] _0530_ _0531_ manchester_baby_instance.CIRCUIT_0.IR.q\[3\]
+ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0862_ _0125_ _0126_ net4 VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0931_ net23 _0447_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nand2_1
X_0793_ _0332_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer1 _0121_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_48_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1130_ clknet_2_0__leaf_clock _0083_ _0034_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ _0536_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0914_ _0274_ _0406_ _0433_ _0436_ _0278_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__a32o_1
X_0845_ _0377_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0776_ net15 _0131_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__or2_1
Xclkbuf_2_0__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_0__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0561_ _0111_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_0630_ net5 net44 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1113_ clknet_2_0__leaf_clock _0066_ _0017_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfrtp_1
X_1044_ net33 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0828_ _0362_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_0759_ _0293_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0613_ net68 _0156_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__or2_1
X_0544_ manchester_baby_instance.CIRCUIT_0.Acc.tick manchester_baby_instance.CIRCUIT_0.IR.q\[15\]
+ _0101_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1027_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\] _0530_ _0531_ manchester_baby_instance.CIRCUIT_0.IR.q\[2\]
+ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__a22o_1
XFILLER_0_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer2 net26 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_15_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0792_ net54 _0331_ _0265_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
X_0861_ _0390_ _0271_ _0369_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and3b_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0930_ net96 _0118_ _0446_ _0450_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0536_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0913_ _0149_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__xnor2_1
X_0775_ net89 _0267_ _0314_ _0316_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__o22a_1
X_0844_ net46 _0376_ _0117_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0560_ net106 net12 _0104_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1112_ clknet_2_2__leaf_clock _0065_ _0016_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfrtp_1
X_1043_ _0534_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0827_ net48 _0361_ _0117_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux2_1
X_0758_ _0246_ _0292_ _0240_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_39_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0689_ _0234_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0612_ _0159_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0543_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] VGND VGND VPWR VPWR
+ _0101_ sky130_fd_sc_hd__and3b_1
X_1026_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0530_ _0531_ manchester_baby_instance.CIRCUIT_0.IR.q\[1\]
+ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__a22o_1
XFILLER_0_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ _0481_ _0512_ _0518_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_120 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput70 net70 VGND VGND VPWR VPWR ram_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ _0278_ _0323_ _0328_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a31o_1
X_0860_ _0178_ _0189_ _0368_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0466_ _0471_ _0470_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0912_ _0434_ _0152_ _0150_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0774_ _0288_ _0310_ _0315_ _0276_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__a31o_1
X_0843_ _0115_ _0372_ _0374_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1042_ _0534_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1111_ clknet_2_2__leaf_clock _0064_ _0015_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0688_ _0235_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__nor2_1
X_0826_ _0274_ _0129_ _0358_ _0360_ _0278_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a32o_1
X_0757_ net19 _0133_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0542_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[0\] VGND VGND VPWR
+ VPWR manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0611_ _0148_ _0150_ _0147_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_36_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1025_ _0501_ _0530_ _0531_ manchester_baby_instance.CIRCUIT_0.IR.q\[0\] VGND VGND
+ VPWR VPWR net35 sky130_fd_sc_hd__a22o_1
XFILLER_0_15_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0809_ _0219_ _0220_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0501_ _0483_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput71 net71 VGND VGND VPWR VPWR ram_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput60 net60 VGND VGND VPWR VPWR ram_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0790_ _0116_ _0317_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ _0466_ _0471_ _0470_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0842_ _0127_ _0128_ _0274_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__o21a_1
X_0911_ _0139_ _0140_ _0146_ _0154_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a31o_1
X_0773_ net17 _0132_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ clknet_2_2__leaf_clock _0063_ _0014_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1041_ _0534_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ _0218_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__xnor2_1
X_0756_ net102 _0267_ _0297_ _0300_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__o22a_1
X_0687_ net58 net19 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_46_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0610_ net68 _0156_ _0157_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__a31o_1
X_1024_ _0101_ _0463_ _0485_ _0525_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0808_ net11 _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nand2_1
X_0739_ _0285_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _0477_ _0519_ _0112_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput72 net72 VGND VGND VPWR VPWR ram_rw_en_o sky130_fd_sc_hd__clkbuf_4
Xoutput61 net61 VGND VGND VPWR VPWR ram_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput50 net50 VGND VGND VPWR VPWR ram_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_clock clknet_0_clock VGND VGND VPWR VPWR clknet_2_3__leaf_clock sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0987_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[1\] _0501_ VGND VGND VPWR
+ VPWR _0502_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0910_ net28 _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nand2_1
X_0772_ _0271_ _0292_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__and3_1
X_0841_ net7 _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1040_ _0534_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0755_ _0288_ _0134_ _0299_ _0276_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0824_ _0213_ _0320_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__nand2_1
X_0686_ net19 net58 VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[2\] manchester_baby_instance.CIRCUIT_0.MEMORY_44.countValue\[1\]
+ manchester_baby_instance.CIRCUIT_0.MEMORY_44.s_nextCounterValue\[0\] VGND VGND VPWR
+ VPWR _0530_ sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_36_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0738_ net61 _0284_ _0265_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0807_ net10 _0129_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0669_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_1006_ _0112_ _0501_ _0464_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_20_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput40 net40 VGND VGND VPWR VPWR ram_data_o[0] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 VGND VGND VPWR VPWR stop_lamp_o sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR ram_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput51 net51 VGND VGND VPWR VPWR ram_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0986_ manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[0\] VGND VGND VPWR VPWR
+ _0501_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0840_ net6 _0127_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_1
X_0771_ _0291_ _0244_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0969_ _0462_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0685_ net59 net20 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0823_ net9 _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__nand2_1
X_0754_ net20 _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nand2_1
X_1099_ clknet_2_3__leaf_clock _0052_ _0003_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.ARITH_38.dataB\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1022_ _0529_ VGND VGND VPWR VPWR manchester_baby_instance.CIRCUIT_0.GATES_13.result
+ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_36_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0737_ _0278_ _0279_ _0280_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a31o_1
X_0806_ net90 _0267_ _0341_ _0343_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__o22a_1
X_0668_ net9 net48 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_0599_ net28 net67 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1005_ net64 _0501_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput41 net41 VGND VGND VPWR VPWR ram_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput52 net52 VGND VGND VPWR VPWR ram_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR ram_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

